module adder(G11, G12, G14);
  wire 00, 01, 02, 03, 04, 05, 06, 07, 08, 09, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55;
  input [7:0] G11;
  input [7:0] G12;
  output [7:0] G14;
  lut lut_gate1(0x96, G11[1], G12[1], 49, G14[1]);
  lut lut_gate2(0x8, G11[0], G12[0], 49);
  lut lut_gate3(0x69, G11[2], G12[2], 50, G14[2]);
  lut lut_gate4(0x17, G11[1], G12[1], 49, 50);
  lut lut_gate5(0x69, G11[3], G12[3], 51, G14[3]);
  lut lut_gate6(0x2b, G11[2], G12[2], 50, 51);
  lut lut_gate7(0x69, G11[4], G12[4], 52, G14[4]);
  lut lut_gate8(0x2b, G11[3], G12[3], 51, 52);
  lut lut_gate9(0x69, G11[5], G12[5], 53, G14[5]);
  lut lut_gate10(0x2b, G11[4], G12[4], 52, 53);
  lut lut_gate11(0x69, G11[6], G12[6], 54, G14[6]);
  lut lut_gate12(0x2b, G11[5], G12[5], 53, 54);
  lut lut_gate13(0x69, G11[7], G12[7], 55, G14[7]);
  lut lut_gate14(0x2b, G11[6], G12[6], 54, 55);
  lut lut_gate15(0x6, G11[0], G12[0], G14[0]);

endmodule
