module c432(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G426, G427, G428, G429, G430, G431, G432, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, G203, G213, G308, G318, G358;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G5, G6, G7, G8, G9;
  output G426, G427, G428, G429, G430, G431, G432;
  lut lut_gate1(0xb, 248, 295, G427);
  lut lut_gate2(0x8, 280, 249, 248);
  lut lut_gate3(0x8, 273, 250, 249);
  lut lut_gate4(0x1, 270, 251, 250);
  lut lut_gate5(0x4, 252, G23, 251);
  lut lut_gate6(0x4, G22, 253, 252);
  lut lut_gate7(0x8, G20, G426, 253);
  lut lut_gate8(0xb, 254, 269, G426);
  lut lut_gate9(0x8, 262, 255, 254);
  lut lut_gate10(0x8, 259, 256, 255);
  lut lut_gate11(0x1, 258, 257, 256);
  lut lut_gate12(0x4, G2, G1, 257);
  lut lut_gate13(0x4, G6, G4, 258);
  lut lut_gate14(0x1, 261, 260, 259);
  lut lut_gate15(0x4, G26, G24, 260);
  lut lut_gate16(0x4, G22, G20, 261);
  lut lut_gate17(0x8, 266, 263, 262);
  lut lut_gate18(0x1, 265, 264, 263);
  lut lut_gate19(0x4, G18, G16, 264);
  lut lut_gate20(0x4, G30, G28, 265);
  lut lut_gate21(0x1, 268, 267, 266);
  lut lut_gate22(0x4, G10, G8, 267);
  lut lut_gate23(0x4, G14, G12, 268);
  lut lut_gate24(0x4, G34, G32, 269);
  lut lut_gate25(0x4, 271, G3, 270);
  lut lut_gate26(0x4, G2, 272, 271);
  lut lut_gate27(0x8, G1, G426, 272);
  lut lut_gate28(0x1, 277, 274, 273);
  lut lut_gate29(0x4, 275, G19, 274);
  lut lut_gate30(0x4, G18, 276, 275);
  lut lut_gate31(0x8, G16, G426, 276);
  lut lut_gate32(0x4, 278, G15, 277);
  lut lut_gate33(0x4, G14, 279, 278);
  lut lut_gate34(0x8, G12, G426, 279);
  lut lut_gate35(0x8, 288, 281, 280);
  lut lut_gate36(0x1, 285, 282, 281);
  lut lut_gate37(0x4, 283, G7, 282);
  lut lut_gate38(0x4, G6, 284, 283);
  lut lut_gate39(0x8, G4, G426, 284);
  lut lut_gate40(0x4, 286, G27, 285);
  lut lut_gate41(0x4, G26, 287, 286);
  lut lut_gate42(0x8, G24, G426, 287);
  lut lut_gate43(0x1, 292, 289, 288);
  lut lut_gate44(0x4, 290, G31, 289);
  lut lut_gate45(0x4, G30, 291, 290);
  lut lut_gate46(0x8, G28, G426, 291);
  lut lut_gate47(0x4, 293, G11, 292);
  lut lut_gate48(0x4, G10, 294, 293);
  lut lut_gate49(0x8, G8, G426, 294);
  lut lut_gate50(0x4, 296, G35, 295);
  lut lut_gate51(0x4, G34, 297, 296);
  lut lut_gate52(0x4, G32, 254, 297);
  lut lut_gate53(0x7, 214, 298, G428);
  lut lut_gate54(0x8, 207, 299, 298);
  lut lut_gate55(0x8, 200, 193, 299);
  lut lut_gate56(0x1, 197, 194, 193);
  lut lut_gate57(0x4, 195, G29, 194);
  lut lut_gate58(0x4, 286, 196, 195);
  lut lut_gate59(0x8, G27, G427, 196);
  lut lut_gate60(0x4, 198, G13, 197);
  lut lut_gate61(0x4, 293, 199, 198);
  lut lut_gate62(0x8, G11, G427, 199);
  lut lut_gate63(0x1, 204, 201, 200);
  lut lut_gate64(0x4, 202, G9, 201);
  lut lut_gate65(0x4, 283, 203, 202);
  lut lut_gate66(0x8, G7, G427, 203);
  lut lut_gate67(0x4, 205, G25, 204);
  lut lut_gate68(0x4, 252, 206, 205);
  lut lut_gate69(0x8, G23, G427, 206);
  lut lut_gate70(0x1, 211, 208, 207);
  lut lut_gate71(0x4, 209, G5, 208);
  lut lut_gate72(0x4, 271, 210, 209);
  lut lut_gate73(0x8, G3, G427, 210);
  lut lut_gate74(0x1, G36, 212, 211);
  lut lut_gate75(0xb, 296, 213, 212);
  lut lut_gate76(0x4, G35, 248, 213);
  lut lut_gate77(0x4, 215, 222, 214);
  lut lut_gate78(0x1, 219, 216, 215);
  lut lut_gate79(0x4, 217, G21, 216);
  lut lut_gate80(0x4, 275, 218, 217);
  lut lut_gate81(0x8, G19, G427, 218);
  lut lut_gate82(0x4, 220, G17, 219);
  lut lut_gate83(0x4, 278, 221, 220);
  lut lut_gate84(0x8, G15, G427, 221);
  lut lut_gate85(0x4, 223, G33, 222);
  lut lut_gate86(0x4, 290, 224, 223);
  lut lut_gate87(0x8, G31, G427, 224);
  lut lut_gate88(0xb, 225, 230, G430);
  lut lut_gate89(0x4, 242, 228, 225);
  lut lut_gate90(0x4, 220, 227, 226);
  lut lut_gate91(0x8, G17, G428, 227);
  lut lut_gate92(0x4, 198, 229, 228);
  lut lut_gate93(0x8, G13, G428, 229);
  lut lut_gate94(0x4, 202, 231, 230);
  lut lut_gate95(0x8, G9, G428, 231);
  lut lut_gate96(0x4, 205, 233, 232);
  lut lut_gate97(0x8, G25, G428, 233);
  lut lut_gate98(0x1, 237, 235, 234);
  lut lut_gate99(0x4, 223, 236, 235);
  lut lut_gate100(0x8, G33, G428, 236);
  lut lut_gate101(0x4, 195, 238, 237);
  lut lut_gate102(0x8, G29, G428, 238);
  lut lut_gate103(0x1, 226, 240, 239);
  lut lut_gate104(0x4, 235, 237, 240);
  lut lut_gate105(0x8f, 217, G21, G428, 241);
  lut lut_gate106(0x4, 241, 226, 242);
  lut lut_gate107(0x1f, 242, 232, 237, 243);
  lut lut_gate108(0xef, 243, 230, 228, G431);
  lut lut_gate109(0x8f, 239, 242, 232, 244);
  lut lut_gate110(0xf4, 230, 244, 228, G432);
  lut lut_gate111(0x8f, 209, G5, G428, 245);
  lut lut_gate112(0xf8, 212, G36, G428, 246);
  lut lut_gate113(0x10, 234, 232, G430, 247);
  lut lut_gate114(0x70, 245, 246, 247, G429);

endmodule
