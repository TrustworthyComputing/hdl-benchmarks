module c1908(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893, G1894, G1895, G1896, G1897, G1898, G1899, G19, G1900, G1901, G1902, G1903, G1904, G1905, G1906, G1907, G1908, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G4, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, G313, G314, G315, G316, G317, G318, G319, G320, G321, G322, G323, G324, G325, G326, G327, G328, G335, G338, G341, G344, G347, G350, G356, G359, G362, G368, G374, G377, G395, G398, G401, G404, G407, G410, G413, G416, G419, G425, G428, G431, G437, G440, G443, G446, G449, G452, G455, G458, G467, G470, G473, G476, G479, G482, G485, G488, G491, G494, G497, G500, G506, G509, G512, G515, G518, G521, G524, G527, G530, G715, G716, G718, G719, G720, G721, G723, G728, G772, G774, G776, G778, G780, G782, G784, G786, G787, G789, G790, G792, G795, G805, G807, G808;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G4, G5, G6, G7, G8, G9;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893, G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903, G1904, G1905, G1906, G1907, G1908;
  lut lut_gate1(0xe01f, 273, 266, 264, 237, G1906);
  lut lut_gate2(0x1000, 259, 238, 252, 248, 237);
  lut lut_gate3(0x9009, 243, 247, G28, 239, 238);
  lut lut_gate4(0x1441, 242, 241, 240, G31, 239);
  lut lut_gate5(0x69, G6, G8, G3, 240);
  lut lut_gate6(0x6, G10, G15, 241);
  lut lut_gate7(0xef10, G12, G19, G23, G33, 242);
  lut lut_gate8(0x4114, 246, 245, 244, G31, 243);
  lut lut_gate9(0x69, G9, G14, G16, 244);
  lut lut_gate10(0x10ef, G13, G20, G23, G33, 245);
  lut lut_gate11(0x69, G4, G7, G10, 246);
  lut lut_gate12(0xe0, G19, G31, G23, 247);
  lut lut_gate13(0xeb14, G27, 251, 249, G31, 248);
  lut lut_gate14(0x9669, G11, G15, 250, 244, 249);
  lut lut_gate15(0x10, G18, G24, G33, 250);
  lut lut_gate16(0x96, G2, G5, G8, 251);
  lut lut_gate17(0xeb14, G26, 256, 253, G31, 252);
  lut lut_gate18(0x9, 255, 254, 253);
  lut lut_gate19(0x69, G13, G11, G12, 254);
  lut lut_gate20(0x69, G16, G10, G15, 255);
  lut lut_gate21(0x9, 258, 257, 256);
  lut lut_gate22(0x96, G7, G5, G6, 257);
  lut lut_gate23(0x10ef, G1, G17, G24, G33, 258);
  lut lut_gate24(0x14eb, 263, 262, 260, G31, 259);
  lut lut_gate25(0x6996, G4, G8, 261, 257, 260);
  lut lut_gate26(0x96, G1, G2, G3, 261);
  lut lut_gate27(0x4bb4, G9, 255, G21, G33, 262);
  lut lut_gate28(0xe0, G17, G31, G24, 263);
  lut lut_gate29(0x0100, 238, 265, 252, 248, 264);
  lut lut_gate30(0xe0, G18, G31, G24, 265);
  lut lut_gate31(0x0, 270, 267, 272, 266);
  lut lut_gate32(0x4b, G25, 268, G31, 267);
  lut lut_gate33(0x9669, 269, 261, 255, 254, 268);
  lut lut_gate34(0xb44b, G4, G14, G22, G33, 269);
  lut lut_gate35(0x0b, 271, G24, G23, 270);
  lut lut_gate36(0xffe0, G33, G32, G31, G29, 271);
  lut lut_gate37(0xe0, G20, G31, G23, 272);
  lut lut_gate38(0x10ea, 260, G29, G21, G33, 273);
  lut lut_gate39(0xe01f, G1, 266, 264, 237, G1884);
  lut lut_gate40(0xe01f, G2, 266, 264, 237, G1885);
  lut lut_gate41(0xe01f, G3, 266, 264, 237, G1886);
  lut lut_gate42(0xe01f, G4, 266, 264, 237, G1887);
  lut lut_gate43(0xe01f, G10, 220, 264, 237, G1888);
  lut lut_gate44(0x0, 221, 267, 272, 220);
  lut lut_gate45(0x0b, 222, G24, G23, 221);
  lut lut_gate46(0xffe0, G33, G32, G30, G31, 222);
  lut lut_gate47(0xe01f, G15, 220, 264, 237, G1889);
  lut lut_gate48(0xe01f, G16, 220, 264, 237, G1890);
  lut lut_gate49(0x9, G5, 223, G1891);
  lut lut_gate50(0xe000, 270, 224, 237, 264, 223);
  lut lut_gate51(0x8, 272, 267, 224);
  lut lut_gate52(0x9, G6, 223, G1892);
  lut lut_gate53(0x9, G7, 223, G1893);
  lut lut_gate54(0x9, G8, 223, G1894);
  lut lut_gate55(0x87, G9, 221, 225, G1895);
  lut lut_gate56(0xe0, 224, 237, 264, 225);
  lut lut_gate57(0x9, G11, 226, G1896);
  lut lut_gate58(0x80, 265, 220, 237, 226);
  lut lut_gate59(0x9, G12, 226, G1897);
  lut lut_gate60(0x9, G13, 226, G1898);
  lut lut_gate61(0x9, G14, 226, G1899);
  lut lut_gate62(0xfff2, 228, G33, 227, G32, G1900);
  lut lut_gate63(0x111f, 264, 237, 220, 266, 227);
  lut lut_gate64(0x4000, 264, 267, 259, 272, 228);
  lut lut_gate65(0xe01f, 229, 220, 264, 237, G1907);
  lut lut_gate66(0x10ea, 230, G30, G22, G33, 229);
  lut lut_gate67(0x69, G9, G14, 253, 230);
  lut lut_gate68(0x0b04, 231, 232, 263, 227, G1901);
  lut lut_gate69(0x6, 262, 260, 231);
  lut lut_gate70(0x1, G32, G33, 232);
  lut lut_gate71(0x0b04, 268, 232, G25, 227, G1902);
  lut lut_gate72(0x07, 232, 233, 227, G1903);
  lut lut_gate73(0x6, 251, 249, 233);
  lut lut_gate74(0x0, 232, 234, 227, G1904);
  lut lut_gate75(0x96, 242, 241, 240, 234);
  lut lut_gate76(0x0, 232, 235, 227, G1905);
  lut lut_gate77(0x69, 246, 245, 244, 235);
  lut lut_gate78(0x40, 236, 227, 232, G1908);
  lut lut_gate79(0x6, 256, 253, 236);

endmodule
