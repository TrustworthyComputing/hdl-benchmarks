module c7552(N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342, N241_O);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, 0950, 0951, 0952, 0953, 0954, 0955, 0956, 0957, 0958, 0959, 0960, 0961, 0962, 0963, 0964, 0965, 0966, 0967, 0968, 0969, 0970, 0971, 0972, 0973, 0974, 0975, 0976, 0977, 0978, 0979, 0980, 0981, 0982, 0983, 0984, 0985, 0986, 0987, 0988, 0989, 0990, 0991, 0992, 0993, 0994, 0995, 0996, 0997, 0998, 0999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165, 1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187, 1188, 1189, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198, 1199, 1200, 1201, 1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209, 1210, 1211, 1212, 1213, 1214, 1215, 1216, 1217, 1218, 1219, 1220, 1221, 1222, 1223, 1224, 1225, 1226, 1227, 1228, 1229, 1230, 1231, 1232, 1233, 1234, 1235, 1236, 1237, 1238, 1239, 1240, 1241, 1242, 1243, 1244, 1245, 1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264, 1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 1274, 1275, 1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 1286, 1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297, 1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308, 1309, 1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319, 1320, 1321, 1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361, 1362, 1363, 1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371, 1372, 1373, 1374, 1375, 1376, 1377, 1378, 1379, 1380, 1381, 1382, 1383, 1384, 1385, 1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 1394, 1395, 1396, 1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 1418, 1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429, 1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440, 1441, 1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451, 1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495, 1496, 1497, 1498, 1499, 1500, 1501, 1502, 1503, 1504, 1505, 1506, 1507, 1508, 1509, 1510, 1511, 1512, 1513, 1514, 1515, 1516, 1517, 1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550, 1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561, 1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572, 1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1601, 1602, 1603, 1604, 1605, 1606, 1607, 1608, 1609, 1610, 1611, 1612, 1613, 1614, 1615, 1616, 1617, 1618, 1619, 1620, 1621, 1622, 1623, 1624, 1625, 1626, 1627, 1628, 1629, 1630, 1631, 1632, 1633, 1634, 1635, 1636, 1637, 1638, 1639, 1640, 1641, 1642, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1651, 1652, 1653, 1654, 1655, 1656, 1657, 1658, 1659, 1660, 1661, 1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 1670, 1671, 1672, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1681, 1682, 1683, 1684, 1685, 1686, 1687, 1688, 1689, 1690, 1691, 1692, 1693, 1694, 1695, 1696, 1697, 1698, 1699, 1700, 1701, 1702, 1703, 1704, 1705, 1706, 1707, 1708, 1709, 1710, 1711, 1712, 1713, 1714, 1715, 1716, 1717, 1718, 1719, 1720, 1721, 1722, 1723, 1724, 1725, 1726, 1727, 1728, 1729, 1730, 1731, 1732, 1733, 1734, 1735, 1736, 1737, 1738, 1739, 1740, 1741, 1742, 1743, 1744, 1745, 1746, 1747, 1748, 1749, 1750, 1751, 1752, 1753, 1754, 1755, 1756, 1757, 1758, 1759, 1760, 1761, 1762, 1763, 1764, 1765, 1766, 1767, 1768, 1769, 1770, 1771, 1772, 1773, 1774, 1775, 1776, 1777, 1778, N10778, N10781, N1116, N1125, N1136, N1147, N1160, N1175, N1182, N1233, N1244, N1249, N1256, N1270, N1277, N1287, N1299, N1308, N1311, N1428, N1431, N1828, N1829, N1830, N1833, N1840, N1841, N1842, N1843, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1913, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1997, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2240, N2267, N2275, N2287, N2293, N2309, N2315, N2331, N2347, N2368, N2384, N2390, N2406, N2412, N590, N614, N625, N636, N657, N676, N682, N689, N750, N871;
  input N1, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N12, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N15, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N18, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N23, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241_I, N242, N245, N248, N251, N254, N257, N26, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N29, N293, N296, N299, N303, N307, N310, N313, N316, N319, N32, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N35, N352, N355, N358, N361, N364, N367, N38, N382, N41, N44, N47, N5, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N9, N94, N97;
  output N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N1110, N1111, N1112, N1113, N1114, N11333, N11334, N11340, N11342, N1489, N1490, N1781, N241_O, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945;
  lut lut_gate1(0xb, N242, N5, N1110);
  lut lut_gate2(0xe, N57, N5, N881);
  lut lut_gate3(0x7fff, N240, N228, N150, N184, N882);
  lut lut_gate4(0x7fff, N230, N218, N210, N152, N883);
  lut lut_gate5(0x7fff, N186, N185, N183, N182, N884);
  lut lut_gate6(0x7fff, N199, N188, N162, N172, N885);
  lut lut_gate7(0xbf, N134, N133, N5, N1113);
  lut lut_gate8(0x6, N367, 1433, N10025);
  lut lut_gate9(0xeb, N310, N41, N18, 1433);
  lut lut_gate10(0x8e71, 1443, 1444, N319, 1434, N10109);
  lut lut_gate11(0x07, 1435, 1440, N367, 1434);
  lut lut_gate12(0x1, 1439, 1436, 1435);
  lut lut_gate13(0x7100, 1441, N313, 1438, 1437, 1436);
  lut lut_gate14(0x10, N41, N310, N18, 1437);
  lut lut_gate15(0xca, N18, N238, N29, 1438);
  lut lut_gate16(0x3500, N316, N18, N237, N26, 1439);
  lut lut_gate17(0x80, 1442, 1441, 1433, 1440);
  lut lut_gate18(0xac53, N316, N18, N26, N237, 1441);
  lut lut_gate19(0xac53, N313, N18, N29, N238, 1442);
  lut lut_gate20(0xac53, N322, N18, N103, N235, 1443);
  lut lut_gate21(0xca, N18, N236, N23, 1444);
  lut lut_gate22(0x9, 1445, 1434, N10110);
  lut lut_gate23(0xac53, N319, N18, N23, N236, 1445);
  lut lut_gate24(0x708f, 1441, 1447, 1442, 1446, N10111);
  lut lut_gate25(0x8, N367, 1433, 1446);
  lut lut_gate26(0x71, N313, 1438, 1437, 1447);
  lut lut_gate27(0x1e, 1442, 1437, 1446, N10112);
  lut lut_gate28(0x8, N12, N9, 1448);
  lut lut_gate29(0x0b, 1448, N18, N157, 1449);
  lut lut_gate30(0xca, N18, N158, N135, 1450);
  lut lut_gate31(0x96, 1455, 1454, 1452, 1451);
  lut lut_gate32(0x53ac, 1453, N18, N141, N161, 1452);
  lut lut_gate33(0x35, N18, N151, N147, 1453);
  lut lut_gate34(0x35, N18, N159, N144, 1454);
  lut lut_gate35(0x35, N18, N160, N138, 1455);
  lut lut_gate36(0x69, N209, N211, N212, 1456);
  lut lut_gate37(0x96, 1464, 1463, 1458, 1457);
  lut lut_gate38(0x96, 1462, 1461, 1459, 1458);
  lut lut_gate39(0x53ac, 1460, N18, N115, N227, 1459);
  lut lut_gate40(0xca, N18, N217, N118, 1460);
  lut lut_gate41(0xca, N18, N223, N47, 1461);
  lut lut_gate42(0xca, N18, N224, N121, 1462);
  lut lut_gate43(0xca, N18, N225, N94, 1463);
  lut lut_gate44(0xca, N18, N226, N97, 1464);
  lut lut_gate45(0x9669, 1475, 1474, 1471, 1466, 1465);
  lut lut_gate46(0x9669, 1444, 1470, 1469, 1467, 1466);
  lut lut_gate47(0x53ac, 1468, N18, N44, N239, 1467);
  lut lut_gate48(0x53, N18, N41, N229, 1468);
  lut lut_gate49(0xac53, 1438, N18, N26, N237, 1469);
  lut lut_gate50(0xca, N18, N235, N103, 1470);
  lut lut_gate51(0x9, 1473, 1472, 1471);
  lut lut_gate52(0x35, N18, N231, N100, 1472);
  lut lut_gate53(0x35, N18, N232, N124, 1473);
  lut lut_gate54(0xca, N18, N233, N127, 1474);
  lut lut_gate55(0xca, N18, N234, N130, 1475);
  lut lut_gate56(0x6996, 1480, 1479, 1478, 1477, 1476);
  lut lut_gate57(0xca, N18, N221, N32, 1477);
  lut lut_gate58(0xca, N18, N222, N35, 1478);
  lut lut_gate59(0xca, N18, N219, N66, 1479);
  lut lut_gate60(0xca, N18, N220, N50, 1480);
  lut lut_gate61(0xbf, 1481, 1505, 1518, N10575);
  lut lut_gate62(0x1441, 1500, 1497, 1492, 1482, 1481);
  lut lut_gate63(0x6996, 1491, 1490, 1488, 1483, 1482);
  lut lut_gate64(0x96, 1487, 1486, 1484, 1483);
  lut lut_gate65(0xa35c, 1485, N18, N114, N248, 1484);
  lut lut_gate66(0x3a, N18, N251, N113, 1485);
  lut lut_gate67(0xc5, N18, N260, N88, 1486);
  lut lut_gate68(0xc5, N18, N257, N112, 1487);
  lut lut_gate69(0xc355, N18, N267, N263, 1489, 1488);
  lut lut_gate70(0x6, N271, N245, 1489);
  lut lut_gate71(0x3a, N18, N106, N87, 1490);
  lut lut_gate72(0x3a, N18, N254, N111, 1491);
  lut lut_gate73(0x96, 1496, 1495, 1493, 1492);
  lut lut_gate74(0xa35c, 1494, N18, N82, N274, 1493);
  lut lut_gate75(0xc5, N18, N277, N65, 1494);
  lut lut_gate76(0xc5, N18, N289, N64, 1495);
  lut lut_gate77(0xc5, N18, N286, N85, 1496);
  lut lut_gate78(0x9, 1499, 1498, 1497);
  lut lut_gate79(0x3a, N18, N283, N84, 1498);
  lut lut_gate80(0xc5, N18, N280, N83, 1499);
  lut lut_gate81(0x9669, 1504, 1503, 1502, 1501, 1500);
  lut lut_gate82(0x3a, N18, N296, N86, 1501);
  lut lut_gate83(0x3a, N18, N293, N63, 1502);
  lut lut_gate84(0x3a, N18, N303, N110, 1503);
  lut lut_gate85(0xc5, N18, N299, N109, 1504);
  lut lut_gate86(0x6996, 1517, 1516, 1514, 1506, 1505);
  lut lut_gate87(0x69, 1513, 1512, 1507, 1506);
  lut lut_gate88(0x9669, 1511, 1510, 1509, 1508, 1507);
  lut lut_gate89(0xc5, N18, N331, N55, 1508);
  lut lut_gate90(0xc5, N18, N328, N54, 1509);
  lut lut_gate91(0xc5, N18, N325, N53, 1510);
  lut lut_gate92(0x3a, N18, N334, N56, 1511);
  lut lut_gate93(0x3a, N18, N322, N73, 1512);
  lut lut_gate94(0xc5, N18, N319, N75, 1513);
  lut lut_gate95(0x5ca3, 1515, N18, N70, N310, 1514);
  lut lut_gate96(0x3a, N18, N307, N69, 1515);
  lut lut_gate97(0x3a, N18, N316, N76, 1516);
  lut lut_gate98(0xc5, N18, N313, N74, 1517);
  lut lut_gate99(0x9669, 1530, 1529, 1528, 1519, 1518);
  lut lut_gate100(0x6996, 1527, 1526, 1524, 1520, 1519);
  lut lut_gate101(0x69, 1523, 1522, 1521, 1520);
  lut lut_gate102(0x3a, N18, N352, N80, 1521);
  lut lut_gate103(0xc5, N18, N349, N81, 1522);
  lut lut_gate104(0xc5, N18, N355, N79, 1523);
  lut lut_gate105(0xa35c, 1525, N18, N58, N337, 1524);
  lut lut_gate106(0xc5, N18, N340, N77, 1525);
  lut lut_gate107(0xc5, N18, N346, N59, 1526);
  lut lut_gate108(0xc5, N18, N343, N78, 1527);
  lut lut_gate109(0xc5, N18, N364, N62, 1528);
  lut lut_gate110(0xc5, N18, N361, N61, 1529);
  lut lut_gate111(0x3a, N18, N358, N60, 1530);
  lut lut_gate112(0x0b, 1448, N18, N177, 1531);
  lut lut_gate113(0xca, N18, N178, N135, 1532);
  lut lut_gate114(0x35, N18, N171, N147, 1533);
  lut lut_gate115(0x35, N18, N179, N144, 1534);
  lut lut_gate116(0x35, N18, N180, N138, 1535);
  lut lut_gate117(0x69, 1547, 1542, 1537, 1536);
  lut lut_gate118(0x6996, 1541, 1540, 1539, 1538, 1537);
  lut lut_gate119(0xca, N18, N193, N47, 1538);
  lut lut_gate120(0xca, N18, N194, N121, 1539);
  lut lut_gate121(0xca, N18, N195, N94, 1540);
  lut lut_gate122(0xca, N18, N196, N97, 1541);
  lut lut_gate123(0x9669, 1546, 1545, 1544, 1543, 1542);
  lut lut_gate124(0xca, N18, N191, N32, 1543);
  lut lut_gate125(0xca, N18, N192, N35, 1544);
  lut lut_gate126(0xca, N18, N189, N66, 1545);
  lut lut_gate127(0xca, N18, N190, N50, 1546);
  lut lut_gate128(0xac53, 1548, N18, N115, N197, 1547);
  lut lut_gate129(0xca, N18, N187, N118, 1548);
  lut lut_gate130(0x6996, 1553, 1552, 1551, 1550, 1549);
  lut lut_gate131(0xca, N18, N206, N26, 1550);
  lut lut_gate132(0xca, N18, N207, N29, 1551);
  lut lut_gate133(0xca, N18, N204, N103, 1552);
  lut lut_gate134(0xca, N18, N205, N23, 1553);
  lut lut_gate135(0x9669, 1558, 1557, 1556, 1555, 1554);
  lut lut_gate136(0xca, N18, N202, N127, 1555);
  lut lut_gate137(0xca, N18, N203, N130, 1556);
  lut lut_gate138(0x35, N18, N200, N100, 1557);
  lut lut_gate139(0x35, N18, N201, N124, 1558);
  lut lut_gate140(0x69, N170, N164, N165, 1559);
  lut lut_gate141(0x6, 1592, 1560, N10632);
  lut lut_gate142(0x222b, 1591, 1561, N364, 1479, 1560);
  lut lut_gate143(0x4f00, 1589, 1587, 1562, 1566, 1561);
  lut lut_gate144(0x71, N352, 1461, 1563, 1562);
  lut lut_gate145(0xb2, 1462, N349, 1564, 1563);
  lut lut_gate146(0xb2, 1463, N346, 1565, 1564);
  lut lut_gate147(0x2b22, 1460, N340, N343, 1464, 1565);
  lut lut_gate148(0x2b00, 1567, N334, 1472, 1574, 1566);
  lut lut_gate149(0x80, 1573, 1572, 1568, 1567);
  lut lut_gate150(0x80, 1571, 1570, 1569, 1568);
  lut lut_gate151(0x9, N340, 1460, 1569);
  lut lut_gate152(0x9, N346, 1463, 1570);
  lut lut_gate153(0x9, N343, 1464, 1571);
  lut lut_gate154(0x9, N352, 1461, 1572);
  lut lut_gate155(0x9, N349, 1462, 1573);
  lut lut_gate156(0x00ef, 1578, 1582, 1586, 1575, 1574);
  lut lut_gate157(0x2b, N331, 1473, 1576, 1575);
  lut lut_gate158(0xb2, 1577, N328, 1474, 1576);
  lut lut_gate159(0x0c0a, N18, N325, N234, N130, 1577);
  lut lut_gate160(0x00, 1579, N331, 1473, 1576, 1578);
  lut lut_gate161(0x9000, 1580, 1581, N325, 1475, 1579);
  lut lut_gate162(0xac53, N331, N18, N124, N232, 1580);
  lut lut_gate163(0xac53, N328, N18, N127, N233, 1581);
  lut lut_gate164(0xef00, 1583, 1585, 1439, 1436, 1582);
  lut lut_gate165(0x71, N322, 1584, 1470, 1583);
  lut lut_gate166(0x0c0a, N18, N319, N236, N23, 1584);
  lut lut_gate167(0x8, 1445, 1443, 1585);
  lut lut_gate168(0x80, N367, 1585, 1440, 1586);
  lut lut_gate169(0x90, 1588, N355, 1478, 1587);
  lut lut_gate170(0x9, N358, 1477, 1588);
  lut lut_gate171(0xb0, 1590, 1480, N361, 1589);
  lut lut_gate172(0x4, 1478, N355, N358, 1477, 1590);
  lut lut_gate173(0x4, N361, 1480, 1591);
  lut lut_gate174(0x6, N277, 1453, 1592);
  lut lut_gate175(0x9, 1618, 1593, N10641);
  lut lut_gate176(0x70, 1613, 1594, 1617, 1593);
  lut lut_gate177(0x0e00, 1605, 1595, 1560, 1596, 1594);
  lut lut_gate178(0x007f, 1596, 1603, 1600, 1604, 1595);
  lut lut_gate179(0xb2, 1449, N289, 1597, 1596);
  lut lut_gate180(0x71, 1450, N286, 1598, 1597);
  lut lut_gate181(0x4, N283, 1454, 1599, 1598);
  lut lut_gate182(0x1117, 1453, N277, N280, 1455, 1599);
  lut lut_gate183(0x80, 1602, 1601, 1592, 1600);
  lut lut_gate184(0x6, N283, 1454, 1601);
  lut lut_gate185(0x6, N280, 1455, 1602);
  lut lut_gate186(0x9, N289, 1449, 1603);
  lut lut_gate187(0x9, N286, 1450, 1604);
  lut lut_gate188(0x80, 1611, 1608, 1606, 1605);
  lut lut_gate189(0x9, N296, 1607, 1606);
  lut lut_gate190(0x0b, 1448, N18, N155, 1607);
  lut lut_gate191(0x1, 1610, 1609, 1608);
  lut lut_gate192(0x000b, N293, 1448, N18, N156, 1609);
  lut lut_gate193(0xf400, N293, 1448, N18, N156, 1610);
  lut lut_gate194(0x9, N299, 1612, 1611);
  lut lut_gate195(0x0b, 1448, N18, N154, 1612);
  lut lut_gate196(0xb2, N303, 1616, 1614, 1613);
  lut lut_gate197(0xb2, N299, 1612, 1615, 1614);
  lut lut_gate198(0x71, N296, 1609, 1607, 1615);
  lut lut_gate199(0x0b, 1448, N18, N153, 1616);
  lut lut_gate200(0x9, N303, 1616, 1617);
  lut lut_gate201(0x1, 1620, 1619, 1618);
  lut lut_gate202(0x000b, N251, 1448, N18, N209, 1619);
  lut lut_gate203(0xf400, N251, 1448, N18, N209, 1620);
  lut lut_gate204(0xf40b, 1604, 1621, 1598, 1560, N10712);
  lut lut_gate205(0x4, 1598, 1600, 1621);
  lut lut_gate206(0xe1, 1603, 1623, 1622, N10711);
  lut lut_gate207(0x0b00, 1598, 1560, 1450, N286, 1622);
  lut lut_gate208(0xb2, N286, 1450, 1621, 1623);
  lut lut_gate209(0x1fe0, 1601, 1624, 1599, 1560, N10713);
  lut lut_gate210(0x17, N280, 1455, 1625, 1624);
  lut lut_gate211(0x8, N277, 1453, 1625);
  lut lut_gate212(0x42b, 1602, N277, 1453, 1560, N10714);
  lut lut_gate213(0x1e, 1637, 1634, 1626, N10715);
  lut lut_gate214(0x8f00, 1627, 1613, 1617, 1594, 1626);
  lut lut_gate215(0x8000, 1632, 1630, 1628, 1618, 1627);
  lut lut_gate216(0x9, N254, 1629, 1628);
  lut lut_gate217(0x0b, 1448, N18, N216, 1629);
  lut lut_gate218(0x9, N106, 1631, 1630);
  lut lut_gate219(0x0b, 1448, N18, N215, 1631);
  lut lut_gate220(0x9, N257, 1633, 1632);
  lut lut_gate221(0x0b, 1448, N18, N214, 1633);
  lut lut_gate222(0x71, 1633, N257, 1635, 1634);
  lut lut_gate223(0x71, N106, 1631, 1636, 1635);
  lut lut_gate224(0xb2, 1619, N254, 1629, 1636);
  lut lut_gate225(0x9, N260, 1638, 1637);
  lut lut_gate226(0x0b, 1448, N18, N213, 1638);
  lut lut_gate227(0xf807, 1632, 1639, 1635, 1593, N10716);
  lut lut_gate228(0x7f00, 1635, 1628, 1618, 1630, 1639);
  lut lut_gate229(0x07f8, 1630, 1636, 1628, 1640, N10717);
  lut lut_gate230(0x4, 1618, 1593, 1640);
  lut lut_gate231(0x1e, 1628, 1619, 1640, N10718);
  lut lut_gate232(0xfeff, 1641, N10576, N10574, N10575, N10729);
  lut lut_gate233(0x0001, N885, N884, N883, N882, 1641);
  lut lut_gate234(0x6, 1569, 1642, N10827);
  lut lut_gate235(0x2b, N334, 1472, 1574, 1642);
  lut lut_gate236(0xb4, 1572, 1644, 1643, N10868);
  lut lut_gate237(0x000b, 1564, 1642, 1462, N349, 1643);
  lut lut_gate238(0xa8fe, N349, 1564, 1568, 1462, 1644);
  lut lut_gate239(0x1e, 1573, 1564, 1645, N10869);
  lut lut_gate240(0x8000, 1571, 1570, 1569, 1642, 1645);
  lut lut_gate241(0xf10e, 1570, 1646, 1565, 1642, N10870);
  lut lut_gate242(0x7150, N340, N343, 1460, 1464, 1646);
  lut lut_gate243(0x4, 1571, 1460, N340, 1642, N10871);
  lut lut_gate244(0x8, N163, N1, N1781);
  lut lut_gate245(0xf710, N38, 1647, 1649, 1648, N10101);
  lut lut_gate246(0xa8fe, N260, 1626, 1634, 1638, 1647);
  lut lut_gate247(0x8, N382, N263, 1648);
  lut lut_gate248(0x8, N382, N267, 1649);
  lut lut_gate249(0xef, 1693, 1699, 1650, N10102);
  lut lut_gate250(0x8f00, 1666, 1686, 1692, N10704, 1650);
  lut lut_gate251(0x01, N89, N70, N18, N41, 1651);
  lut lut_gate252(0xbbb0, 1552, 1512, 1513, 1553, 1652);
  lut lut_gate253(0x4, 1553, 1552, 1513, 1512, 1653);
  lut lut_gate254(0x6, 1558, 1508, 1654);
  lut lut_gate255(0x4f00, 1662, 1661, 1656, 1658, 1655);
  lut lut_gate256(0x60, 1657, 1538, 1521, 1656);
  lut lut_gate257(0xb00b, 1539, 1522, 1526, 1540, 1657);
  lut lut_gate258(0x0071, 1660, 1527, 1541, 1659, 1658);
  lut lut_gate259(0x4, 1548, 1525, 1659);
  lut lut_gate260(0x4, 1540, 1526, 1660);
  lut lut_gate261(0x4, 1539, 1538, 1522, 1521, 1661);
  lut lut_gate262(0x0990, 1543, 1530, 1544, 1523, 1662);
  lut lut_gate263(0x4, 1544, 1543, 1523, 1530, 1663);
  lut lut_gate264(0x41, 1541, 1527, 1660, 1664);
  lut lut_gate265(0x222b, 1558, 1508, 1557, 1511, 1665);
  lut lut_gate266(0x80, 1683, 1680, 1667, 1666);
  lut lut_gate267(0x8000, 1678, 1677, 1673, 1668, 1667);
  lut lut_gate268(0x90, 1669, 1487, 1672, 1668);
  lut lut_gate269(0xeee0, 1490, 1670, 1491, 1671, 1669);
  lut lut_gate270(0x0b, 1448, N18, N168, 1670);
  lut lut_gate271(0x0b, 1448, N18, N169, 1671);
  lut lut_gate272(0x0b, 1448, N18, N167, 1672);
  lut lut_gate273(0x000b, 1675, 1674, 1448, 1485, 1673);
  lut lut_gate274(0x8, 1490, 1670, 1674);
  lut lut_gate275(0x4, 1676, 1486, 1675);
  lut lut_gate276(0x0b, 1448, N18, N166, 1676);
  lut lut_gate277(0x0bbb, 1491, 1671, 1485, 1448, 1677);
  lut lut_gate278(0x0, 1679, 1676, 1486, 1678);
  lut lut_gate279(0x108f, N38, N382, N271, N245, 1679);
  lut lut_gate280(0x4182, 1503, 1504, 1682, 1681, 1680);
  lut lut_gate281(0x0b, 1448, N18, N173, 1681);
  lut lut_gate282(0x0b, 1448, N18, N174, 1682);
  lut lut_gate283(0x1428, 1501, 1502, 1685, 1684, 1683);
  lut lut_gate284(0x0b, 1448, N18, N175, 1684);
  lut lut_gate285(0x0b, 1448, N18, N176, 1685);
  lut lut_gate286(0xb0, 1691, 1687, 1688, 1686);
  lut lut_gate287(0x9009, 1532, 1496, 1495, 1531, 1687);
  lut lut_gate288(0x00ef, 1690, 1689, 1533, 1494, 1688);
  lut lut_gate289(0x0990, 1535, 1499, 1534, 1498, 1689);
  lut lut_gate290(0x222b, 1535, 1499, 1534, 1498, 1690);
  lut lut_gate291(0x4, 1532, 1496, 1495, 1531, 1691);
  lut lut_gate292(0x6000, 1689, 1687, 1533, 1494, 1692);
  lut lut_gate293(0x0, 1694, 1697, 1678, 1693);
  lut lut_gate294(0xf800, 1667, 1695, 1696, 1680, 1694);
  lut lut_gate295(0xb2a0, 1682, 1503, 1504, 1681, 1695);
  lut lut_gate296(0xe888, 1502, 1685, 1501, 1684, 1696);
  lut lut_gate297(0x00b2, 1675, 1487, 1672, 1698, 1697);
  lut lut_gate298(0x0, 1674, 1677, 1669, 1698);
  lut lut_gate299(0xef00, N38, N382, N245, N271, 1699);
  lut lut_gate300(0x6, 1700, 1574, N10350);
  lut lut_gate301(0x6, N334, 1472, 1700);
  lut lut_gate302(0x1e, 1580, 1576, 1701, N10351);
  lut lut_gate303(0x4100, 1581, N325, 1475, 1702, 1701);
  lut lut_gate304(0x4, 1582, 1586, 1702);
  lut lut_gate305(0xb24, 1581, N325, 1475, 1702, N10352);
  lut lut_gate306(0x96, N325, 1475, 1702, N10353);
  lut lut_gate307(0x4b, 1617, 1614, 1594, N10760);
  lut lut_gate308(0x4b, 1611, 1615, 1703, N10761);
  lut lut_gate309(0x40, 1608, 1606, 1704, 1703);
  lut lut_gate310(0xf1, 1595, 1596, 1560, 1704);
  lut lut_gate311(0xf20, 1606, 1610, 1609, 1704, N10762);
  lut lut_gate312(0x9, 1608, 1704, N10763);
  lut lut_gate313(0x35, 1647, 1706, 1705, N10837);
  lut lut_gate314(0x78, 1649, N38, 1648, 1705);
  lut lut_gate315(0xe1, 1649, N38, 1648, 1706);
  lut lut_gate316(0x69, N38, 1648, 1647, N10839);
  lut lut_gate317(0xe1, 1707, 1591, 1561, N10905);
  lut lut_gate318(0x9, N364, 1479, 1707);
  lut lut_gate319(0x96, N361, 1480, 1708, N10906);
  lut lut_gate320(0x70, 1590, 1709, 1587, 1708);
  lut lut_gate321(0xb, 1562, 1566, 1709);
  lut lut_gate322(0x4, 1588, 1478, N355, 1709, N10907);
  lut lut_gate323(0x69, N355, 1478, 1709, N10908);
  lut lut_gate324(0xe7, N296, 1610, 1607, 1710);
  lut lut_gate325(0x6996, 1604, 1602, 1601, 1603, 1711);
  lut lut_gate326(0x42b, 1621, N280, 1455, 1625, 1712);
  lut lut_gate327(0x96, 1599, 1598, 1597, 1713);
  lut lut_gate328(0xa35c, 1714, 1647, 1706, 1705, N11334);
  lut lut_gate329(0x5ca3, 1721, 1593, 1715, 1718, 1714);
  lut lut_gate330(0x69, 1618, 1717, 1716, 1715);
  lut lut_gate331(0x1, 1627, 1634, 1716);
  lut lut_gate332(0xe178, N254, 1639, 1620, 1629, 1717);
  lut lut_gate333(0x55c3, 1618, 1716, 1717, 1719, 1718);
  lut lut_gate334(0x9, 1720, 1634, 1719);
  lut lut_gate335(0x4b, 1635, 1629, N254, 1720);
  lut lut_gate336(0x9669, 1632, 1630, 1628, 1637, 1721);
  lut lut_gate337(0x9669, 1573, 1572, 1571, 1570, 1722);
  lut lut_gate338(0x69, 1646, 1724, 1644, 1723);
  lut lut_gate339(0xaf, 1564, N340, 1568, 1460, 1724);
  lut lut_gate340(0x6, 1726, 1563, 1725);
  lut lut_gate341(0x4b, 1564, 1464, N343, 1726);
  lut lut_gate342(0xa33c, N367, 1433, 1728, 1731, 1727);
  lut lut_gate343(0x96, 1730, 1435, 1729, 1728);
  lut lut_gate344(0x71, N319, 1444, 1435, 1729);
  lut lut_gate345(0x18, 1438, N313, 1437, 1730);
  lut lut_gate346(0x708f, 1732, 1729, 1445, 1440, 1731);
  lut lut_gate347(0xc1, 1733, 1435, 1440, 1732);
  lut lut_gate348(0x70, 1447, 1433, 1442, 1733);
  lut lut_gate349(0x6, 1580, 1700, 1734);
  lut lut_gate350(0xb42b, N325, 1475, N328, 1474, 1735);
  lut lut_gate351(0x2b, N325, 1475, N328, 1474, 1736);
  lut lut_gate352(0x9669, 1445, 1442, 1441, 1443, 1737);
  lut lut_gate353(0x1, N15, N1111);
  lut lut_gate354(0xf710, N38, 1647, 1649, 1648, N10104);
  lut lut_gate355(0xf710, N38, 1647, 1649, 1648, N10706);
  lut lut_gate356(0xf710, N38, 1647, 1649, 1648, N10759);
  lut lut_gate357(0x6996, N213, N214, N215, N216, 1738);
  lut lut_gate358(0xebff, N18, 1456, 1738, 1448, 1739);
  lut lut_gate359(0x1400, 1739, 1476, 1457, 1465, 1740);
  lut lut_gate360(0x6996, N166, N167, N168, N169, 1741);
  lut lut_gate361(0xebff, N18, 1559, 1741, 1448, 1742);
  lut lut_gate362(0x6996, 1535, 1534, 1533, 1532, 1743);
  lut lut_gate363(0x5ca3, 1743, N18, N141, N181, 1744);
  lut lut_gate364(0x6996, N177, N173, N174, N175, 1745);
  lut lut_gate365(0xb2, 1749, 1556, 1510, 1746);
  lut lut_gate366(0xb0ff, 1768, 1752, 1765, 1665, N10704);
  lut lut_gate367(0x8e71, 1516, 1551, 1651, 1517, 1747);
  lut lut_gate368(0x53ff, 1652, 1747, 1516, 1550, 1748);
  lut lut_gate369(0x8, 1653, 1748, 1749);
  lut lut_gate370(0x9009, 1546, 1529, 1545, 1528, 1750);
  lut lut_gate371(0x9000, 1662, 1750, 1548, 1525, 1751);
  lut lut_gate372(0x80, 1664, 1656, 1751, 1752);
  lut lut_gate373(0xc5, 1560, 1595, 1596, 1753);
  lut lut_gate374(0x6, 1712, 1623, 1754);
  lut lut_gate375(0x3ac3, 1592, 1560, 1754, 1713, 1755);
  lut lut_gate376(0x3caa, 1702, 1735, 1575, 1736, 1756);
  lut lut_gate377(0x96, 1737, 1734, 1727, 1757);
  lut lut_gate378(0x1ee1, 1757, 1756, 1702, 1578, N11342);
  lut lut_gate379(0x6996, N153, N154, N155, N156, 1758);
  lut lut_gate380(0xbf40, 1450, 1758, N18, 1448, 1759);
  lut lut_gate381(0x96ff, 1740, 1451, 1449, 1759, N10574);
  lut lut_gate382(0x3caa, N18, N198, N208, N44, 1760);
  lut lut_gate383(0x96, 1554, 1549, 1760, 1761);
  lut lut_gate384(0x06f0, N18, 1448, 1745, N176, 1762);
  lut lut_gate385(0x4100, 1742, 1744, 1762, 1536, 1763);
  lut lut_gate386(0xb4ff, 1763, 1761, N41, N18, N10576);
  lut lut_gate387(0x7100, 1654, 1555, 1746, 1509, 1764);
  lut lut_gate388(0x6f, 1764, 1557, 1511, 1765);
  lut lut_gate389(0x4, 1663, 1655, 1766);
  lut lut_gate390(0x4, 1528, 1766, 1546, 1529, 1767);
  lut lut_gate391(0x5c, 1767, 1528, 1545, 1768);
  lut lut_gate392(0x4b3c, 1710, 1608, 1614, 1605, 1769);
  lut lut_gate393(0xe73c, 1753, 1612, N299, 1615, 1770);
  lut lut_gate394(0x6996, 1755, 1711, 1617, 1606, 1771);
  lut lut_gate395(0x5ac3, 1753, 1771, 1769, 1610, 1772);
  lut lut_gate396(0x6, 1772, 1770, N11333);
  lut lut_gate397(0x70, 1562, 1567, 1642, 1773);
  lut lut_gate398(0x0, 1590, 1773, 1587, 1774);
  lut lut_gate399(0x3ca3, 1642, 1569, 1723, 1725, 1775);
  lut lut_gate400(0x6996, 1775, 1722, 1707, 1588, 1776);
  lut lut_gate401(0x2b4, 1774, 1776, 1480, N361, 1777);
  lut lut_gate402(0x18, 1478, 1773, N355, 1778);
  lut lut_gate403(0x6, 1778, 1777, N11340);

endmodule
