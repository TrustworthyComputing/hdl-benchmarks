module c2670(G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, G1014, G1017, G1021, G1026, G1030, G1033, G1036, G1148, G1152, G1159, G1193, G1231, G1237, G1240, G1329, G1336, G1342, G1345, G1348, G1351, G1377, G1478, G1540, G1546, G1563, G1578, G1584, G1650, G1653, G1661, G1663, G1675, G1682, G1683, G1720, G1721, G1722, G1723, G1724, G1725, G1726, G1727, G1734, G1735, G1946, G2418, G2488, G2512, G2515, G2516, G2517, G2520, G2523, G2524, G291, G292, G598, G603, G614, G631, G636, G647, G663, G674, G701, G703, G704, G705, G706, G707, G718, G734, G739, G745, G747, G748, G749, G750, G751, G756, G761, G766, G771, G772, G773, G774, G775, G776, G780, G783, G786, G789, G792, G795, G798, G801, G804, G807, G810, G811, G812, G815, G818, G821, G824, G827;
  input G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594;
  lut lut_gate1(0x6, 0620, 0615, G2583);
  lut lut_gate2(0x6, 0619, 0616, 0615);
  lut lut_gate3(0x9, 0618, 0617, 0616);
  lut lut_gate4(0x6, G131, G132, 0617);
  lut lut_gate5(0x9, G156, G128, 0618);
  lut lut_gate6(0x6, G129, G130, 0619);
  lut lut_gate7(0x9, 0622, 0621, 0620);
  lut lut_gate8(0x9, G133, G134, 0621);
  lut lut_gate9(0x9, G135, G136, 0622);
  lut lut_gate10(0x9, 0626, 0623, G2582);
  lut lut_gate11(0x9, 0625, 0624, 0623);
  lut lut_gate12(0x6, G139, G140, 0624);
  lut lut_gate13(0x6, G141, G142, 0625);
  lut lut_gate14(0x6, 0628, 0627, 0626);
  lut lut_gate15(0x9, G143, G144, 0627);
  lut lut_gate16(0x6, G157, G138, 0628);
  lut lut_gate17(0x9, 0716, 0713, 0629);
  lut lut_gate18(0x9, 0722, 0719, 0630);
  lut lut_gate19(0x6, 0725, 0632, 0631);
  lut lut_gate20(0x6, G2558, G2557, 0632);
  lut lut_gate21(0x6, 0637, 0634, 0633);
  lut lut_gate22(0x6, 0636, 0635, 0634);
  lut lut_gate23(0x9, 0738, 0735, 0635);
  lut lut_gate24(0x9, G2561, G2562, 0636);
  lut lut_gate25(0x9, 0741, G2566, 0637);
  lut lut_gate26(0x9, 0640, 0639, 0638);
  lut lut_gate27(0x6, G2571, G2570, 0639);
  lut lut_gate28(0x9, G2560, G2572, 0640);
  lut lut_gate29(0x8, 0643, 0642, 0641);
  lut lut_gate30(0x1, G127, G2559, 0642);
  lut lut_gate31(0x8, G30, G2557, 0643);
  lut lut_gate32(0x8, G2571, G2570, 0644);
  lut lut_gate33(0x8, G132, G133, 0645);
  lut lut_gate34(0x4, 0643, 0642, 0646);
  lut lut_gate35(0x7, 0648, 0647, G2547);
  lut lut_gate36(0x8, G139, G140, 0647);
  lut lut_gate37(0x8, G141, G142, 0648);
  lut lut_gate38(0x7, G121, 0649, G2548);
  lut lut_gate39(0x8, G2, G11, 0649);
  lut lut_gate40(0x7, G7, G121, G2551);
  lut lut_gate41(0xb, G119, G2551, G2552);
  lut lut_gate42(0xb, G147, G2551, G2553);
  lut lut_gate43(0x7, 0653, 0650, G2554);
  lut lut_gate44(0x8, 0652, 0651, 0650);
  lut lut_gate45(0x8, G106, G32, 0651);
  lut lut_gate46(0x8, G76, G64, 0652);
  lut lut_gate47(0x8, 0655, 0654, 0653);
  lut lut_gate48(0x8, G96, G53, 0654);
  lut lut_gate49(0x8, G86, G43, 0655);
  lut lut_gate50(0xe, 0657, 0656, G2556);
  lut lut_gate51(0x4, G147, 0650, 0656);
  lut lut_gate52(0x4, G119, 0653, 0657);
  lut lut_gate53(0x7, G28, 0658, G2564);
  lut lut_gate54(0x4, 0659, G2556, 0658);
  lut lut_gate55(0x4, G116, G121, 0659);
  lut lut_gate56(0xb, 0658, 0660, G2565);
  lut lut_gate57(0x8, G1, G3, 0660);
  lut lut_gate58(0xe, G144, 0661, G2580);
  lut lut_gate59(0x6, G143, 0725, 0661);
  lut lut_gate60(0x6, 0666, 0663, 0662);
  lut lut_gate61(0x6, 0665, 0664, 0663);
  lut lut_gate62(0x6, G152, G153, 0664);
  lut lut_gate63(0x9, G148, G149, 0665);
  lut lut_gate64(0x6, G150, G151, 0666);
  lut lut_gate65(0x9, 0669, 0668, 0667);
  lut lut_gate66(0x6, G154, G155, 0668);
  lut lut_gate67(0x9, G125, G126, 0669);
  lut lut_gate68(0x4, G142, 0762, 0670);
  lut lut_gate69(0x1, G134, 0768, 0671);
  lut lut_gate70(0x1, 0674, 0673, 0672);
  lut lut_gate71(0x1, G130, 0769, 0673);
  lut lut_gate72(0x1, G128, 0770, 0674);
  lut lut_gate73(0x4, G141, 0771, 0675);
  lut lut_gate74(0x1, 0678, 0677, 0676);
  lut lut_gate75(0x4, 0771, G141, 0677);
  lut lut_gate76(0x8, G130, 0769, 0678);
  lut lut_gate77(0x4, 0680, 0683, 0679);
  lut lut_gate78(0x1, 0682, 0681, 0680);
  lut lut_gate79(0x4, 0762, G142, 0681);
  lut lut_gate80(0x8, G128, 0770, 0682);
  lut lut_gate81(0x8, G134, 0768, 0683);
  lut lut_gate82(0x9, 0638, 0685, 0684);
  lut lut_gate83(0x9, G2566, 0686, 0685);
  lut lut_gate84(0x6, 0687, 0635, 0686);
  lut lut_gate85(0x8, G118, 0741, 0687);
  lut lut_gate86(0x7, G2590, 0688, G2593);
  lut lut_gate87(0x8, 0689, G2587, 0688);
  lut lut_gate88(0x8, 0690, G2581, 0689);
  lut lut_gate89(0x4, 0691, G2583, 0690);
  lut lut_gate90(0x1, G2582, G2556, 0691);
  lut lut_gate91(0x4, G74, G115, G2550);
  lut lut_gate92(0x7, G122, 0735, G2563);
  lut lut_gate93(0xb, 0741, 0692, G2577);
  lut lut_gate94(0x4, G118, G122, 0692);
  lut lut_gate95(0x1, G2562, G2567);
  lut lut_gate96(0x1, G115, G2531);
  lut lut_gate97(0x1, G124, G2534);
  lut lut_gate98(0x1, G137, G2536);
  lut lut_gate99(0x1, G32, G2539);
  lut lut_gate100(0x1, G106, G2540);
  lut lut_gate101(0x1, G64, G2541);
  lut lut_gate102(0x1, G76, G2542);
  lut lut_gate103(0x1, G53, G2543);
  lut lut_gate104(0x1, G96, G2544);
  lut lut_gate105(0x1, G43, G2545);
  lut lut_gate106(0x1, G86, G2546);
  lut lut_gate107(0x1, G2560, G2569);
  lut lut_gate108(0x1, G2561, G2568);
  lut lut_gate109(0xca, G120, G71, G49, 0693);
  lut lut_gate110(0xca, G120, G39, G60, 0694);
  lut lut_gate111(0xca, G117, 0693, 0694, G2566);
  lut lut_gate112(0xbc, G120, G117, G67, 0695);
  lut lut_gate113(0xc5, G120, G35, G56, 0696);
  lut lut_gate114(0xe1, 0695, 0696, G117, G2570);
  lut lut_gate115(0xca, G120, G66, G45, 0697);
  lut lut_gate116(0xca, G120, G34, G55, 0698);
  lut lut_gate117(0xca, G117, 0697, 0698, G2571);
  lut lut_gate118(0xca, G120, G65, G44, 0699);
  lut lut_gate119(0xca, G120, G33, G54, 0700);
  lut lut_gate120(0xca, G117, 0699, 0700, G2572);
  lut lut_gate121(0xca, G145, G109, G79, 0701);
  lut lut_gate122(0x3a, G146, 0701, 0702, G2557);
  lut lut_gate123(0x35, G145, G99, G89, 0702);
  lut lut_gate124(0xca, G145, G108, G78, 0703);
  lut lut_gate125(0x3a, G146, 0703, 0704, G2558);
  lut lut_gate126(0x35, G145, G98, G88, 0704);
  lut lut_gate127(0xca, G145, G110, G80, 0705);
  lut lut_gate128(0x3a, G146, 0705, 0706, G2559);
  lut lut_gate129(0x35, G145, G100, G90, 0706);
  lut lut_gate130(0xbe, 0631, 0711, G29, G2587);
  lut lut_gate131(0xca, G146, G114, G104, 0707);
  lut lut_gate132(0xca, G146, G84, G94, 0708);
  lut lut_gate133(0xca, G145, 0707, 0708, 0709);
  lut lut_gate134(0x96, G2559, 0630, 0629, 0710);
  lut lut_gate135(0x6, 0710, 0709, 0711);
  lut lut_gate136(0xca, G145, G112, G82, 0712);
  lut lut_gate137(0x3a, G146, 0712, 0714, 0713);
  lut lut_gate138(0x35, G145, G102, G92, 0714);
  lut lut_gate139(0xca, G145, G113, G83, 0715);
  lut lut_gate140(0x3a, G146, 0715, 0717, 0716);
  lut lut_gate141(0x35, G145, G103, G93, 0717);
  lut lut_gate142(0xca, G145, G105, G75, 0718);
  lut lut_gate143(0xca, G146, 0718, 0720, 0719);
  lut lut_gate144(0xca, G145, G95, G85, 0720);
  lut lut_gate145(0xca, G145, G111, G81, 0721);
  lut lut_gate146(0x3a, G146, 0721, 0723, 0722);
  lut lut_gate147(0x35, G145, G101, G91, 0723);
  lut lut_gate148(0xca, G145, G107, G77, 0724);
  lut lut_gate149(0x3a, G146, 0724, 0726, 0725);
  lut lut_gate150(0x35, G145, G97, G87, 0726);
  lut lut_gate151(0xca, G120, G68, G46, 0727);
  lut lut_gate152(0xca, G120, G36, G57, 0728);
  lut lut_gate153(0x35, G117, 0727, 0728, G2560);
  lut lut_gate154(0xca, G120, G70, G48, 0729);
  lut lut_gate155(0xca, G120, G38, G59, 0730);
  lut lut_gate156(0x35, G117, 0729, 0730, G2562);
  lut lut_gate157(0xca, G120, G69, G47, 0731);
  lut lut_gate158(0xca, G120, G37, G58, 0732);
  lut lut_gate159(0x35, G117, 0731, 0732, G2561);
  lut lut_gate160(0xbe, 0638, 0633, G29, G2590);
  lut lut_gate161(0xca, G120, G63, G42, 0733);
  lut lut_gate162(0xca, G120, G31, G52, 0734);
  lut lut_gate163(0x35, G117, 0733, 0734, 0735);
  lut lut_gate164(0xca, G120, G73, G51, 0736);
  lut lut_gate165(0xca, G120, G41, G62, 0737);
  lut lut_gate166(0x35, G117, 0736, 0737, 0738);
  lut lut_gate167(0xca, G120, G72, G50, 0739);
  lut lut_gate168(0xca, G120, G40, G61, 0740);
  lut lut_gate169(0x35, G117, 0739, 0740, 0741);
  lut lut_gate170(0xe8, G2566, 0746, 0789, 0742);
  lut lut_gate171(0x35, 0641, G138, G126, 0743);
  lut lut_gate172(0x35, 0641, G136, G125, 0744);
  lut lut_gate173(0x8, 0735, 0744, 0745);
  lut lut_gate174(0x53, 0641, G128, G139, 0746);
  lut lut_gate175(0x53, 0641, G129, G140, 0747);
  lut lut_gate176(0xac, 0641, G130, G141, 0748);
  lut lut_gate177(0x3a, G123, G2562, 0741, G2573);
  lut lut_gate178(0xca, G123, G2561, G2566, G2575);
  lut lut_gate179(0x4, 0741, G118, 0749);
  lut lut_gate180(0xca, G123, 0749, 0735, G2578);
  lut lut_gate181(0x6f, G10, 0667, 0662, G2581);
  lut lut_gate182(0x90, 0676, 0775, G135, 0750);
  lut lut_gate183(0x60, 0777, 0774, G129, 0751);
  lut lut_gate184(0x80, 0679, 0751, 0750, 0752);
  lut lut_gate185(0xb4, G138, G23, G20, 0753);
  lut lut_gate186(0xb4, 0753, 0713, G23, 0754);
  lut lut_gate187(0xb4, G139, G23, G25, 0755);
  lut lut_gate188(0xb4, 0755, 0722, G23, 0756);
  lut lut_gate189(0x8, 0766, 0759, 0757);
  lut lut_gate190(0xca, G12, G17, G2570, 0758);
  lut lut_gate191(0x90, 0761, 0758, G132, 0759);
  lut lut_gate192(0xc5, G23, G22, 0725, 0760);
  lut lut_gate193(0x40, 0760, G9, 0670, 0761);
  lut lut_gate194(0xc5, G23, G27, G2558, 0762);
  lut lut_gate195(0x14, 0767, G131, 0671, 0763);
  lut lut_gate196(0xc5, G12, G4, 0741, 0764);
  lut lut_gate197(0x41, G126, 0764, 0675, 0765);
  lut lut_gate198(0x80, 0672, 0765, 0763, 0766);
  lut lut_gate199(0x3a, G12, G16, G2560, 0767);
  lut lut_gate200(0x35, G12, G18, G2572, 0768);
  lut lut_gate201(0x3a, G12, G15, G2561, 0769);
  lut lut_gate202(0x35, G12, G14, G2566, 0770);
  lut lut_gate203(0xc5, G23, G26, G2557, 0771);
  lut lut_gate204(0xca, G12, G6, G2571, 0772);
  lut lut_gate205(0x6, 0772, G133, 0773);
  lut lut_gate206(0x3a, G12, G5, G2562, 0774);
  lut lut_gate207(0xca, G23, G19, 0719, 0775);
  lut lut_gate208(0xc5, G12, G13, 0735, 0776);
  lut lut_gate209(0x9, 0776, G125, 0777);
  lut lut_gate210(0xc5, G123, 0684, 0738, G2588);
  lut lut_gate211(0x35, G122, 0738, 0686, G2586);
  lut lut_gate212(0x71, G2572, 0788, G134, 0778);
  lut lut_gate213(0xca, 0646, 0778, 0788, 0779);
  lut lut_gate214(0xb2, 0719, 0779, G135, 0780);
  lut lut_gate215(0x71, 0716, 0780, G136, 0781);
  lut lut_gate216(0xb2, 0713, 0781, G138, 0782);
  lut lut_gate217(0xca, 0646, 0782, 0779, G2591);
  lut lut_gate218(0x17, 0748, G2561, 0795, 0783);
  lut lut_gate219(0xac, 0641, G131, G142, 0784);
  lut lut_gate220(0xca, 0641, 0644, 0645, 0785);
  lut lut_gate221(0xb2, 0784, 0783, G2560, 0786);
  lut lut_gate222(0xac, 0785, 0641, 0786, 0787);
  lut lut_gate223(0xca, G8, 0787, 0795, 0788);
  lut lut_gate224(0xe8, 0745, 0743, 0741, 0789);
  lut lut_gate225(0xc5, G23, G24, 0716, 0790);
  lut lut_gate226(0x90, 0754, 0790, G136, 0791);
  lut lut_gate227(0x7f, 0794, 0752, 0791, G2584);
  lut lut_gate228(0xc5, G23, G21, G2559, 0792);
  lut lut_gate229(0x90, 0756, 0792, G140, 0793);
  lut lut_gate230(0x40, 0793, 0757, 0773, 0794);
  lut lut_gate231(0x2b, 0747, 0742, G2562, 0795);

endmodule
