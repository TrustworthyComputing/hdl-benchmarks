module mmult (a_0_0, b_0_0, a_0_1, b_0_1, a_0_2, b_0_2, a_0_3, b_0_3, a_0_4, b_0_4, a_0_5, b_0_5, a_0_6, b_0_6, a_0_7, b_0_7, a_0_8, b_0_8, a_0_9, b_0_9, a_1_0, b_1_0, a_1_1, b_1_1, a_1_2, b_1_2, a_1_3, b_1_3, a_1_4, b_1_4, a_1_5, b_1_5, a_1_6, b_1_6, a_1_7, b_1_7, a_1_8, b_1_8, a_1_9, b_1_9, a_2_0, b_2_0, a_2_1, b_2_1, a_2_2, b_2_2, a_2_3, b_2_3, a_2_4, b_2_4, a_2_5, b_2_5, a_2_6, b_2_6, a_2_7, b_2_7, a_2_8, b_2_8, a_2_9, b_2_9, a_3_0, b_3_0, a_3_1, b_3_1, a_3_2, b_3_2, a_3_3, b_3_3, a_3_4, b_3_4, a_3_5, b_3_5, a_3_6, b_3_6, a_3_7, b_3_7, a_3_8, b_3_8, a_3_9, b_3_9, a_4_0, b_4_0, a_4_1, b_4_1, a_4_2, b_4_2, a_4_3, b_4_3, a_4_4, b_4_4, a_4_5, b_4_5, a_4_6, b_4_6, a_4_7, b_4_7, a_4_8, b_4_8, a_4_9, b_4_9, a_5_0, b_5_0, a_5_1, b_5_1, a_5_2, b_5_2, a_5_3, b_5_3, a_5_4, b_5_4, a_5_5, b_5_5, a_5_6, b_5_6, a_5_7, b_5_7, a_5_8, b_5_8, a_5_9, b_5_9, a_6_0, b_6_0, a_6_1, b_6_1, a_6_2, b_6_2, a_6_3, b_6_3, a_6_4, b_6_4, a_6_5, b_6_5, a_6_6, b_6_6, a_6_7, b_6_7, a_6_8, b_6_8, a_6_9, b_6_9, a_7_0, b_7_0, a_7_1, b_7_1, a_7_2, b_7_2, a_7_3, b_7_3, a_7_4, b_7_4, a_7_5, b_7_5, a_7_6, b_7_6, a_7_7, b_7_7, a_7_8, b_7_8, a_7_9, b_7_9, a_8_0, b_8_0, a_8_1, b_8_1, a_8_2, b_8_2, a_8_3, b_8_3, a_8_4, b_8_4, a_8_5, b_8_5, a_8_6, b_8_6, a_8_7, b_8_7, a_8_8, b_8_8, a_8_9, b_8_9, a_9_0, b_9_0, a_9_1, b_9_1, a_9_2, b_9_2, a_9_3, b_9_3, a_9_4, b_9_4, a_9_5, b_9_5, a_9_6, b_9_6, a_9_7, b_9_7, a_9_8, b_9_8, a_9_9, b_9_9, c_0_0, c_0_1, c_0_2, c_0_3, c_0_4, c_0_5, c_0_6, c_0_7, c_0_8, c_0_9, c_1_0, c_1_1, c_1_2, c_1_3, c_1_4, c_1_5, c_1_6, c_1_7, c_1_8, c_1_9, c_2_0, c_2_1, c_2_2, c_2_3, c_2_4, c_2_5, c_2_6, c_2_7, c_2_8, c_2_9, c_3_0, c_3_1, c_3_2, c_3_3, c_3_4, c_3_5, c_3_6, c_3_7, c_3_8, c_3_9, c_4_0, c_4_1, c_4_2, c_4_3, c_4_4, c_4_5, c_4_6, c_4_7, c_4_8, c_4_9, c_5_0, c_5_1, c_5_2, c_5_3, c_5_4, c_5_5, c_5_6, c_5_7, c_5_8, c_5_9, c_6_0, c_6_1, c_6_2, c_6_3, c_6_4, c_6_5, c_6_6, c_6_7, c_6_8, c_6_9, c_7_0, c_7_1, c_7_2, c_7_3, c_7_4, c_7_5, c_7_6, c_7_7, c_7_8, c_7_9, c_8_0, c_8_1, c_8_2, c_8_3, c_8_4, c_8_5, c_8_6, c_8_7, c_8_8, c_8_9, c_9_0, c_9_1, c_9_2, c_9_3, c_9_4, c_9_5, c_9_6, c_9_7, c_9_8, c_9_9);

  input [15:0] a_0_0;
  input [15:0] b_0_0;
  input [15:0] a_0_1;
  input [15:0] b_0_1;
  input [15:0] a_0_2;
  input [15:0] b_0_2;
  input [15:0] a_0_3;
  input [15:0] b_0_3;
  input [15:0] a_0_4;
  input [15:0] b_0_4;
  input [15:0] a_0_5;
  input [15:0] b_0_5;
  input [15:0] a_0_6;
  input [15:0] b_0_6;
  input [15:0] a_0_7;
  input [15:0] b_0_7;
  input [15:0] a_0_8;
  input [15:0] b_0_8;
  input [15:0] a_0_9;
  input [15:0] b_0_9;
  input [15:0] a_1_0;
  input [15:0] b_1_0;
  input [15:0] a_1_1;
  input [15:0] b_1_1;
  input [15:0] a_1_2;
  input [15:0] b_1_2;
  input [15:0] a_1_3;
  input [15:0] b_1_3;
  input [15:0] a_1_4;
  input [15:0] b_1_4;
  input [15:0] a_1_5;
  input [15:0] b_1_5;
  input [15:0] a_1_6;
  input [15:0] b_1_6;
  input [15:0] a_1_7;
  input [15:0] b_1_7;
  input [15:0] a_1_8;
  input [15:0] b_1_8;
  input [15:0] a_1_9;
  input [15:0] b_1_9;
  input [15:0] a_2_0;
  input [15:0] b_2_0;
  input [15:0] a_2_1;
  input [15:0] b_2_1;
  input [15:0] a_2_2;
  input [15:0] b_2_2;
  input [15:0] a_2_3;
  input [15:0] b_2_3;
  input [15:0] a_2_4;
  input [15:0] b_2_4;
  input [15:0] a_2_5;
  input [15:0] b_2_5;
  input [15:0] a_2_6;
  input [15:0] b_2_6;
  input [15:0] a_2_7;
  input [15:0] b_2_7;
  input [15:0] a_2_8;
  input [15:0] b_2_8;
  input [15:0] a_2_9;
  input [15:0] b_2_9;
  input [15:0] a_3_0;
  input [15:0] b_3_0;
  input [15:0] a_3_1;
  input [15:0] b_3_1;
  input [15:0] a_3_2;
  input [15:0] b_3_2;
  input [15:0] a_3_3;
  input [15:0] b_3_3;
  input [15:0] a_3_4;
  input [15:0] b_3_4;
  input [15:0] a_3_5;
  input [15:0] b_3_5;
  input [15:0] a_3_6;
  input [15:0] b_3_6;
  input [15:0] a_3_7;
  input [15:0] b_3_7;
  input [15:0] a_3_8;
  input [15:0] b_3_8;
  input [15:0] a_3_9;
  input [15:0] b_3_9;
  input [15:0] a_4_0;
  input [15:0] b_4_0;
  input [15:0] a_4_1;
  input [15:0] b_4_1;
  input [15:0] a_4_2;
  input [15:0] b_4_2;
  input [15:0] a_4_3;
  input [15:0] b_4_3;
  input [15:0] a_4_4;
  input [15:0] b_4_4;
  input [15:0] a_4_5;
  input [15:0] b_4_5;
  input [15:0] a_4_6;
  input [15:0] b_4_6;
  input [15:0] a_4_7;
  input [15:0] b_4_7;
  input [15:0] a_4_8;
  input [15:0] b_4_8;
  input [15:0] a_4_9;
  input [15:0] b_4_9;
  input [15:0] a_5_0;
  input [15:0] b_5_0;
  input [15:0] a_5_1;
  input [15:0] b_5_1;
  input [15:0] a_5_2;
  input [15:0] b_5_2;
  input [15:0] a_5_3;
  input [15:0] b_5_3;
  input [15:0] a_5_4;
  input [15:0] b_5_4;
  input [15:0] a_5_5;
  input [15:0] b_5_5;
  input [15:0] a_5_6;
  input [15:0] b_5_6;
  input [15:0] a_5_7;
  input [15:0] b_5_7;
  input [15:0] a_5_8;
  input [15:0] b_5_8;
  input [15:0] a_5_9;
  input [15:0] b_5_9;
  input [15:0] a_6_0;
  input [15:0] b_6_0;
  input [15:0] a_6_1;
  input [15:0] b_6_1;
  input [15:0] a_6_2;
  input [15:0] b_6_2;
  input [15:0] a_6_3;
  input [15:0] b_6_3;
  input [15:0] a_6_4;
  input [15:0] b_6_4;
  input [15:0] a_6_5;
  input [15:0] b_6_5;
  input [15:0] a_6_6;
  input [15:0] b_6_6;
  input [15:0] a_6_7;
  input [15:0] b_6_7;
  input [15:0] a_6_8;
  input [15:0] b_6_8;
  input [15:0] a_6_9;
  input [15:0] b_6_9;
  input [15:0] a_7_0;
  input [15:0] b_7_0;
  input [15:0] a_7_1;
  input [15:0] b_7_1;
  input [15:0] a_7_2;
  input [15:0] b_7_2;
  input [15:0] a_7_3;
  input [15:0] b_7_3;
  input [15:0] a_7_4;
  input [15:0] b_7_4;
  input [15:0] a_7_5;
  input [15:0] b_7_5;
  input [15:0] a_7_6;
  input [15:0] b_7_6;
  input [15:0] a_7_7;
  input [15:0] b_7_7;
  input [15:0] a_7_8;
  input [15:0] b_7_8;
  input [15:0] a_7_9;
  input [15:0] b_7_9;
  input [15:0] a_8_0;
  input [15:0] b_8_0;
  input [15:0] a_8_1;
  input [15:0] b_8_1;
  input [15:0] a_8_2;
  input [15:0] b_8_2;
  input [15:0] a_8_3;
  input [15:0] b_8_3;
  input [15:0] a_8_4;
  input [15:0] b_8_4;
  input [15:0] a_8_5;
  input [15:0] b_8_5;
  input [15:0] a_8_6;
  input [15:0] b_8_6;
  input [15:0] a_8_7;
  input [15:0] b_8_7;
  input [15:0] a_8_8;
  input [15:0] b_8_8;
  input [15:0] a_8_9;
  input [15:0] b_8_9;
  input [15:0] a_9_0;
  input [15:0] b_9_0;
  input [15:0] a_9_1;
  input [15:0] b_9_1;
  input [15:0] a_9_2;
  input [15:0] b_9_2;
  input [15:0] a_9_3;
  input [15:0] b_9_3;
  input [15:0] a_9_4;
  input [15:0] b_9_4;
  input [15:0] a_9_5;
  input [15:0] b_9_5;
  input [15:0] a_9_6;
  input [15:0] b_9_6;
  input [15:0] a_9_7;
  input [15:0] b_9_7;
  input [15:0] a_9_8;
  input [15:0] b_9_8;
  input [15:0] a_9_9;
  input [15:0] b_9_9;

  output [15:0] c_0_0;
  output [15:0] c_0_1;
  output [15:0] c_0_2;
  output [15:0] c_0_3;
  output [15:0] c_0_4;
  output [15:0] c_0_5;
  output [15:0] c_0_6;
  output [15:0] c_0_7;
  output [15:0] c_0_8;
  output [15:0] c_0_9;
  output [15:0] c_1_0;
  output [15:0] c_1_1;
  output [15:0] c_1_2;
  output [15:0] c_1_3;
  output [15:0] c_1_4;
  output [15:0] c_1_5;
  output [15:0] c_1_6;
  output [15:0] c_1_7;
  output [15:0] c_1_8;
  output [15:0] c_1_9;
  output [15:0] c_2_0;
  output [15:0] c_2_1;
  output [15:0] c_2_2;
  output [15:0] c_2_3;
  output [15:0] c_2_4;
  output [15:0] c_2_5;
  output [15:0] c_2_6;
  output [15:0] c_2_7;
  output [15:0] c_2_8;
  output [15:0] c_2_9;
  output [15:0] c_3_0;
  output [15:0] c_3_1;
  output [15:0] c_3_2;
  output [15:0] c_3_3;
  output [15:0] c_3_4;
  output [15:0] c_3_5;
  output [15:0] c_3_6;
  output [15:0] c_3_7;
  output [15:0] c_3_8;
  output [15:0] c_3_9;
  output [15:0] c_4_0;
  output [15:0] c_4_1;
  output [15:0] c_4_2;
  output [15:0] c_4_3;
  output [15:0] c_4_4;
  output [15:0] c_4_5;
  output [15:0] c_4_6;
  output [15:0] c_4_7;
  output [15:0] c_4_8;
  output [15:0] c_4_9;
  output [15:0] c_5_0;
  output [15:0] c_5_1;
  output [15:0] c_5_2;
  output [15:0] c_5_3;
  output [15:0] c_5_4;
  output [15:0] c_5_5;
  output [15:0] c_5_6;
  output [15:0] c_5_7;
  output [15:0] c_5_8;
  output [15:0] c_5_9;
  output [15:0] c_6_0;
  output [15:0] c_6_1;
  output [15:0] c_6_2;
  output [15:0] c_6_3;
  output [15:0] c_6_4;
  output [15:0] c_6_5;
  output [15:0] c_6_6;
  output [15:0] c_6_7;
  output [15:0] c_6_8;
  output [15:0] c_6_9;
  output [15:0] c_7_0;
  output [15:0] c_7_1;
  output [15:0] c_7_2;
  output [15:0] c_7_3;
  output [15:0] c_7_4;
  output [15:0] c_7_5;
  output [15:0] c_7_6;
  output [15:0] c_7_7;
  output [15:0] c_7_8;
  output [15:0] c_7_9;
  output [15:0] c_8_0;
  output [15:0] c_8_1;
  output [15:0] c_8_2;
  output [15:0] c_8_3;
  output [15:0] c_8_4;
  output [15:0] c_8_5;
  output [15:0] c_8_6;
  output [15:0] c_8_7;
  output [15:0] c_8_8;
  output [15:0] c_8_9;
  output [15:0] c_9_0;
  output [15:0] c_9_1;
  output [15:0] c_9_2;
  output [15:0] c_9_3;
  output [15:0] c_9_4;
  output [15:0] c_9_5;
  output [15:0] c_9_6;
  output [15:0] c_9_7;
  output [15:0] c_9_8;
  output [15:0] c_9_9;

  wire [15:0] t0_r0_c0_rr0;
  wire [15:0] t0_r0_c0_rr1;
  wire [15:0] t0_r0_c0_rr2;
  wire [15:0] t0_r0_c0_rr3;
  wire [15:0] t0_r0_c0_rr4;
  wire [15:0] t0_r0_c0_rr5;
  wire [15:0] t0_r0_c0_rr6;
  wire [15:0] t0_r0_c0_rr7;
  wire [15:0] t0_r0_c0_rr8;
  wire [15:0] t0_r0_c0_rr9;
  wire [15:0] t1_r0_c0_rr0;
  wire [15:0] t1_r0_c0_rr1;
  wire [15:0] t1_r0_c0_rr2;
  wire [15:0] t1_r0_c0_rr3;
  wire [15:0] t1_r0_c0_rr4;
  wire [15:0] t2_r0_c0_rr0;
  wire [15:0] t2_r0_c0_rr1;
  wire [15:0] t2_r0_c0_rr2;
  wire [15:0] t3_r0_c0_rr0;
  wire [15:0] t3_r0_c0_rr1;
  wire [15:0] t4_r0_c0_rr0;
  wire [15:0] t0_r0_c1_rr0;
  wire [15:0] t0_r0_c1_rr1;
  wire [15:0] t0_r0_c1_rr2;
  wire [15:0] t0_r0_c1_rr3;
  wire [15:0] t0_r0_c1_rr4;
  wire [15:0] t0_r0_c1_rr5;
  wire [15:0] t0_r0_c1_rr6;
  wire [15:0] t0_r0_c1_rr7;
  wire [15:0] t0_r0_c1_rr8;
  wire [15:0] t0_r0_c1_rr9;
  wire [15:0] t1_r0_c1_rr0;
  wire [15:0] t1_r0_c1_rr1;
  wire [15:0] t1_r0_c1_rr2;
  wire [15:0] t1_r0_c1_rr3;
  wire [15:0] t1_r0_c1_rr4;
  wire [15:0] t2_r0_c1_rr0;
  wire [15:0] t2_r0_c1_rr1;
  wire [15:0] t2_r0_c1_rr2;
  wire [15:0] t3_r0_c1_rr0;
  wire [15:0] t3_r0_c1_rr1;
  wire [15:0] t4_r0_c1_rr0;
  wire [15:0] t0_r0_c2_rr0;
  wire [15:0] t0_r0_c2_rr1;
  wire [15:0] t0_r0_c2_rr2;
  wire [15:0] t0_r0_c2_rr3;
  wire [15:0] t0_r0_c2_rr4;
  wire [15:0] t0_r0_c2_rr5;
  wire [15:0] t0_r0_c2_rr6;
  wire [15:0] t0_r0_c2_rr7;
  wire [15:0] t0_r0_c2_rr8;
  wire [15:0] t0_r0_c2_rr9;
  wire [15:0] t1_r0_c2_rr0;
  wire [15:0] t1_r0_c2_rr1;
  wire [15:0] t1_r0_c2_rr2;
  wire [15:0] t1_r0_c2_rr3;
  wire [15:0] t1_r0_c2_rr4;
  wire [15:0] t2_r0_c2_rr0;
  wire [15:0] t2_r0_c2_rr1;
  wire [15:0] t2_r0_c2_rr2;
  wire [15:0] t3_r0_c2_rr0;
  wire [15:0] t3_r0_c2_rr1;
  wire [15:0] t4_r0_c2_rr0;
  wire [15:0] t0_r0_c3_rr0;
  wire [15:0] t0_r0_c3_rr1;
  wire [15:0] t0_r0_c3_rr2;
  wire [15:0] t0_r0_c3_rr3;
  wire [15:0] t0_r0_c3_rr4;
  wire [15:0] t0_r0_c3_rr5;
  wire [15:0] t0_r0_c3_rr6;
  wire [15:0] t0_r0_c3_rr7;
  wire [15:0] t0_r0_c3_rr8;
  wire [15:0] t0_r0_c3_rr9;
  wire [15:0] t1_r0_c3_rr0;
  wire [15:0] t1_r0_c3_rr1;
  wire [15:0] t1_r0_c3_rr2;
  wire [15:0] t1_r0_c3_rr3;
  wire [15:0] t1_r0_c3_rr4;
  wire [15:0] t2_r0_c3_rr0;
  wire [15:0] t2_r0_c3_rr1;
  wire [15:0] t2_r0_c3_rr2;
  wire [15:0] t3_r0_c3_rr0;
  wire [15:0] t3_r0_c3_rr1;
  wire [15:0] t4_r0_c3_rr0;
  wire [15:0] t0_r0_c4_rr0;
  wire [15:0] t0_r0_c4_rr1;
  wire [15:0] t0_r0_c4_rr2;
  wire [15:0] t0_r0_c4_rr3;
  wire [15:0] t0_r0_c4_rr4;
  wire [15:0] t0_r0_c4_rr5;
  wire [15:0] t0_r0_c4_rr6;
  wire [15:0] t0_r0_c4_rr7;
  wire [15:0] t0_r0_c4_rr8;
  wire [15:0] t0_r0_c4_rr9;
  wire [15:0] t1_r0_c4_rr0;
  wire [15:0] t1_r0_c4_rr1;
  wire [15:0] t1_r0_c4_rr2;
  wire [15:0] t1_r0_c4_rr3;
  wire [15:0] t1_r0_c4_rr4;
  wire [15:0] t2_r0_c4_rr0;
  wire [15:0] t2_r0_c4_rr1;
  wire [15:0] t2_r0_c4_rr2;
  wire [15:0] t3_r0_c4_rr0;
  wire [15:0] t3_r0_c4_rr1;
  wire [15:0] t4_r0_c4_rr0;
  wire [15:0] t0_r0_c5_rr0;
  wire [15:0] t0_r0_c5_rr1;
  wire [15:0] t0_r0_c5_rr2;
  wire [15:0] t0_r0_c5_rr3;
  wire [15:0] t0_r0_c5_rr4;
  wire [15:0] t0_r0_c5_rr5;
  wire [15:0] t0_r0_c5_rr6;
  wire [15:0] t0_r0_c5_rr7;
  wire [15:0] t0_r0_c5_rr8;
  wire [15:0] t0_r0_c5_rr9;
  wire [15:0] t1_r0_c5_rr0;
  wire [15:0] t1_r0_c5_rr1;
  wire [15:0] t1_r0_c5_rr2;
  wire [15:0] t1_r0_c5_rr3;
  wire [15:0] t1_r0_c5_rr4;
  wire [15:0] t2_r0_c5_rr0;
  wire [15:0] t2_r0_c5_rr1;
  wire [15:0] t2_r0_c5_rr2;
  wire [15:0] t3_r0_c5_rr0;
  wire [15:0] t3_r0_c5_rr1;
  wire [15:0] t4_r0_c5_rr0;
  wire [15:0] t0_r0_c6_rr0;
  wire [15:0] t0_r0_c6_rr1;
  wire [15:0] t0_r0_c6_rr2;
  wire [15:0] t0_r0_c6_rr3;
  wire [15:0] t0_r0_c6_rr4;
  wire [15:0] t0_r0_c6_rr5;
  wire [15:0] t0_r0_c6_rr6;
  wire [15:0] t0_r0_c6_rr7;
  wire [15:0] t0_r0_c6_rr8;
  wire [15:0] t0_r0_c6_rr9;
  wire [15:0] t1_r0_c6_rr0;
  wire [15:0] t1_r0_c6_rr1;
  wire [15:0] t1_r0_c6_rr2;
  wire [15:0] t1_r0_c6_rr3;
  wire [15:0] t1_r0_c6_rr4;
  wire [15:0] t2_r0_c6_rr0;
  wire [15:0] t2_r0_c6_rr1;
  wire [15:0] t2_r0_c6_rr2;
  wire [15:0] t3_r0_c6_rr0;
  wire [15:0] t3_r0_c6_rr1;
  wire [15:0] t4_r0_c6_rr0;
  wire [15:0] t0_r0_c7_rr0;
  wire [15:0] t0_r0_c7_rr1;
  wire [15:0] t0_r0_c7_rr2;
  wire [15:0] t0_r0_c7_rr3;
  wire [15:0] t0_r0_c7_rr4;
  wire [15:0] t0_r0_c7_rr5;
  wire [15:0] t0_r0_c7_rr6;
  wire [15:0] t0_r0_c7_rr7;
  wire [15:0] t0_r0_c7_rr8;
  wire [15:0] t0_r0_c7_rr9;
  wire [15:0] t1_r0_c7_rr0;
  wire [15:0] t1_r0_c7_rr1;
  wire [15:0] t1_r0_c7_rr2;
  wire [15:0] t1_r0_c7_rr3;
  wire [15:0] t1_r0_c7_rr4;
  wire [15:0] t2_r0_c7_rr0;
  wire [15:0] t2_r0_c7_rr1;
  wire [15:0] t2_r0_c7_rr2;
  wire [15:0] t3_r0_c7_rr0;
  wire [15:0] t3_r0_c7_rr1;
  wire [15:0] t4_r0_c7_rr0;
  wire [15:0] t0_r0_c8_rr0;
  wire [15:0] t0_r0_c8_rr1;
  wire [15:0] t0_r0_c8_rr2;
  wire [15:0] t0_r0_c8_rr3;
  wire [15:0] t0_r0_c8_rr4;
  wire [15:0] t0_r0_c8_rr5;
  wire [15:0] t0_r0_c8_rr6;
  wire [15:0] t0_r0_c8_rr7;
  wire [15:0] t0_r0_c8_rr8;
  wire [15:0] t0_r0_c8_rr9;
  wire [15:0] t1_r0_c8_rr0;
  wire [15:0] t1_r0_c8_rr1;
  wire [15:0] t1_r0_c8_rr2;
  wire [15:0] t1_r0_c8_rr3;
  wire [15:0] t1_r0_c8_rr4;
  wire [15:0] t2_r0_c8_rr0;
  wire [15:0] t2_r0_c8_rr1;
  wire [15:0] t2_r0_c8_rr2;
  wire [15:0] t3_r0_c8_rr0;
  wire [15:0] t3_r0_c8_rr1;
  wire [15:0] t4_r0_c8_rr0;
  wire [15:0] t0_r0_c9_rr0;
  wire [15:0] t0_r0_c9_rr1;
  wire [15:0] t0_r0_c9_rr2;
  wire [15:0] t0_r0_c9_rr3;
  wire [15:0] t0_r0_c9_rr4;
  wire [15:0] t0_r0_c9_rr5;
  wire [15:0] t0_r0_c9_rr6;
  wire [15:0] t0_r0_c9_rr7;
  wire [15:0] t0_r0_c9_rr8;
  wire [15:0] t0_r0_c9_rr9;
  wire [15:0] t1_r0_c9_rr0;
  wire [15:0] t1_r0_c9_rr1;
  wire [15:0] t1_r0_c9_rr2;
  wire [15:0] t1_r0_c9_rr3;
  wire [15:0] t1_r0_c9_rr4;
  wire [15:0] t2_r0_c9_rr0;
  wire [15:0] t2_r0_c9_rr1;
  wire [15:0] t2_r0_c9_rr2;
  wire [15:0] t3_r0_c9_rr0;
  wire [15:0] t3_r0_c9_rr1;
  wire [15:0] t4_r0_c9_rr0;
  wire [15:0] t0_r1_c0_rr0;
  wire [15:0] t0_r1_c0_rr1;
  wire [15:0] t0_r1_c0_rr2;
  wire [15:0] t0_r1_c0_rr3;
  wire [15:0] t0_r1_c0_rr4;
  wire [15:0] t0_r1_c0_rr5;
  wire [15:0] t0_r1_c0_rr6;
  wire [15:0] t0_r1_c0_rr7;
  wire [15:0] t0_r1_c0_rr8;
  wire [15:0] t0_r1_c0_rr9;
  wire [15:0] t1_r1_c0_rr0;
  wire [15:0] t1_r1_c0_rr1;
  wire [15:0] t1_r1_c0_rr2;
  wire [15:0] t1_r1_c0_rr3;
  wire [15:0] t1_r1_c0_rr4;
  wire [15:0] t2_r1_c0_rr0;
  wire [15:0] t2_r1_c0_rr1;
  wire [15:0] t2_r1_c0_rr2;
  wire [15:0] t3_r1_c0_rr0;
  wire [15:0] t3_r1_c0_rr1;
  wire [15:0] t4_r1_c0_rr0;
  wire [15:0] t0_r1_c1_rr0;
  wire [15:0] t0_r1_c1_rr1;
  wire [15:0] t0_r1_c1_rr2;
  wire [15:0] t0_r1_c1_rr3;
  wire [15:0] t0_r1_c1_rr4;
  wire [15:0] t0_r1_c1_rr5;
  wire [15:0] t0_r1_c1_rr6;
  wire [15:0] t0_r1_c1_rr7;
  wire [15:0] t0_r1_c1_rr8;
  wire [15:0] t0_r1_c1_rr9;
  wire [15:0] t1_r1_c1_rr0;
  wire [15:0] t1_r1_c1_rr1;
  wire [15:0] t1_r1_c1_rr2;
  wire [15:0] t1_r1_c1_rr3;
  wire [15:0] t1_r1_c1_rr4;
  wire [15:0] t2_r1_c1_rr0;
  wire [15:0] t2_r1_c1_rr1;
  wire [15:0] t2_r1_c1_rr2;
  wire [15:0] t3_r1_c1_rr0;
  wire [15:0] t3_r1_c1_rr1;
  wire [15:0] t4_r1_c1_rr0;
  wire [15:0] t0_r1_c2_rr0;
  wire [15:0] t0_r1_c2_rr1;
  wire [15:0] t0_r1_c2_rr2;
  wire [15:0] t0_r1_c2_rr3;
  wire [15:0] t0_r1_c2_rr4;
  wire [15:0] t0_r1_c2_rr5;
  wire [15:0] t0_r1_c2_rr6;
  wire [15:0] t0_r1_c2_rr7;
  wire [15:0] t0_r1_c2_rr8;
  wire [15:0] t0_r1_c2_rr9;
  wire [15:0] t1_r1_c2_rr0;
  wire [15:0] t1_r1_c2_rr1;
  wire [15:0] t1_r1_c2_rr2;
  wire [15:0] t1_r1_c2_rr3;
  wire [15:0] t1_r1_c2_rr4;
  wire [15:0] t2_r1_c2_rr0;
  wire [15:0] t2_r1_c2_rr1;
  wire [15:0] t2_r1_c2_rr2;
  wire [15:0] t3_r1_c2_rr0;
  wire [15:0] t3_r1_c2_rr1;
  wire [15:0] t4_r1_c2_rr0;
  wire [15:0] t0_r1_c3_rr0;
  wire [15:0] t0_r1_c3_rr1;
  wire [15:0] t0_r1_c3_rr2;
  wire [15:0] t0_r1_c3_rr3;
  wire [15:0] t0_r1_c3_rr4;
  wire [15:0] t0_r1_c3_rr5;
  wire [15:0] t0_r1_c3_rr6;
  wire [15:0] t0_r1_c3_rr7;
  wire [15:0] t0_r1_c3_rr8;
  wire [15:0] t0_r1_c3_rr9;
  wire [15:0] t1_r1_c3_rr0;
  wire [15:0] t1_r1_c3_rr1;
  wire [15:0] t1_r1_c3_rr2;
  wire [15:0] t1_r1_c3_rr3;
  wire [15:0] t1_r1_c3_rr4;
  wire [15:0] t2_r1_c3_rr0;
  wire [15:0] t2_r1_c3_rr1;
  wire [15:0] t2_r1_c3_rr2;
  wire [15:0] t3_r1_c3_rr0;
  wire [15:0] t3_r1_c3_rr1;
  wire [15:0] t4_r1_c3_rr0;
  wire [15:0] t0_r1_c4_rr0;
  wire [15:0] t0_r1_c4_rr1;
  wire [15:0] t0_r1_c4_rr2;
  wire [15:0] t0_r1_c4_rr3;
  wire [15:0] t0_r1_c4_rr4;
  wire [15:0] t0_r1_c4_rr5;
  wire [15:0] t0_r1_c4_rr6;
  wire [15:0] t0_r1_c4_rr7;
  wire [15:0] t0_r1_c4_rr8;
  wire [15:0] t0_r1_c4_rr9;
  wire [15:0] t1_r1_c4_rr0;
  wire [15:0] t1_r1_c4_rr1;
  wire [15:0] t1_r1_c4_rr2;
  wire [15:0] t1_r1_c4_rr3;
  wire [15:0] t1_r1_c4_rr4;
  wire [15:0] t2_r1_c4_rr0;
  wire [15:0] t2_r1_c4_rr1;
  wire [15:0] t2_r1_c4_rr2;
  wire [15:0] t3_r1_c4_rr0;
  wire [15:0] t3_r1_c4_rr1;
  wire [15:0] t4_r1_c4_rr0;
  wire [15:0] t0_r1_c5_rr0;
  wire [15:0] t0_r1_c5_rr1;
  wire [15:0] t0_r1_c5_rr2;
  wire [15:0] t0_r1_c5_rr3;
  wire [15:0] t0_r1_c5_rr4;
  wire [15:0] t0_r1_c5_rr5;
  wire [15:0] t0_r1_c5_rr6;
  wire [15:0] t0_r1_c5_rr7;
  wire [15:0] t0_r1_c5_rr8;
  wire [15:0] t0_r1_c5_rr9;
  wire [15:0] t1_r1_c5_rr0;
  wire [15:0] t1_r1_c5_rr1;
  wire [15:0] t1_r1_c5_rr2;
  wire [15:0] t1_r1_c5_rr3;
  wire [15:0] t1_r1_c5_rr4;
  wire [15:0] t2_r1_c5_rr0;
  wire [15:0] t2_r1_c5_rr1;
  wire [15:0] t2_r1_c5_rr2;
  wire [15:0] t3_r1_c5_rr0;
  wire [15:0] t3_r1_c5_rr1;
  wire [15:0] t4_r1_c5_rr0;
  wire [15:0] t0_r1_c6_rr0;
  wire [15:0] t0_r1_c6_rr1;
  wire [15:0] t0_r1_c6_rr2;
  wire [15:0] t0_r1_c6_rr3;
  wire [15:0] t0_r1_c6_rr4;
  wire [15:0] t0_r1_c6_rr5;
  wire [15:0] t0_r1_c6_rr6;
  wire [15:0] t0_r1_c6_rr7;
  wire [15:0] t0_r1_c6_rr8;
  wire [15:0] t0_r1_c6_rr9;
  wire [15:0] t1_r1_c6_rr0;
  wire [15:0] t1_r1_c6_rr1;
  wire [15:0] t1_r1_c6_rr2;
  wire [15:0] t1_r1_c6_rr3;
  wire [15:0] t1_r1_c6_rr4;
  wire [15:0] t2_r1_c6_rr0;
  wire [15:0] t2_r1_c6_rr1;
  wire [15:0] t2_r1_c6_rr2;
  wire [15:0] t3_r1_c6_rr0;
  wire [15:0] t3_r1_c6_rr1;
  wire [15:0] t4_r1_c6_rr0;
  wire [15:0] t0_r1_c7_rr0;
  wire [15:0] t0_r1_c7_rr1;
  wire [15:0] t0_r1_c7_rr2;
  wire [15:0] t0_r1_c7_rr3;
  wire [15:0] t0_r1_c7_rr4;
  wire [15:0] t0_r1_c7_rr5;
  wire [15:0] t0_r1_c7_rr6;
  wire [15:0] t0_r1_c7_rr7;
  wire [15:0] t0_r1_c7_rr8;
  wire [15:0] t0_r1_c7_rr9;
  wire [15:0] t1_r1_c7_rr0;
  wire [15:0] t1_r1_c7_rr1;
  wire [15:0] t1_r1_c7_rr2;
  wire [15:0] t1_r1_c7_rr3;
  wire [15:0] t1_r1_c7_rr4;
  wire [15:0] t2_r1_c7_rr0;
  wire [15:0] t2_r1_c7_rr1;
  wire [15:0] t2_r1_c7_rr2;
  wire [15:0] t3_r1_c7_rr0;
  wire [15:0] t3_r1_c7_rr1;
  wire [15:0] t4_r1_c7_rr0;
  wire [15:0] t0_r1_c8_rr0;
  wire [15:0] t0_r1_c8_rr1;
  wire [15:0] t0_r1_c8_rr2;
  wire [15:0] t0_r1_c8_rr3;
  wire [15:0] t0_r1_c8_rr4;
  wire [15:0] t0_r1_c8_rr5;
  wire [15:0] t0_r1_c8_rr6;
  wire [15:0] t0_r1_c8_rr7;
  wire [15:0] t0_r1_c8_rr8;
  wire [15:0] t0_r1_c8_rr9;
  wire [15:0] t1_r1_c8_rr0;
  wire [15:0] t1_r1_c8_rr1;
  wire [15:0] t1_r1_c8_rr2;
  wire [15:0] t1_r1_c8_rr3;
  wire [15:0] t1_r1_c8_rr4;
  wire [15:0] t2_r1_c8_rr0;
  wire [15:0] t2_r1_c8_rr1;
  wire [15:0] t2_r1_c8_rr2;
  wire [15:0] t3_r1_c8_rr0;
  wire [15:0] t3_r1_c8_rr1;
  wire [15:0] t4_r1_c8_rr0;
  wire [15:0] t0_r1_c9_rr0;
  wire [15:0] t0_r1_c9_rr1;
  wire [15:0] t0_r1_c9_rr2;
  wire [15:0] t0_r1_c9_rr3;
  wire [15:0] t0_r1_c9_rr4;
  wire [15:0] t0_r1_c9_rr5;
  wire [15:0] t0_r1_c9_rr6;
  wire [15:0] t0_r1_c9_rr7;
  wire [15:0] t0_r1_c9_rr8;
  wire [15:0] t0_r1_c9_rr9;
  wire [15:0] t1_r1_c9_rr0;
  wire [15:0] t1_r1_c9_rr1;
  wire [15:0] t1_r1_c9_rr2;
  wire [15:0] t1_r1_c9_rr3;
  wire [15:0] t1_r1_c9_rr4;
  wire [15:0] t2_r1_c9_rr0;
  wire [15:0] t2_r1_c9_rr1;
  wire [15:0] t2_r1_c9_rr2;
  wire [15:0] t3_r1_c9_rr0;
  wire [15:0] t3_r1_c9_rr1;
  wire [15:0] t4_r1_c9_rr0;
  wire [15:0] t0_r2_c0_rr0;
  wire [15:0] t0_r2_c0_rr1;
  wire [15:0] t0_r2_c0_rr2;
  wire [15:0] t0_r2_c0_rr3;
  wire [15:0] t0_r2_c0_rr4;
  wire [15:0] t0_r2_c0_rr5;
  wire [15:0] t0_r2_c0_rr6;
  wire [15:0] t0_r2_c0_rr7;
  wire [15:0] t0_r2_c0_rr8;
  wire [15:0] t0_r2_c0_rr9;
  wire [15:0] t1_r2_c0_rr0;
  wire [15:0] t1_r2_c0_rr1;
  wire [15:0] t1_r2_c0_rr2;
  wire [15:0] t1_r2_c0_rr3;
  wire [15:0] t1_r2_c0_rr4;
  wire [15:0] t2_r2_c0_rr0;
  wire [15:0] t2_r2_c0_rr1;
  wire [15:0] t2_r2_c0_rr2;
  wire [15:0] t3_r2_c0_rr0;
  wire [15:0] t3_r2_c0_rr1;
  wire [15:0] t4_r2_c0_rr0;
  wire [15:0] t0_r2_c1_rr0;
  wire [15:0] t0_r2_c1_rr1;
  wire [15:0] t0_r2_c1_rr2;
  wire [15:0] t0_r2_c1_rr3;
  wire [15:0] t0_r2_c1_rr4;
  wire [15:0] t0_r2_c1_rr5;
  wire [15:0] t0_r2_c1_rr6;
  wire [15:0] t0_r2_c1_rr7;
  wire [15:0] t0_r2_c1_rr8;
  wire [15:0] t0_r2_c1_rr9;
  wire [15:0] t1_r2_c1_rr0;
  wire [15:0] t1_r2_c1_rr1;
  wire [15:0] t1_r2_c1_rr2;
  wire [15:0] t1_r2_c1_rr3;
  wire [15:0] t1_r2_c1_rr4;
  wire [15:0] t2_r2_c1_rr0;
  wire [15:0] t2_r2_c1_rr1;
  wire [15:0] t2_r2_c1_rr2;
  wire [15:0] t3_r2_c1_rr0;
  wire [15:0] t3_r2_c1_rr1;
  wire [15:0] t4_r2_c1_rr0;
  wire [15:0] t0_r2_c2_rr0;
  wire [15:0] t0_r2_c2_rr1;
  wire [15:0] t0_r2_c2_rr2;
  wire [15:0] t0_r2_c2_rr3;
  wire [15:0] t0_r2_c2_rr4;
  wire [15:0] t0_r2_c2_rr5;
  wire [15:0] t0_r2_c2_rr6;
  wire [15:0] t0_r2_c2_rr7;
  wire [15:0] t0_r2_c2_rr8;
  wire [15:0] t0_r2_c2_rr9;
  wire [15:0] t1_r2_c2_rr0;
  wire [15:0] t1_r2_c2_rr1;
  wire [15:0] t1_r2_c2_rr2;
  wire [15:0] t1_r2_c2_rr3;
  wire [15:0] t1_r2_c2_rr4;
  wire [15:0] t2_r2_c2_rr0;
  wire [15:0] t2_r2_c2_rr1;
  wire [15:0] t2_r2_c2_rr2;
  wire [15:0] t3_r2_c2_rr0;
  wire [15:0] t3_r2_c2_rr1;
  wire [15:0] t4_r2_c2_rr0;
  wire [15:0] t0_r2_c3_rr0;
  wire [15:0] t0_r2_c3_rr1;
  wire [15:0] t0_r2_c3_rr2;
  wire [15:0] t0_r2_c3_rr3;
  wire [15:0] t0_r2_c3_rr4;
  wire [15:0] t0_r2_c3_rr5;
  wire [15:0] t0_r2_c3_rr6;
  wire [15:0] t0_r2_c3_rr7;
  wire [15:0] t0_r2_c3_rr8;
  wire [15:0] t0_r2_c3_rr9;
  wire [15:0] t1_r2_c3_rr0;
  wire [15:0] t1_r2_c3_rr1;
  wire [15:0] t1_r2_c3_rr2;
  wire [15:0] t1_r2_c3_rr3;
  wire [15:0] t1_r2_c3_rr4;
  wire [15:0] t2_r2_c3_rr0;
  wire [15:0] t2_r2_c3_rr1;
  wire [15:0] t2_r2_c3_rr2;
  wire [15:0] t3_r2_c3_rr0;
  wire [15:0] t3_r2_c3_rr1;
  wire [15:0] t4_r2_c3_rr0;
  wire [15:0] t0_r2_c4_rr0;
  wire [15:0] t0_r2_c4_rr1;
  wire [15:0] t0_r2_c4_rr2;
  wire [15:0] t0_r2_c4_rr3;
  wire [15:0] t0_r2_c4_rr4;
  wire [15:0] t0_r2_c4_rr5;
  wire [15:0] t0_r2_c4_rr6;
  wire [15:0] t0_r2_c4_rr7;
  wire [15:0] t0_r2_c4_rr8;
  wire [15:0] t0_r2_c4_rr9;
  wire [15:0] t1_r2_c4_rr0;
  wire [15:0] t1_r2_c4_rr1;
  wire [15:0] t1_r2_c4_rr2;
  wire [15:0] t1_r2_c4_rr3;
  wire [15:0] t1_r2_c4_rr4;
  wire [15:0] t2_r2_c4_rr0;
  wire [15:0] t2_r2_c4_rr1;
  wire [15:0] t2_r2_c4_rr2;
  wire [15:0] t3_r2_c4_rr0;
  wire [15:0] t3_r2_c4_rr1;
  wire [15:0] t4_r2_c4_rr0;
  wire [15:0] t0_r2_c5_rr0;
  wire [15:0] t0_r2_c5_rr1;
  wire [15:0] t0_r2_c5_rr2;
  wire [15:0] t0_r2_c5_rr3;
  wire [15:0] t0_r2_c5_rr4;
  wire [15:0] t0_r2_c5_rr5;
  wire [15:0] t0_r2_c5_rr6;
  wire [15:0] t0_r2_c5_rr7;
  wire [15:0] t0_r2_c5_rr8;
  wire [15:0] t0_r2_c5_rr9;
  wire [15:0] t1_r2_c5_rr0;
  wire [15:0] t1_r2_c5_rr1;
  wire [15:0] t1_r2_c5_rr2;
  wire [15:0] t1_r2_c5_rr3;
  wire [15:0] t1_r2_c5_rr4;
  wire [15:0] t2_r2_c5_rr0;
  wire [15:0] t2_r2_c5_rr1;
  wire [15:0] t2_r2_c5_rr2;
  wire [15:0] t3_r2_c5_rr0;
  wire [15:0] t3_r2_c5_rr1;
  wire [15:0] t4_r2_c5_rr0;
  wire [15:0] t0_r2_c6_rr0;
  wire [15:0] t0_r2_c6_rr1;
  wire [15:0] t0_r2_c6_rr2;
  wire [15:0] t0_r2_c6_rr3;
  wire [15:0] t0_r2_c6_rr4;
  wire [15:0] t0_r2_c6_rr5;
  wire [15:0] t0_r2_c6_rr6;
  wire [15:0] t0_r2_c6_rr7;
  wire [15:0] t0_r2_c6_rr8;
  wire [15:0] t0_r2_c6_rr9;
  wire [15:0] t1_r2_c6_rr0;
  wire [15:0] t1_r2_c6_rr1;
  wire [15:0] t1_r2_c6_rr2;
  wire [15:0] t1_r2_c6_rr3;
  wire [15:0] t1_r2_c6_rr4;
  wire [15:0] t2_r2_c6_rr0;
  wire [15:0] t2_r2_c6_rr1;
  wire [15:0] t2_r2_c6_rr2;
  wire [15:0] t3_r2_c6_rr0;
  wire [15:0] t3_r2_c6_rr1;
  wire [15:0] t4_r2_c6_rr0;
  wire [15:0] t0_r2_c7_rr0;
  wire [15:0] t0_r2_c7_rr1;
  wire [15:0] t0_r2_c7_rr2;
  wire [15:0] t0_r2_c7_rr3;
  wire [15:0] t0_r2_c7_rr4;
  wire [15:0] t0_r2_c7_rr5;
  wire [15:0] t0_r2_c7_rr6;
  wire [15:0] t0_r2_c7_rr7;
  wire [15:0] t0_r2_c7_rr8;
  wire [15:0] t0_r2_c7_rr9;
  wire [15:0] t1_r2_c7_rr0;
  wire [15:0] t1_r2_c7_rr1;
  wire [15:0] t1_r2_c7_rr2;
  wire [15:0] t1_r2_c7_rr3;
  wire [15:0] t1_r2_c7_rr4;
  wire [15:0] t2_r2_c7_rr0;
  wire [15:0] t2_r2_c7_rr1;
  wire [15:0] t2_r2_c7_rr2;
  wire [15:0] t3_r2_c7_rr0;
  wire [15:0] t3_r2_c7_rr1;
  wire [15:0] t4_r2_c7_rr0;
  wire [15:0] t0_r2_c8_rr0;
  wire [15:0] t0_r2_c8_rr1;
  wire [15:0] t0_r2_c8_rr2;
  wire [15:0] t0_r2_c8_rr3;
  wire [15:0] t0_r2_c8_rr4;
  wire [15:0] t0_r2_c8_rr5;
  wire [15:0] t0_r2_c8_rr6;
  wire [15:0] t0_r2_c8_rr7;
  wire [15:0] t0_r2_c8_rr8;
  wire [15:0] t0_r2_c8_rr9;
  wire [15:0] t1_r2_c8_rr0;
  wire [15:0] t1_r2_c8_rr1;
  wire [15:0] t1_r2_c8_rr2;
  wire [15:0] t1_r2_c8_rr3;
  wire [15:0] t1_r2_c8_rr4;
  wire [15:0] t2_r2_c8_rr0;
  wire [15:0] t2_r2_c8_rr1;
  wire [15:0] t2_r2_c8_rr2;
  wire [15:0] t3_r2_c8_rr0;
  wire [15:0] t3_r2_c8_rr1;
  wire [15:0] t4_r2_c8_rr0;
  wire [15:0] t0_r2_c9_rr0;
  wire [15:0] t0_r2_c9_rr1;
  wire [15:0] t0_r2_c9_rr2;
  wire [15:0] t0_r2_c9_rr3;
  wire [15:0] t0_r2_c9_rr4;
  wire [15:0] t0_r2_c9_rr5;
  wire [15:0] t0_r2_c9_rr6;
  wire [15:0] t0_r2_c9_rr7;
  wire [15:0] t0_r2_c9_rr8;
  wire [15:0] t0_r2_c9_rr9;
  wire [15:0] t1_r2_c9_rr0;
  wire [15:0] t1_r2_c9_rr1;
  wire [15:0] t1_r2_c9_rr2;
  wire [15:0] t1_r2_c9_rr3;
  wire [15:0] t1_r2_c9_rr4;
  wire [15:0] t2_r2_c9_rr0;
  wire [15:0] t2_r2_c9_rr1;
  wire [15:0] t2_r2_c9_rr2;
  wire [15:0] t3_r2_c9_rr0;
  wire [15:0] t3_r2_c9_rr1;
  wire [15:0] t4_r2_c9_rr0;
  wire [15:0] t0_r3_c0_rr0;
  wire [15:0] t0_r3_c0_rr1;
  wire [15:0] t0_r3_c0_rr2;
  wire [15:0] t0_r3_c0_rr3;
  wire [15:0] t0_r3_c0_rr4;
  wire [15:0] t0_r3_c0_rr5;
  wire [15:0] t0_r3_c0_rr6;
  wire [15:0] t0_r3_c0_rr7;
  wire [15:0] t0_r3_c0_rr8;
  wire [15:0] t0_r3_c0_rr9;
  wire [15:0] t1_r3_c0_rr0;
  wire [15:0] t1_r3_c0_rr1;
  wire [15:0] t1_r3_c0_rr2;
  wire [15:0] t1_r3_c0_rr3;
  wire [15:0] t1_r3_c0_rr4;
  wire [15:0] t2_r3_c0_rr0;
  wire [15:0] t2_r3_c0_rr1;
  wire [15:0] t2_r3_c0_rr2;
  wire [15:0] t3_r3_c0_rr0;
  wire [15:0] t3_r3_c0_rr1;
  wire [15:0] t4_r3_c0_rr0;
  wire [15:0] t0_r3_c1_rr0;
  wire [15:0] t0_r3_c1_rr1;
  wire [15:0] t0_r3_c1_rr2;
  wire [15:0] t0_r3_c1_rr3;
  wire [15:0] t0_r3_c1_rr4;
  wire [15:0] t0_r3_c1_rr5;
  wire [15:0] t0_r3_c1_rr6;
  wire [15:0] t0_r3_c1_rr7;
  wire [15:0] t0_r3_c1_rr8;
  wire [15:0] t0_r3_c1_rr9;
  wire [15:0] t1_r3_c1_rr0;
  wire [15:0] t1_r3_c1_rr1;
  wire [15:0] t1_r3_c1_rr2;
  wire [15:0] t1_r3_c1_rr3;
  wire [15:0] t1_r3_c1_rr4;
  wire [15:0] t2_r3_c1_rr0;
  wire [15:0] t2_r3_c1_rr1;
  wire [15:0] t2_r3_c1_rr2;
  wire [15:0] t3_r3_c1_rr0;
  wire [15:0] t3_r3_c1_rr1;
  wire [15:0] t4_r3_c1_rr0;
  wire [15:0] t0_r3_c2_rr0;
  wire [15:0] t0_r3_c2_rr1;
  wire [15:0] t0_r3_c2_rr2;
  wire [15:0] t0_r3_c2_rr3;
  wire [15:0] t0_r3_c2_rr4;
  wire [15:0] t0_r3_c2_rr5;
  wire [15:0] t0_r3_c2_rr6;
  wire [15:0] t0_r3_c2_rr7;
  wire [15:0] t0_r3_c2_rr8;
  wire [15:0] t0_r3_c2_rr9;
  wire [15:0] t1_r3_c2_rr0;
  wire [15:0] t1_r3_c2_rr1;
  wire [15:0] t1_r3_c2_rr2;
  wire [15:0] t1_r3_c2_rr3;
  wire [15:0] t1_r3_c2_rr4;
  wire [15:0] t2_r3_c2_rr0;
  wire [15:0] t2_r3_c2_rr1;
  wire [15:0] t2_r3_c2_rr2;
  wire [15:0] t3_r3_c2_rr0;
  wire [15:0] t3_r3_c2_rr1;
  wire [15:0] t4_r3_c2_rr0;
  wire [15:0] t0_r3_c3_rr0;
  wire [15:0] t0_r3_c3_rr1;
  wire [15:0] t0_r3_c3_rr2;
  wire [15:0] t0_r3_c3_rr3;
  wire [15:0] t0_r3_c3_rr4;
  wire [15:0] t0_r3_c3_rr5;
  wire [15:0] t0_r3_c3_rr6;
  wire [15:0] t0_r3_c3_rr7;
  wire [15:0] t0_r3_c3_rr8;
  wire [15:0] t0_r3_c3_rr9;
  wire [15:0] t1_r3_c3_rr0;
  wire [15:0] t1_r3_c3_rr1;
  wire [15:0] t1_r3_c3_rr2;
  wire [15:0] t1_r3_c3_rr3;
  wire [15:0] t1_r3_c3_rr4;
  wire [15:0] t2_r3_c3_rr0;
  wire [15:0] t2_r3_c3_rr1;
  wire [15:0] t2_r3_c3_rr2;
  wire [15:0] t3_r3_c3_rr0;
  wire [15:0] t3_r3_c3_rr1;
  wire [15:0] t4_r3_c3_rr0;
  wire [15:0] t0_r3_c4_rr0;
  wire [15:0] t0_r3_c4_rr1;
  wire [15:0] t0_r3_c4_rr2;
  wire [15:0] t0_r3_c4_rr3;
  wire [15:0] t0_r3_c4_rr4;
  wire [15:0] t0_r3_c4_rr5;
  wire [15:0] t0_r3_c4_rr6;
  wire [15:0] t0_r3_c4_rr7;
  wire [15:0] t0_r3_c4_rr8;
  wire [15:0] t0_r3_c4_rr9;
  wire [15:0] t1_r3_c4_rr0;
  wire [15:0] t1_r3_c4_rr1;
  wire [15:0] t1_r3_c4_rr2;
  wire [15:0] t1_r3_c4_rr3;
  wire [15:0] t1_r3_c4_rr4;
  wire [15:0] t2_r3_c4_rr0;
  wire [15:0] t2_r3_c4_rr1;
  wire [15:0] t2_r3_c4_rr2;
  wire [15:0] t3_r3_c4_rr0;
  wire [15:0] t3_r3_c4_rr1;
  wire [15:0] t4_r3_c4_rr0;
  wire [15:0] t0_r3_c5_rr0;
  wire [15:0] t0_r3_c5_rr1;
  wire [15:0] t0_r3_c5_rr2;
  wire [15:0] t0_r3_c5_rr3;
  wire [15:0] t0_r3_c5_rr4;
  wire [15:0] t0_r3_c5_rr5;
  wire [15:0] t0_r3_c5_rr6;
  wire [15:0] t0_r3_c5_rr7;
  wire [15:0] t0_r3_c5_rr8;
  wire [15:0] t0_r3_c5_rr9;
  wire [15:0] t1_r3_c5_rr0;
  wire [15:0] t1_r3_c5_rr1;
  wire [15:0] t1_r3_c5_rr2;
  wire [15:0] t1_r3_c5_rr3;
  wire [15:0] t1_r3_c5_rr4;
  wire [15:0] t2_r3_c5_rr0;
  wire [15:0] t2_r3_c5_rr1;
  wire [15:0] t2_r3_c5_rr2;
  wire [15:0] t3_r3_c5_rr0;
  wire [15:0] t3_r3_c5_rr1;
  wire [15:0] t4_r3_c5_rr0;
  wire [15:0] t0_r3_c6_rr0;
  wire [15:0] t0_r3_c6_rr1;
  wire [15:0] t0_r3_c6_rr2;
  wire [15:0] t0_r3_c6_rr3;
  wire [15:0] t0_r3_c6_rr4;
  wire [15:0] t0_r3_c6_rr5;
  wire [15:0] t0_r3_c6_rr6;
  wire [15:0] t0_r3_c6_rr7;
  wire [15:0] t0_r3_c6_rr8;
  wire [15:0] t0_r3_c6_rr9;
  wire [15:0] t1_r3_c6_rr0;
  wire [15:0] t1_r3_c6_rr1;
  wire [15:0] t1_r3_c6_rr2;
  wire [15:0] t1_r3_c6_rr3;
  wire [15:0] t1_r3_c6_rr4;
  wire [15:0] t2_r3_c6_rr0;
  wire [15:0] t2_r3_c6_rr1;
  wire [15:0] t2_r3_c6_rr2;
  wire [15:0] t3_r3_c6_rr0;
  wire [15:0] t3_r3_c6_rr1;
  wire [15:0] t4_r3_c6_rr0;
  wire [15:0] t0_r3_c7_rr0;
  wire [15:0] t0_r3_c7_rr1;
  wire [15:0] t0_r3_c7_rr2;
  wire [15:0] t0_r3_c7_rr3;
  wire [15:0] t0_r3_c7_rr4;
  wire [15:0] t0_r3_c7_rr5;
  wire [15:0] t0_r3_c7_rr6;
  wire [15:0] t0_r3_c7_rr7;
  wire [15:0] t0_r3_c7_rr8;
  wire [15:0] t0_r3_c7_rr9;
  wire [15:0] t1_r3_c7_rr0;
  wire [15:0] t1_r3_c7_rr1;
  wire [15:0] t1_r3_c7_rr2;
  wire [15:0] t1_r3_c7_rr3;
  wire [15:0] t1_r3_c7_rr4;
  wire [15:0] t2_r3_c7_rr0;
  wire [15:0] t2_r3_c7_rr1;
  wire [15:0] t2_r3_c7_rr2;
  wire [15:0] t3_r3_c7_rr0;
  wire [15:0] t3_r3_c7_rr1;
  wire [15:0] t4_r3_c7_rr0;
  wire [15:0] t0_r3_c8_rr0;
  wire [15:0] t0_r3_c8_rr1;
  wire [15:0] t0_r3_c8_rr2;
  wire [15:0] t0_r3_c8_rr3;
  wire [15:0] t0_r3_c8_rr4;
  wire [15:0] t0_r3_c8_rr5;
  wire [15:0] t0_r3_c8_rr6;
  wire [15:0] t0_r3_c8_rr7;
  wire [15:0] t0_r3_c8_rr8;
  wire [15:0] t0_r3_c8_rr9;
  wire [15:0] t1_r3_c8_rr0;
  wire [15:0] t1_r3_c8_rr1;
  wire [15:0] t1_r3_c8_rr2;
  wire [15:0] t1_r3_c8_rr3;
  wire [15:0] t1_r3_c8_rr4;
  wire [15:0] t2_r3_c8_rr0;
  wire [15:0] t2_r3_c8_rr1;
  wire [15:0] t2_r3_c8_rr2;
  wire [15:0] t3_r3_c8_rr0;
  wire [15:0] t3_r3_c8_rr1;
  wire [15:0] t4_r3_c8_rr0;
  wire [15:0] t0_r3_c9_rr0;
  wire [15:0] t0_r3_c9_rr1;
  wire [15:0] t0_r3_c9_rr2;
  wire [15:0] t0_r3_c9_rr3;
  wire [15:0] t0_r3_c9_rr4;
  wire [15:0] t0_r3_c9_rr5;
  wire [15:0] t0_r3_c9_rr6;
  wire [15:0] t0_r3_c9_rr7;
  wire [15:0] t0_r3_c9_rr8;
  wire [15:0] t0_r3_c9_rr9;
  wire [15:0] t1_r3_c9_rr0;
  wire [15:0] t1_r3_c9_rr1;
  wire [15:0] t1_r3_c9_rr2;
  wire [15:0] t1_r3_c9_rr3;
  wire [15:0] t1_r3_c9_rr4;
  wire [15:0] t2_r3_c9_rr0;
  wire [15:0] t2_r3_c9_rr1;
  wire [15:0] t2_r3_c9_rr2;
  wire [15:0] t3_r3_c9_rr0;
  wire [15:0] t3_r3_c9_rr1;
  wire [15:0] t4_r3_c9_rr0;
  wire [15:0] t0_r4_c0_rr0;
  wire [15:0] t0_r4_c0_rr1;
  wire [15:0] t0_r4_c0_rr2;
  wire [15:0] t0_r4_c0_rr3;
  wire [15:0] t0_r4_c0_rr4;
  wire [15:0] t0_r4_c0_rr5;
  wire [15:0] t0_r4_c0_rr6;
  wire [15:0] t0_r4_c0_rr7;
  wire [15:0] t0_r4_c0_rr8;
  wire [15:0] t0_r4_c0_rr9;
  wire [15:0] t1_r4_c0_rr0;
  wire [15:0] t1_r4_c0_rr1;
  wire [15:0] t1_r4_c0_rr2;
  wire [15:0] t1_r4_c0_rr3;
  wire [15:0] t1_r4_c0_rr4;
  wire [15:0] t2_r4_c0_rr0;
  wire [15:0] t2_r4_c0_rr1;
  wire [15:0] t2_r4_c0_rr2;
  wire [15:0] t3_r4_c0_rr0;
  wire [15:0] t3_r4_c0_rr1;
  wire [15:0] t4_r4_c0_rr0;
  wire [15:0] t0_r4_c1_rr0;
  wire [15:0] t0_r4_c1_rr1;
  wire [15:0] t0_r4_c1_rr2;
  wire [15:0] t0_r4_c1_rr3;
  wire [15:0] t0_r4_c1_rr4;
  wire [15:0] t0_r4_c1_rr5;
  wire [15:0] t0_r4_c1_rr6;
  wire [15:0] t0_r4_c1_rr7;
  wire [15:0] t0_r4_c1_rr8;
  wire [15:0] t0_r4_c1_rr9;
  wire [15:0] t1_r4_c1_rr0;
  wire [15:0] t1_r4_c1_rr1;
  wire [15:0] t1_r4_c1_rr2;
  wire [15:0] t1_r4_c1_rr3;
  wire [15:0] t1_r4_c1_rr4;
  wire [15:0] t2_r4_c1_rr0;
  wire [15:0] t2_r4_c1_rr1;
  wire [15:0] t2_r4_c1_rr2;
  wire [15:0] t3_r4_c1_rr0;
  wire [15:0] t3_r4_c1_rr1;
  wire [15:0] t4_r4_c1_rr0;
  wire [15:0] t0_r4_c2_rr0;
  wire [15:0] t0_r4_c2_rr1;
  wire [15:0] t0_r4_c2_rr2;
  wire [15:0] t0_r4_c2_rr3;
  wire [15:0] t0_r4_c2_rr4;
  wire [15:0] t0_r4_c2_rr5;
  wire [15:0] t0_r4_c2_rr6;
  wire [15:0] t0_r4_c2_rr7;
  wire [15:0] t0_r4_c2_rr8;
  wire [15:0] t0_r4_c2_rr9;
  wire [15:0] t1_r4_c2_rr0;
  wire [15:0] t1_r4_c2_rr1;
  wire [15:0] t1_r4_c2_rr2;
  wire [15:0] t1_r4_c2_rr3;
  wire [15:0] t1_r4_c2_rr4;
  wire [15:0] t2_r4_c2_rr0;
  wire [15:0] t2_r4_c2_rr1;
  wire [15:0] t2_r4_c2_rr2;
  wire [15:0] t3_r4_c2_rr0;
  wire [15:0] t3_r4_c2_rr1;
  wire [15:0] t4_r4_c2_rr0;
  wire [15:0] t0_r4_c3_rr0;
  wire [15:0] t0_r4_c3_rr1;
  wire [15:0] t0_r4_c3_rr2;
  wire [15:0] t0_r4_c3_rr3;
  wire [15:0] t0_r4_c3_rr4;
  wire [15:0] t0_r4_c3_rr5;
  wire [15:0] t0_r4_c3_rr6;
  wire [15:0] t0_r4_c3_rr7;
  wire [15:0] t0_r4_c3_rr8;
  wire [15:0] t0_r4_c3_rr9;
  wire [15:0] t1_r4_c3_rr0;
  wire [15:0] t1_r4_c3_rr1;
  wire [15:0] t1_r4_c3_rr2;
  wire [15:0] t1_r4_c3_rr3;
  wire [15:0] t1_r4_c3_rr4;
  wire [15:0] t2_r4_c3_rr0;
  wire [15:0] t2_r4_c3_rr1;
  wire [15:0] t2_r4_c3_rr2;
  wire [15:0] t3_r4_c3_rr0;
  wire [15:0] t3_r4_c3_rr1;
  wire [15:0] t4_r4_c3_rr0;
  wire [15:0] t0_r4_c4_rr0;
  wire [15:0] t0_r4_c4_rr1;
  wire [15:0] t0_r4_c4_rr2;
  wire [15:0] t0_r4_c4_rr3;
  wire [15:0] t0_r4_c4_rr4;
  wire [15:0] t0_r4_c4_rr5;
  wire [15:0] t0_r4_c4_rr6;
  wire [15:0] t0_r4_c4_rr7;
  wire [15:0] t0_r4_c4_rr8;
  wire [15:0] t0_r4_c4_rr9;
  wire [15:0] t1_r4_c4_rr0;
  wire [15:0] t1_r4_c4_rr1;
  wire [15:0] t1_r4_c4_rr2;
  wire [15:0] t1_r4_c4_rr3;
  wire [15:0] t1_r4_c4_rr4;
  wire [15:0] t2_r4_c4_rr0;
  wire [15:0] t2_r4_c4_rr1;
  wire [15:0] t2_r4_c4_rr2;
  wire [15:0] t3_r4_c4_rr0;
  wire [15:0] t3_r4_c4_rr1;
  wire [15:0] t4_r4_c4_rr0;
  wire [15:0] t0_r4_c5_rr0;
  wire [15:0] t0_r4_c5_rr1;
  wire [15:0] t0_r4_c5_rr2;
  wire [15:0] t0_r4_c5_rr3;
  wire [15:0] t0_r4_c5_rr4;
  wire [15:0] t0_r4_c5_rr5;
  wire [15:0] t0_r4_c5_rr6;
  wire [15:0] t0_r4_c5_rr7;
  wire [15:0] t0_r4_c5_rr8;
  wire [15:0] t0_r4_c5_rr9;
  wire [15:0] t1_r4_c5_rr0;
  wire [15:0] t1_r4_c5_rr1;
  wire [15:0] t1_r4_c5_rr2;
  wire [15:0] t1_r4_c5_rr3;
  wire [15:0] t1_r4_c5_rr4;
  wire [15:0] t2_r4_c5_rr0;
  wire [15:0] t2_r4_c5_rr1;
  wire [15:0] t2_r4_c5_rr2;
  wire [15:0] t3_r4_c5_rr0;
  wire [15:0] t3_r4_c5_rr1;
  wire [15:0] t4_r4_c5_rr0;
  wire [15:0] t0_r4_c6_rr0;
  wire [15:0] t0_r4_c6_rr1;
  wire [15:0] t0_r4_c6_rr2;
  wire [15:0] t0_r4_c6_rr3;
  wire [15:0] t0_r4_c6_rr4;
  wire [15:0] t0_r4_c6_rr5;
  wire [15:0] t0_r4_c6_rr6;
  wire [15:0] t0_r4_c6_rr7;
  wire [15:0] t0_r4_c6_rr8;
  wire [15:0] t0_r4_c6_rr9;
  wire [15:0] t1_r4_c6_rr0;
  wire [15:0] t1_r4_c6_rr1;
  wire [15:0] t1_r4_c6_rr2;
  wire [15:0] t1_r4_c6_rr3;
  wire [15:0] t1_r4_c6_rr4;
  wire [15:0] t2_r4_c6_rr0;
  wire [15:0] t2_r4_c6_rr1;
  wire [15:0] t2_r4_c6_rr2;
  wire [15:0] t3_r4_c6_rr0;
  wire [15:0] t3_r4_c6_rr1;
  wire [15:0] t4_r4_c6_rr0;
  wire [15:0] t0_r4_c7_rr0;
  wire [15:0] t0_r4_c7_rr1;
  wire [15:0] t0_r4_c7_rr2;
  wire [15:0] t0_r4_c7_rr3;
  wire [15:0] t0_r4_c7_rr4;
  wire [15:0] t0_r4_c7_rr5;
  wire [15:0] t0_r4_c7_rr6;
  wire [15:0] t0_r4_c7_rr7;
  wire [15:0] t0_r4_c7_rr8;
  wire [15:0] t0_r4_c7_rr9;
  wire [15:0] t1_r4_c7_rr0;
  wire [15:0] t1_r4_c7_rr1;
  wire [15:0] t1_r4_c7_rr2;
  wire [15:0] t1_r4_c7_rr3;
  wire [15:0] t1_r4_c7_rr4;
  wire [15:0] t2_r4_c7_rr0;
  wire [15:0] t2_r4_c7_rr1;
  wire [15:0] t2_r4_c7_rr2;
  wire [15:0] t3_r4_c7_rr0;
  wire [15:0] t3_r4_c7_rr1;
  wire [15:0] t4_r4_c7_rr0;
  wire [15:0] t0_r4_c8_rr0;
  wire [15:0] t0_r4_c8_rr1;
  wire [15:0] t0_r4_c8_rr2;
  wire [15:0] t0_r4_c8_rr3;
  wire [15:0] t0_r4_c8_rr4;
  wire [15:0] t0_r4_c8_rr5;
  wire [15:0] t0_r4_c8_rr6;
  wire [15:0] t0_r4_c8_rr7;
  wire [15:0] t0_r4_c8_rr8;
  wire [15:0] t0_r4_c8_rr9;
  wire [15:0] t1_r4_c8_rr0;
  wire [15:0] t1_r4_c8_rr1;
  wire [15:0] t1_r4_c8_rr2;
  wire [15:0] t1_r4_c8_rr3;
  wire [15:0] t1_r4_c8_rr4;
  wire [15:0] t2_r4_c8_rr0;
  wire [15:0] t2_r4_c8_rr1;
  wire [15:0] t2_r4_c8_rr2;
  wire [15:0] t3_r4_c8_rr0;
  wire [15:0] t3_r4_c8_rr1;
  wire [15:0] t4_r4_c8_rr0;
  wire [15:0] t0_r4_c9_rr0;
  wire [15:0] t0_r4_c9_rr1;
  wire [15:0] t0_r4_c9_rr2;
  wire [15:0] t0_r4_c9_rr3;
  wire [15:0] t0_r4_c9_rr4;
  wire [15:0] t0_r4_c9_rr5;
  wire [15:0] t0_r4_c9_rr6;
  wire [15:0] t0_r4_c9_rr7;
  wire [15:0] t0_r4_c9_rr8;
  wire [15:0] t0_r4_c9_rr9;
  wire [15:0] t1_r4_c9_rr0;
  wire [15:0] t1_r4_c9_rr1;
  wire [15:0] t1_r4_c9_rr2;
  wire [15:0] t1_r4_c9_rr3;
  wire [15:0] t1_r4_c9_rr4;
  wire [15:0] t2_r4_c9_rr0;
  wire [15:0] t2_r4_c9_rr1;
  wire [15:0] t2_r4_c9_rr2;
  wire [15:0] t3_r4_c9_rr0;
  wire [15:0] t3_r4_c9_rr1;
  wire [15:0] t4_r4_c9_rr0;
  wire [15:0] t0_r5_c0_rr0;
  wire [15:0] t0_r5_c0_rr1;
  wire [15:0] t0_r5_c0_rr2;
  wire [15:0] t0_r5_c0_rr3;
  wire [15:0] t0_r5_c0_rr4;
  wire [15:0] t0_r5_c0_rr5;
  wire [15:0] t0_r5_c0_rr6;
  wire [15:0] t0_r5_c0_rr7;
  wire [15:0] t0_r5_c0_rr8;
  wire [15:0] t0_r5_c0_rr9;
  wire [15:0] t1_r5_c0_rr0;
  wire [15:0] t1_r5_c0_rr1;
  wire [15:0] t1_r5_c0_rr2;
  wire [15:0] t1_r5_c0_rr3;
  wire [15:0] t1_r5_c0_rr4;
  wire [15:0] t2_r5_c0_rr0;
  wire [15:0] t2_r5_c0_rr1;
  wire [15:0] t2_r5_c0_rr2;
  wire [15:0] t3_r5_c0_rr0;
  wire [15:0] t3_r5_c0_rr1;
  wire [15:0] t4_r5_c0_rr0;
  wire [15:0] t0_r5_c1_rr0;
  wire [15:0] t0_r5_c1_rr1;
  wire [15:0] t0_r5_c1_rr2;
  wire [15:0] t0_r5_c1_rr3;
  wire [15:0] t0_r5_c1_rr4;
  wire [15:0] t0_r5_c1_rr5;
  wire [15:0] t0_r5_c1_rr6;
  wire [15:0] t0_r5_c1_rr7;
  wire [15:0] t0_r5_c1_rr8;
  wire [15:0] t0_r5_c1_rr9;
  wire [15:0] t1_r5_c1_rr0;
  wire [15:0] t1_r5_c1_rr1;
  wire [15:0] t1_r5_c1_rr2;
  wire [15:0] t1_r5_c1_rr3;
  wire [15:0] t1_r5_c1_rr4;
  wire [15:0] t2_r5_c1_rr0;
  wire [15:0] t2_r5_c1_rr1;
  wire [15:0] t2_r5_c1_rr2;
  wire [15:0] t3_r5_c1_rr0;
  wire [15:0] t3_r5_c1_rr1;
  wire [15:0] t4_r5_c1_rr0;
  wire [15:0] t0_r5_c2_rr0;
  wire [15:0] t0_r5_c2_rr1;
  wire [15:0] t0_r5_c2_rr2;
  wire [15:0] t0_r5_c2_rr3;
  wire [15:0] t0_r5_c2_rr4;
  wire [15:0] t0_r5_c2_rr5;
  wire [15:0] t0_r5_c2_rr6;
  wire [15:0] t0_r5_c2_rr7;
  wire [15:0] t0_r5_c2_rr8;
  wire [15:0] t0_r5_c2_rr9;
  wire [15:0] t1_r5_c2_rr0;
  wire [15:0] t1_r5_c2_rr1;
  wire [15:0] t1_r5_c2_rr2;
  wire [15:0] t1_r5_c2_rr3;
  wire [15:0] t1_r5_c2_rr4;
  wire [15:0] t2_r5_c2_rr0;
  wire [15:0] t2_r5_c2_rr1;
  wire [15:0] t2_r5_c2_rr2;
  wire [15:0] t3_r5_c2_rr0;
  wire [15:0] t3_r5_c2_rr1;
  wire [15:0] t4_r5_c2_rr0;
  wire [15:0] t0_r5_c3_rr0;
  wire [15:0] t0_r5_c3_rr1;
  wire [15:0] t0_r5_c3_rr2;
  wire [15:0] t0_r5_c3_rr3;
  wire [15:0] t0_r5_c3_rr4;
  wire [15:0] t0_r5_c3_rr5;
  wire [15:0] t0_r5_c3_rr6;
  wire [15:0] t0_r5_c3_rr7;
  wire [15:0] t0_r5_c3_rr8;
  wire [15:0] t0_r5_c3_rr9;
  wire [15:0] t1_r5_c3_rr0;
  wire [15:0] t1_r5_c3_rr1;
  wire [15:0] t1_r5_c3_rr2;
  wire [15:0] t1_r5_c3_rr3;
  wire [15:0] t1_r5_c3_rr4;
  wire [15:0] t2_r5_c3_rr0;
  wire [15:0] t2_r5_c3_rr1;
  wire [15:0] t2_r5_c3_rr2;
  wire [15:0] t3_r5_c3_rr0;
  wire [15:0] t3_r5_c3_rr1;
  wire [15:0] t4_r5_c3_rr0;
  wire [15:0] t0_r5_c4_rr0;
  wire [15:0] t0_r5_c4_rr1;
  wire [15:0] t0_r5_c4_rr2;
  wire [15:0] t0_r5_c4_rr3;
  wire [15:0] t0_r5_c4_rr4;
  wire [15:0] t0_r5_c4_rr5;
  wire [15:0] t0_r5_c4_rr6;
  wire [15:0] t0_r5_c4_rr7;
  wire [15:0] t0_r5_c4_rr8;
  wire [15:0] t0_r5_c4_rr9;
  wire [15:0] t1_r5_c4_rr0;
  wire [15:0] t1_r5_c4_rr1;
  wire [15:0] t1_r5_c4_rr2;
  wire [15:0] t1_r5_c4_rr3;
  wire [15:0] t1_r5_c4_rr4;
  wire [15:0] t2_r5_c4_rr0;
  wire [15:0] t2_r5_c4_rr1;
  wire [15:0] t2_r5_c4_rr2;
  wire [15:0] t3_r5_c4_rr0;
  wire [15:0] t3_r5_c4_rr1;
  wire [15:0] t4_r5_c4_rr0;
  wire [15:0] t0_r5_c5_rr0;
  wire [15:0] t0_r5_c5_rr1;
  wire [15:0] t0_r5_c5_rr2;
  wire [15:0] t0_r5_c5_rr3;
  wire [15:0] t0_r5_c5_rr4;
  wire [15:0] t0_r5_c5_rr5;
  wire [15:0] t0_r5_c5_rr6;
  wire [15:0] t0_r5_c5_rr7;
  wire [15:0] t0_r5_c5_rr8;
  wire [15:0] t0_r5_c5_rr9;
  wire [15:0] t1_r5_c5_rr0;
  wire [15:0] t1_r5_c5_rr1;
  wire [15:0] t1_r5_c5_rr2;
  wire [15:0] t1_r5_c5_rr3;
  wire [15:0] t1_r5_c5_rr4;
  wire [15:0] t2_r5_c5_rr0;
  wire [15:0] t2_r5_c5_rr1;
  wire [15:0] t2_r5_c5_rr2;
  wire [15:0] t3_r5_c5_rr0;
  wire [15:0] t3_r5_c5_rr1;
  wire [15:0] t4_r5_c5_rr0;
  wire [15:0] t0_r5_c6_rr0;
  wire [15:0] t0_r5_c6_rr1;
  wire [15:0] t0_r5_c6_rr2;
  wire [15:0] t0_r5_c6_rr3;
  wire [15:0] t0_r5_c6_rr4;
  wire [15:0] t0_r5_c6_rr5;
  wire [15:0] t0_r5_c6_rr6;
  wire [15:0] t0_r5_c6_rr7;
  wire [15:0] t0_r5_c6_rr8;
  wire [15:0] t0_r5_c6_rr9;
  wire [15:0] t1_r5_c6_rr0;
  wire [15:0] t1_r5_c6_rr1;
  wire [15:0] t1_r5_c6_rr2;
  wire [15:0] t1_r5_c6_rr3;
  wire [15:0] t1_r5_c6_rr4;
  wire [15:0] t2_r5_c6_rr0;
  wire [15:0] t2_r5_c6_rr1;
  wire [15:0] t2_r5_c6_rr2;
  wire [15:0] t3_r5_c6_rr0;
  wire [15:0] t3_r5_c6_rr1;
  wire [15:0] t4_r5_c6_rr0;
  wire [15:0] t0_r5_c7_rr0;
  wire [15:0] t0_r5_c7_rr1;
  wire [15:0] t0_r5_c7_rr2;
  wire [15:0] t0_r5_c7_rr3;
  wire [15:0] t0_r5_c7_rr4;
  wire [15:0] t0_r5_c7_rr5;
  wire [15:0] t0_r5_c7_rr6;
  wire [15:0] t0_r5_c7_rr7;
  wire [15:0] t0_r5_c7_rr8;
  wire [15:0] t0_r5_c7_rr9;
  wire [15:0] t1_r5_c7_rr0;
  wire [15:0] t1_r5_c7_rr1;
  wire [15:0] t1_r5_c7_rr2;
  wire [15:0] t1_r5_c7_rr3;
  wire [15:0] t1_r5_c7_rr4;
  wire [15:0] t2_r5_c7_rr0;
  wire [15:0] t2_r5_c7_rr1;
  wire [15:0] t2_r5_c7_rr2;
  wire [15:0] t3_r5_c7_rr0;
  wire [15:0] t3_r5_c7_rr1;
  wire [15:0] t4_r5_c7_rr0;
  wire [15:0] t0_r5_c8_rr0;
  wire [15:0] t0_r5_c8_rr1;
  wire [15:0] t0_r5_c8_rr2;
  wire [15:0] t0_r5_c8_rr3;
  wire [15:0] t0_r5_c8_rr4;
  wire [15:0] t0_r5_c8_rr5;
  wire [15:0] t0_r5_c8_rr6;
  wire [15:0] t0_r5_c8_rr7;
  wire [15:0] t0_r5_c8_rr8;
  wire [15:0] t0_r5_c8_rr9;
  wire [15:0] t1_r5_c8_rr0;
  wire [15:0] t1_r5_c8_rr1;
  wire [15:0] t1_r5_c8_rr2;
  wire [15:0] t1_r5_c8_rr3;
  wire [15:0] t1_r5_c8_rr4;
  wire [15:0] t2_r5_c8_rr0;
  wire [15:0] t2_r5_c8_rr1;
  wire [15:0] t2_r5_c8_rr2;
  wire [15:0] t3_r5_c8_rr0;
  wire [15:0] t3_r5_c8_rr1;
  wire [15:0] t4_r5_c8_rr0;
  wire [15:0] t0_r5_c9_rr0;
  wire [15:0] t0_r5_c9_rr1;
  wire [15:0] t0_r5_c9_rr2;
  wire [15:0] t0_r5_c9_rr3;
  wire [15:0] t0_r5_c9_rr4;
  wire [15:0] t0_r5_c9_rr5;
  wire [15:0] t0_r5_c9_rr6;
  wire [15:0] t0_r5_c9_rr7;
  wire [15:0] t0_r5_c9_rr8;
  wire [15:0] t0_r5_c9_rr9;
  wire [15:0] t1_r5_c9_rr0;
  wire [15:0] t1_r5_c9_rr1;
  wire [15:0] t1_r5_c9_rr2;
  wire [15:0] t1_r5_c9_rr3;
  wire [15:0] t1_r5_c9_rr4;
  wire [15:0] t2_r5_c9_rr0;
  wire [15:0] t2_r5_c9_rr1;
  wire [15:0] t2_r5_c9_rr2;
  wire [15:0] t3_r5_c9_rr0;
  wire [15:0] t3_r5_c9_rr1;
  wire [15:0] t4_r5_c9_rr0;
  wire [15:0] t0_r6_c0_rr0;
  wire [15:0] t0_r6_c0_rr1;
  wire [15:0] t0_r6_c0_rr2;
  wire [15:0] t0_r6_c0_rr3;
  wire [15:0] t0_r6_c0_rr4;
  wire [15:0] t0_r6_c0_rr5;
  wire [15:0] t0_r6_c0_rr6;
  wire [15:0] t0_r6_c0_rr7;
  wire [15:0] t0_r6_c0_rr8;
  wire [15:0] t0_r6_c0_rr9;
  wire [15:0] t1_r6_c0_rr0;
  wire [15:0] t1_r6_c0_rr1;
  wire [15:0] t1_r6_c0_rr2;
  wire [15:0] t1_r6_c0_rr3;
  wire [15:0] t1_r6_c0_rr4;
  wire [15:0] t2_r6_c0_rr0;
  wire [15:0] t2_r6_c0_rr1;
  wire [15:0] t2_r6_c0_rr2;
  wire [15:0] t3_r6_c0_rr0;
  wire [15:0] t3_r6_c0_rr1;
  wire [15:0] t4_r6_c0_rr0;
  wire [15:0] t0_r6_c1_rr0;
  wire [15:0] t0_r6_c1_rr1;
  wire [15:0] t0_r6_c1_rr2;
  wire [15:0] t0_r6_c1_rr3;
  wire [15:0] t0_r6_c1_rr4;
  wire [15:0] t0_r6_c1_rr5;
  wire [15:0] t0_r6_c1_rr6;
  wire [15:0] t0_r6_c1_rr7;
  wire [15:0] t0_r6_c1_rr8;
  wire [15:0] t0_r6_c1_rr9;
  wire [15:0] t1_r6_c1_rr0;
  wire [15:0] t1_r6_c1_rr1;
  wire [15:0] t1_r6_c1_rr2;
  wire [15:0] t1_r6_c1_rr3;
  wire [15:0] t1_r6_c1_rr4;
  wire [15:0] t2_r6_c1_rr0;
  wire [15:0] t2_r6_c1_rr1;
  wire [15:0] t2_r6_c1_rr2;
  wire [15:0] t3_r6_c1_rr0;
  wire [15:0] t3_r6_c1_rr1;
  wire [15:0] t4_r6_c1_rr0;
  wire [15:0] t0_r6_c2_rr0;
  wire [15:0] t0_r6_c2_rr1;
  wire [15:0] t0_r6_c2_rr2;
  wire [15:0] t0_r6_c2_rr3;
  wire [15:0] t0_r6_c2_rr4;
  wire [15:0] t0_r6_c2_rr5;
  wire [15:0] t0_r6_c2_rr6;
  wire [15:0] t0_r6_c2_rr7;
  wire [15:0] t0_r6_c2_rr8;
  wire [15:0] t0_r6_c2_rr9;
  wire [15:0] t1_r6_c2_rr0;
  wire [15:0] t1_r6_c2_rr1;
  wire [15:0] t1_r6_c2_rr2;
  wire [15:0] t1_r6_c2_rr3;
  wire [15:0] t1_r6_c2_rr4;
  wire [15:0] t2_r6_c2_rr0;
  wire [15:0] t2_r6_c2_rr1;
  wire [15:0] t2_r6_c2_rr2;
  wire [15:0] t3_r6_c2_rr0;
  wire [15:0] t3_r6_c2_rr1;
  wire [15:0] t4_r6_c2_rr0;
  wire [15:0] t0_r6_c3_rr0;
  wire [15:0] t0_r6_c3_rr1;
  wire [15:0] t0_r6_c3_rr2;
  wire [15:0] t0_r6_c3_rr3;
  wire [15:0] t0_r6_c3_rr4;
  wire [15:0] t0_r6_c3_rr5;
  wire [15:0] t0_r6_c3_rr6;
  wire [15:0] t0_r6_c3_rr7;
  wire [15:0] t0_r6_c3_rr8;
  wire [15:0] t0_r6_c3_rr9;
  wire [15:0] t1_r6_c3_rr0;
  wire [15:0] t1_r6_c3_rr1;
  wire [15:0] t1_r6_c3_rr2;
  wire [15:0] t1_r6_c3_rr3;
  wire [15:0] t1_r6_c3_rr4;
  wire [15:0] t2_r6_c3_rr0;
  wire [15:0] t2_r6_c3_rr1;
  wire [15:0] t2_r6_c3_rr2;
  wire [15:0] t3_r6_c3_rr0;
  wire [15:0] t3_r6_c3_rr1;
  wire [15:0] t4_r6_c3_rr0;
  wire [15:0] t0_r6_c4_rr0;
  wire [15:0] t0_r6_c4_rr1;
  wire [15:0] t0_r6_c4_rr2;
  wire [15:0] t0_r6_c4_rr3;
  wire [15:0] t0_r6_c4_rr4;
  wire [15:0] t0_r6_c4_rr5;
  wire [15:0] t0_r6_c4_rr6;
  wire [15:0] t0_r6_c4_rr7;
  wire [15:0] t0_r6_c4_rr8;
  wire [15:0] t0_r6_c4_rr9;
  wire [15:0] t1_r6_c4_rr0;
  wire [15:0] t1_r6_c4_rr1;
  wire [15:0] t1_r6_c4_rr2;
  wire [15:0] t1_r6_c4_rr3;
  wire [15:0] t1_r6_c4_rr4;
  wire [15:0] t2_r6_c4_rr0;
  wire [15:0] t2_r6_c4_rr1;
  wire [15:0] t2_r6_c4_rr2;
  wire [15:0] t3_r6_c4_rr0;
  wire [15:0] t3_r6_c4_rr1;
  wire [15:0] t4_r6_c4_rr0;
  wire [15:0] t0_r6_c5_rr0;
  wire [15:0] t0_r6_c5_rr1;
  wire [15:0] t0_r6_c5_rr2;
  wire [15:0] t0_r6_c5_rr3;
  wire [15:0] t0_r6_c5_rr4;
  wire [15:0] t0_r6_c5_rr5;
  wire [15:0] t0_r6_c5_rr6;
  wire [15:0] t0_r6_c5_rr7;
  wire [15:0] t0_r6_c5_rr8;
  wire [15:0] t0_r6_c5_rr9;
  wire [15:0] t1_r6_c5_rr0;
  wire [15:0] t1_r6_c5_rr1;
  wire [15:0] t1_r6_c5_rr2;
  wire [15:0] t1_r6_c5_rr3;
  wire [15:0] t1_r6_c5_rr4;
  wire [15:0] t2_r6_c5_rr0;
  wire [15:0] t2_r6_c5_rr1;
  wire [15:0] t2_r6_c5_rr2;
  wire [15:0] t3_r6_c5_rr0;
  wire [15:0] t3_r6_c5_rr1;
  wire [15:0] t4_r6_c5_rr0;
  wire [15:0] t0_r6_c6_rr0;
  wire [15:0] t0_r6_c6_rr1;
  wire [15:0] t0_r6_c6_rr2;
  wire [15:0] t0_r6_c6_rr3;
  wire [15:0] t0_r6_c6_rr4;
  wire [15:0] t0_r6_c6_rr5;
  wire [15:0] t0_r6_c6_rr6;
  wire [15:0] t0_r6_c6_rr7;
  wire [15:0] t0_r6_c6_rr8;
  wire [15:0] t0_r6_c6_rr9;
  wire [15:0] t1_r6_c6_rr0;
  wire [15:0] t1_r6_c6_rr1;
  wire [15:0] t1_r6_c6_rr2;
  wire [15:0] t1_r6_c6_rr3;
  wire [15:0] t1_r6_c6_rr4;
  wire [15:0] t2_r6_c6_rr0;
  wire [15:0] t2_r6_c6_rr1;
  wire [15:0] t2_r6_c6_rr2;
  wire [15:0] t3_r6_c6_rr0;
  wire [15:0] t3_r6_c6_rr1;
  wire [15:0] t4_r6_c6_rr0;
  wire [15:0] t0_r6_c7_rr0;
  wire [15:0] t0_r6_c7_rr1;
  wire [15:0] t0_r6_c7_rr2;
  wire [15:0] t0_r6_c7_rr3;
  wire [15:0] t0_r6_c7_rr4;
  wire [15:0] t0_r6_c7_rr5;
  wire [15:0] t0_r6_c7_rr6;
  wire [15:0] t0_r6_c7_rr7;
  wire [15:0] t0_r6_c7_rr8;
  wire [15:0] t0_r6_c7_rr9;
  wire [15:0] t1_r6_c7_rr0;
  wire [15:0] t1_r6_c7_rr1;
  wire [15:0] t1_r6_c7_rr2;
  wire [15:0] t1_r6_c7_rr3;
  wire [15:0] t1_r6_c7_rr4;
  wire [15:0] t2_r6_c7_rr0;
  wire [15:0] t2_r6_c7_rr1;
  wire [15:0] t2_r6_c7_rr2;
  wire [15:0] t3_r6_c7_rr0;
  wire [15:0] t3_r6_c7_rr1;
  wire [15:0] t4_r6_c7_rr0;
  wire [15:0] t0_r6_c8_rr0;
  wire [15:0] t0_r6_c8_rr1;
  wire [15:0] t0_r6_c8_rr2;
  wire [15:0] t0_r6_c8_rr3;
  wire [15:0] t0_r6_c8_rr4;
  wire [15:0] t0_r6_c8_rr5;
  wire [15:0] t0_r6_c8_rr6;
  wire [15:0] t0_r6_c8_rr7;
  wire [15:0] t0_r6_c8_rr8;
  wire [15:0] t0_r6_c8_rr9;
  wire [15:0] t1_r6_c8_rr0;
  wire [15:0] t1_r6_c8_rr1;
  wire [15:0] t1_r6_c8_rr2;
  wire [15:0] t1_r6_c8_rr3;
  wire [15:0] t1_r6_c8_rr4;
  wire [15:0] t2_r6_c8_rr0;
  wire [15:0] t2_r6_c8_rr1;
  wire [15:0] t2_r6_c8_rr2;
  wire [15:0] t3_r6_c8_rr0;
  wire [15:0] t3_r6_c8_rr1;
  wire [15:0] t4_r6_c8_rr0;
  wire [15:0] t0_r6_c9_rr0;
  wire [15:0] t0_r6_c9_rr1;
  wire [15:0] t0_r6_c9_rr2;
  wire [15:0] t0_r6_c9_rr3;
  wire [15:0] t0_r6_c9_rr4;
  wire [15:0] t0_r6_c9_rr5;
  wire [15:0] t0_r6_c9_rr6;
  wire [15:0] t0_r6_c9_rr7;
  wire [15:0] t0_r6_c9_rr8;
  wire [15:0] t0_r6_c9_rr9;
  wire [15:0] t1_r6_c9_rr0;
  wire [15:0] t1_r6_c9_rr1;
  wire [15:0] t1_r6_c9_rr2;
  wire [15:0] t1_r6_c9_rr3;
  wire [15:0] t1_r6_c9_rr4;
  wire [15:0] t2_r6_c9_rr0;
  wire [15:0] t2_r6_c9_rr1;
  wire [15:0] t2_r6_c9_rr2;
  wire [15:0] t3_r6_c9_rr0;
  wire [15:0] t3_r6_c9_rr1;
  wire [15:0] t4_r6_c9_rr0;
  wire [15:0] t0_r7_c0_rr0;
  wire [15:0] t0_r7_c0_rr1;
  wire [15:0] t0_r7_c0_rr2;
  wire [15:0] t0_r7_c0_rr3;
  wire [15:0] t0_r7_c0_rr4;
  wire [15:0] t0_r7_c0_rr5;
  wire [15:0] t0_r7_c0_rr6;
  wire [15:0] t0_r7_c0_rr7;
  wire [15:0] t0_r7_c0_rr8;
  wire [15:0] t0_r7_c0_rr9;
  wire [15:0] t1_r7_c0_rr0;
  wire [15:0] t1_r7_c0_rr1;
  wire [15:0] t1_r7_c0_rr2;
  wire [15:0] t1_r7_c0_rr3;
  wire [15:0] t1_r7_c0_rr4;
  wire [15:0] t2_r7_c0_rr0;
  wire [15:0] t2_r7_c0_rr1;
  wire [15:0] t2_r7_c0_rr2;
  wire [15:0] t3_r7_c0_rr0;
  wire [15:0] t3_r7_c0_rr1;
  wire [15:0] t4_r7_c0_rr0;
  wire [15:0] t0_r7_c1_rr0;
  wire [15:0] t0_r7_c1_rr1;
  wire [15:0] t0_r7_c1_rr2;
  wire [15:0] t0_r7_c1_rr3;
  wire [15:0] t0_r7_c1_rr4;
  wire [15:0] t0_r7_c1_rr5;
  wire [15:0] t0_r7_c1_rr6;
  wire [15:0] t0_r7_c1_rr7;
  wire [15:0] t0_r7_c1_rr8;
  wire [15:0] t0_r7_c1_rr9;
  wire [15:0] t1_r7_c1_rr0;
  wire [15:0] t1_r7_c1_rr1;
  wire [15:0] t1_r7_c1_rr2;
  wire [15:0] t1_r7_c1_rr3;
  wire [15:0] t1_r7_c1_rr4;
  wire [15:0] t2_r7_c1_rr0;
  wire [15:0] t2_r7_c1_rr1;
  wire [15:0] t2_r7_c1_rr2;
  wire [15:0] t3_r7_c1_rr0;
  wire [15:0] t3_r7_c1_rr1;
  wire [15:0] t4_r7_c1_rr0;
  wire [15:0] t0_r7_c2_rr0;
  wire [15:0] t0_r7_c2_rr1;
  wire [15:0] t0_r7_c2_rr2;
  wire [15:0] t0_r7_c2_rr3;
  wire [15:0] t0_r7_c2_rr4;
  wire [15:0] t0_r7_c2_rr5;
  wire [15:0] t0_r7_c2_rr6;
  wire [15:0] t0_r7_c2_rr7;
  wire [15:0] t0_r7_c2_rr8;
  wire [15:0] t0_r7_c2_rr9;
  wire [15:0] t1_r7_c2_rr0;
  wire [15:0] t1_r7_c2_rr1;
  wire [15:0] t1_r7_c2_rr2;
  wire [15:0] t1_r7_c2_rr3;
  wire [15:0] t1_r7_c2_rr4;
  wire [15:0] t2_r7_c2_rr0;
  wire [15:0] t2_r7_c2_rr1;
  wire [15:0] t2_r7_c2_rr2;
  wire [15:0] t3_r7_c2_rr0;
  wire [15:0] t3_r7_c2_rr1;
  wire [15:0] t4_r7_c2_rr0;
  wire [15:0] t0_r7_c3_rr0;
  wire [15:0] t0_r7_c3_rr1;
  wire [15:0] t0_r7_c3_rr2;
  wire [15:0] t0_r7_c3_rr3;
  wire [15:0] t0_r7_c3_rr4;
  wire [15:0] t0_r7_c3_rr5;
  wire [15:0] t0_r7_c3_rr6;
  wire [15:0] t0_r7_c3_rr7;
  wire [15:0] t0_r7_c3_rr8;
  wire [15:0] t0_r7_c3_rr9;
  wire [15:0] t1_r7_c3_rr0;
  wire [15:0] t1_r7_c3_rr1;
  wire [15:0] t1_r7_c3_rr2;
  wire [15:0] t1_r7_c3_rr3;
  wire [15:0] t1_r7_c3_rr4;
  wire [15:0] t2_r7_c3_rr0;
  wire [15:0] t2_r7_c3_rr1;
  wire [15:0] t2_r7_c3_rr2;
  wire [15:0] t3_r7_c3_rr0;
  wire [15:0] t3_r7_c3_rr1;
  wire [15:0] t4_r7_c3_rr0;
  wire [15:0] t0_r7_c4_rr0;
  wire [15:0] t0_r7_c4_rr1;
  wire [15:0] t0_r7_c4_rr2;
  wire [15:0] t0_r7_c4_rr3;
  wire [15:0] t0_r7_c4_rr4;
  wire [15:0] t0_r7_c4_rr5;
  wire [15:0] t0_r7_c4_rr6;
  wire [15:0] t0_r7_c4_rr7;
  wire [15:0] t0_r7_c4_rr8;
  wire [15:0] t0_r7_c4_rr9;
  wire [15:0] t1_r7_c4_rr0;
  wire [15:0] t1_r7_c4_rr1;
  wire [15:0] t1_r7_c4_rr2;
  wire [15:0] t1_r7_c4_rr3;
  wire [15:0] t1_r7_c4_rr4;
  wire [15:0] t2_r7_c4_rr0;
  wire [15:0] t2_r7_c4_rr1;
  wire [15:0] t2_r7_c4_rr2;
  wire [15:0] t3_r7_c4_rr0;
  wire [15:0] t3_r7_c4_rr1;
  wire [15:0] t4_r7_c4_rr0;
  wire [15:0] t0_r7_c5_rr0;
  wire [15:0] t0_r7_c5_rr1;
  wire [15:0] t0_r7_c5_rr2;
  wire [15:0] t0_r7_c5_rr3;
  wire [15:0] t0_r7_c5_rr4;
  wire [15:0] t0_r7_c5_rr5;
  wire [15:0] t0_r7_c5_rr6;
  wire [15:0] t0_r7_c5_rr7;
  wire [15:0] t0_r7_c5_rr8;
  wire [15:0] t0_r7_c5_rr9;
  wire [15:0] t1_r7_c5_rr0;
  wire [15:0] t1_r7_c5_rr1;
  wire [15:0] t1_r7_c5_rr2;
  wire [15:0] t1_r7_c5_rr3;
  wire [15:0] t1_r7_c5_rr4;
  wire [15:0] t2_r7_c5_rr0;
  wire [15:0] t2_r7_c5_rr1;
  wire [15:0] t2_r7_c5_rr2;
  wire [15:0] t3_r7_c5_rr0;
  wire [15:0] t3_r7_c5_rr1;
  wire [15:0] t4_r7_c5_rr0;
  wire [15:0] t0_r7_c6_rr0;
  wire [15:0] t0_r7_c6_rr1;
  wire [15:0] t0_r7_c6_rr2;
  wire [15:0] t0_r7_c6_rr3;
  wire [15:0] t0_r7_c6_rr4;
  wire [15:0] t0_r7_c6_rr5;
  wire [15:0] t0_r7_c6_rr6;
  wire [15:0] t0_r7_c6_rr7;
  wire [15:0] t0_r7_c6_rr8;
  wire [15:0] t0_r7_c6_rr9;
  wire [15:0] t1_r7_c6_rr0;
  wire [15:0] t1_r7_c6_rr1;
  wire [15:0] t1_r7_c6_rr2;
  wire [15:0] t1_r7_c6_rr3;
  wire [15:0] t1_r7_c6_rr4;
  wire [15:0] t2_r7_c6_rr0;
  wire [15:0] t2_r7_c6_rr1;
  wire [15:0] t2_r7_c6_rr2;
  wire [15:0] t3_r7_c6_rr0;
  wire [15:0] t3_r7_c6_rr1;
  wire [15:0] t4_r7_c6_rr0;
  wire [15:0] t0_r7_c7_rr0;
  wire [15:0] t0_r7_c7_rr1;
  wire [15:0] t0_r7_c7_rr2;
  wire [15:0] t0_r7_c7_rr3;
  wire [15:0] t0_r7_c7_rr4;
  wire [15:0] t0_r7_c7_rr5;
  wire [15:0] t0_r7_c7_rr6;
  wire [15:0] t0_r7_c7_rr7;
  wire [15:0] t0_r7_c7_rr8;
  wire [15:0] t0_r7_c7_rr9;
  wire [15:0] t1_r7_c7_rr0;
  wire [15:0] t1_r7_c7_rr1;
  wire [15:0] t1_r7_c7_rr2;
  wire [15:0] t1_r7_c7_rr3;
  wire [15:0] t1_r7_c7_rr4;
  wire [15:0] t2_r7_c7_rr0;
  wire [15:0] t2_r7_c7_rr1;
  wire [15:0] t2_r7_c7_rr2;
  wire [15:0] t3_r7_c7_rr0;
  wire [15:0] t3_r7_c7_rr1;
  wire [15:0] t4_r7_c7_rr0;
  wire [15:0] t0_r7_c8_rr0;
  wire [15:0] t0_r7_c8_rr1;
  wire [15:0] t0_r7_c8_rr2;
  wire [15:0] t0_r7_c8_rr3;
  wire [15:0] t0_r7_c8_rr4;
  wire [15:0] t0_r7_c8_rr5;
  wire [15:0] t0_r7_c8_rr6;
  wire [15:0] t0_r7_c8_rr7;
  wire [15:0] t0_r7_c8_rr8;
  wire [15:0] t0_r7_c8_rr9;
  wire [15:0] t1_r7_c8_rr0;
  wire [15:0] t1_r7_c8_rr1;
  wire [15:0] t1_r7_c8_rr2;
  wire [15:0] t1_r7_c8_rr3;
  wire [15:0] t1_r7_c8_rr4;
  wire [15:0] t2_r7_c8_rr0;
  wire [15:0] t2_r7_c8_rr1;
  wire [15:0] t2_r7_c8_rr2;
  wire [15:0] t3_r7_c8_rr0;
  wire [15:0] t3_r7_c8_rr1;
  wire [15:0] t4_r7_c8_rr0;
  wire [15:0] t0_r7_c9_rr0;
  wire [15:0] t0_r7_c9_rr1;
  wire [15:0] t0_r7_c9_rr2;
  wire [15:0] t0_r7_c9_rr3;
  wire [15:0] t0_r7_c9_rr4;
  wire [15:0] t0_r7_c9_rr5;
  wire [15:0] t0_r7_c9_rr6;
  wire [15:0] t0_r7_c9_rr7;
  wire [15:0] t0_r7_c9_rr8;
  wire [15:0] t0_r7_c9_rr9;
  wire [15:0] t1_r7_c9_rr0;
  wire [15:0] t1_r7_c9_rr1;
  wire [15:0] t1_r7_c9_rr2;
  wire [15:0] t1_r7_c9_rr3;
  wire [15:0] t1_r7_c9_rr4;
  wire [15:0] t2_r7_c9_rr0;
  wire [15:0] t2_r7_c9_rr1;
  wire [15:0] t2_r7_c9_rr2;
  wire [15:0] t3_r7_c9_rr0;
  wire [15:0] t3_r7_c9_rr1;
  wire [15:0] t4_r7_c9_rr0;
  wire [15:0] t0_r8_c0_rr0;
  wire [15:0] t0_r8_c0_rr1;
  wire [15:0] t0_r8_c0_rr2;
  wire [15:0] t0_r8_c0_rr3;
  wire [15:0] t0_r8_c0_rr4;
  wire [15:0] t0_r8_c0_rr5;
  wire [15:0] t0_r8_c0_rr6;
  wire [15:0] t0_r8_c0_rr7;
  wire [15:0] t0_r8_c0_rr8;
  wire [15:0] t0_r8_c0_rr9;
  wire [15:0] t1_r8_c0_rr0;
  wire [15:0] t1_r8_c0_rr1;
  wire [15:0] t1_r8_c0_rr2;
  wire [15:0] t1_r8_c0_rr3;
  wire [15:0] t1_r8_c0_rr4;
  wire [15:0] t2_r8_c0_rr0;
  wire [15:0] t2_r8_c0_rr1;
  wire [15:0] t2_r8_c0_rr2;
  wire [15:0] t3_r8_c0_rr0;
  wire [15:0] t3_r8_c0_rr1;
  wire [15:0] t4_r8_c0_rr0;
  wire [15:0] t0_r8_c1_rr0;
  wire [15:0] t0_r8_c1_rr1;
  wire [15:0] t0_r8_c1_rr2;
  wire [15:0] t0_r8_c1_rr3;
  wire [15:0] t0_r8_c1_rr4;
  wire [15:0] t0_r8_c1_rr5;
  wire [15:0] t0_r8_c1_rr6;
  wire [15:0] t0_r8_c1_rr7;
  wire [15:0] t0_r8_c1_rr8;
  wire [15:0] t0_r8_c1_rr9;
  wire [15:0] t1_r8_c1_rr0;
  wire [15:0] t1_r8_c1_rr1;
  wire [15:0] t1_r8_c1_rr2;
  wire [15:0] t1_r8_c1_rr3;
  wire [15:0] t1_r8_c1_rr4;
  wire [15:0] t2_r8_c1_rr0;
  wire [15:0] t2_r8_c1_rr1;
  wire [15:0] t2_r8_c1_rr2;
  wire [15:0] t3_r8_c1_rr0;
  wire [15:0] t3_r8_c1_rr1;
  wire [15:0] t4_r8_c1_rr0;
  wire [15:0] t0_r8_c2_rr0;
  wire [15:0] t0_r8_c2_rr1;
  wire [15:0] t0_r8_c2_rr2;
  wire [15:0] t0_r8_c2_rr3;
  wire [15:0] t0_r8_c2_rr4;
  wire [15:0] t0_r8_c2_rr5;
  wire [15:0] t0_r8_c2_rr6;
  wire [15:0] t0_r8_c2_rr7;
  wire [15:0] t0_r8_c2_rr8;
  wire [15:0] t0_r8_c2_rr9;
  wire [15:0] t1_r8_c2_rr0;
  wire [15:0] t1_r8_c2_rr1;
  wire [15:0] t1_r8_c2_rr2;
  wire [15:0] t1_r8_c2_rr3;
  wire [15:0] t1_r8_c2_rr4;
  wire [15:0] t2_r8_c2_rr0;
  wire [15:0] t2_r8_c2_rr1;
  wire [15:0] t2_r8_c2_rr2;
  wire [15:0] t3_r8_c2_rr0;
  wire [15:0] t3_r8_c2_rr1;
  wire [15:0] t4_r8_c2_rr0;
  wire [15:0] t0_r8_c3_rr0;
  wire [15:0] t0_r8_c3_rr1;
  wire [15:0] t0_r8_c3_rr2;
  wire [15:0] t0_r8_c3_rr3;
  wire [15:0] t0_r8_c3_rr4;
  wire [15:0] t0_r8_c3_rr5;
  wire [15:0] t0_r8_c3_rr6;
  wire [15:0] t0_r8_c3_rr7;
  wire [15:0] t0_r8_c3_rr8;
  wire [15:0] t0_r8_c3_rr9;
  wire [15:0] t1_r8_c3_rr0;
  wire [15:0] t1_r8_c3_rr1;
  wire [15:0] t1_r8_c3_rr2;
  wire [15:0] t1_r8_c3_rr3;
  wire [15:0] t1_r8_c3_rr4;
  wire [15:0] t2_r8_c3_rr0;
  wire [15:0] t2_r8_c3_rr1;
  wire [15:0] t2_r8_c3_rr2;
  wire [15:0] t3_r8_c3_rr0;
  wire [15:0] t3_r8_c3_rr1;
  wire [15:0] t4_r8_c3_rr0;
  wire [15:0] t0_r8_c4_rr0;
  wire [15:0] t0_r8_c4_rr1;
  wire [15:0] t0_r8_c4_rr2;
  wire [15:0] t0_r8_c4_rr3;
  wire [15:0] t0_r8_c4_rr4;
  wire [15:0] t0_r8_c4_rr5;
  wire [15:0] t0_r8_c4_rr6;
  wire [15:0] t0_r8_c4_rr7;
  wire [15:0] t0_r8_c4_rr8;
  wire [15:0] t0_r8_c4_rr9;
  wire [15:0] t1_r8_c4_rr0;
  wire [15:0] t1_r8_c4_rr1;
  wire [15:0] t1_r8_c4_rr2;
  wire [15:0] t1_r8_c4_rr3;
  wire [15:0] t1_r8_c4_rr4;
  wire [15:0] t2_r8_c4_rr0;
  wire [15:0] t2_r8_c4_rr1;
  wire [15:0] t2_r8_c4_rr2;
  wire [15:0] t3_r8_c4_rr0;
  wire [15:0] t3_r8_c4_rr1;
  wire [15:0] t4_r8_c4_rr0;
  wire [15:0] t0_r8_c5_rr0;
  wire [15:0] t0_r8_c5_rr1;
  wire [15:0] t0_r8_c5_rr2;
  wire [15:0] t0_r8_c5_rr3;
  wire [15:0] t0_r8_c5_rr4;
  wire [15:0] t0_r8_c5_rr5;
  wire [15:0] t0_r8_c5_rr6;
  wire [15:0] t0_r8_c5_rr7;
  wire [15:0] t0_r8_c5_rr8;
  wire [15:0] t0_r8_c5_rr9;
  wire [15:0] t1_r8_c5_rr0;
  wire [15:0] t1_r8_c5_rr1;
  wire [15:0] t1_r8_c5_rr2;
  wire [15:0] t1_r8_c5_rr3;
  wire [15:0] t1_r8_c5_rr4;
  wire [15:0] t2_r8_c5_rr0;
  wire [15:0] t2_r8_c5_rr1;
  wire [15:0] t2_r8_c5_rr2;
  wire [15:0] t3_r8_c5_rr0;
  wire [15:0] t3_r8_c5_rr1;
  wire [15:0] t4_r8_c5_rr0;
  wire [15:0] t0_r8_c6_rr0;
  wire [15:0] t0_r8_c6_rr1;
  wire [15:0] t0_r8_c6_rr2;
  wire [15:0] t0_r8_c6_rr3;
  wire [15:0] t0_r8_c6_rr4;
  wire [15:0] t0_r8_c6_rr5;
  wire [15:0] t0_r8_c6_rr6;
  wire [15:0] t0_r8_c6_rr7;
  wire [15:0] t0_r8_c6_rr8;
  wire [15:0] t0_r8_c6_rr9;
  wire [15:0] t1_r8_c6_rr0;
  wire [15:0] t1_r8_c6_rr1;
  wire [15:0] t1_r8_c6_rr2;
  wire [15:0] t1_r8_c6_rr3;
  wire [15:0] t1_r8_c6_rr4;
  wire [15:0] t2_r8_c6_rr0;
  wire [15:0] t2_r8_c6_rr1;
  wire [15:0] t2_r8_c6_rr2;
  wire [15:0] t3_r8_c6_rr0;
  wire [15:0] t3_r8_c6_rr1;
  wire [15:0] t4_r8_c6_rr0;
  wire [15:0] t0_r8_c7_rr0;
  wire [15:0] t0_r8_c7_rr1;
  wire [15:0] t0_r8_c7_rr2;
  wire [15:0] t0_r8_c7_rr3;
  wire [15:0] t0_r8_c7_rr4;
  wire [15:0] t0_r8_c7_rr5;
  wire [15:0] t0_r8_c7_rr6;
  wire [15:0] t0_r8_c7_rr7;
  wire [15:0] t0_r8_c7_rr8;
  wire [15:0] t0_r8_c7_rr9;
  wire [15:0] t1_r8_c7_rr0;
  wire [15:0] t1_r8_c7_rr1;
  wire [15:0] t1_r8_c7_rr2;
  wire [15:0] t1_r8_c7_rr3;
  wire [15:0] t1_r8_c7_rr4;
  wire [15:0] t2_r8_c7_rr0;
  wire [15:0] t2_r8_c7_rr1;
  wire [15:0] t2_r8_c7_rr2;
  wire [15:0] t3_r8_c7_rr0;
  wire [15:0] t3_r8_c7_rr1;
  wire [15:0] t4_r8_c7_rr0;
  wire [15:0] t0_r8_c8_rr0;
  wire [15:0] t0_r8_c8_rr1;
  wire [15:0] t0_r8_c8_rr2;
  wire [15:0] t0_r8_c8_rr3;
  wire [15:0] t0_r8_c8_rr4;
  wire [15:0] t0_r8_c8_rr5;
  wire [15:0] t0_r8_c8_rr6;
  wire [15:0] t0_r8_c8_rr7;
  wire [15:0] t0_r8_c8_rr8;
  wire [15:0] t0_r8_c8_rr9;
  wire [15:0] t1_r8_c8_rr0;
  wire [15:0] t1_r8_c8_rr1;
  wire [15:0] t1_r8_c8_rr2;
  wire [15:0] t1_r8_c8_rr3;
  wire [15:0] t1_r8_c8_rr4;
  wire [15:0] t2_r8_c8_rr0;
  wire [15:0] t2_r8_c8_rr1;
  wire [15:0] t2_r8_c8_rr2;
  wire [15:0] t3_r8_c8_rr0;
  wire [15:0] t3_r8_c8_rr1;
  wire [15:0] t4_r8_c8_rr0;
  wire [15:0] t0_r8_c9_rr0;
  wire [15:0] t0_r8_c9_rr1;
  wire [15:0] t0_r8_c9_rr2;
  wire [15:0] t0_r8_c9_rr3;
  wire [15:0] t0_r8_c9_rr4;
  wire [15:0] t0_r8_c9_rr5;
  wire [15:0] t0_r8_c9_rr6;
  wire [15:0] t0_r8_c9_rr7;
  wire [15:0] t0_r8_c9_rr8;
  wire [15:0] t0_r8_c9_rr9;
  wire [15:0] t1_r8_c9_rr0;
  wire [15:0] t1_r8_c9_rr1;
  wire [15:0] t1_r8_c9_rr2;
  wire [15:0] t1_r8_c9_rr3;
  wire [15:0] t1_r8_c9_rr4;
  wire [15:0] t2_r8_c9_rr0;
  wire [15:0] t2_r8_c9_rr1;
  wire [15:0] t2_r8_c9_rr2;
  wire [15:0] t3_r8_c9_rr0;
  wire [15:0] t3_r8_c9_rr1;
  wire [15:0] t4_r8_c9_rr0;
  wire [15:0] t0_r9_c0_rr0;
  wire [15:0] t0_r9_c0_rr1;
  wire [15:0] t0_r9_c0_rr2;
  wire [15:0] t0_r9_c0_rr3;
  wire [15:0] t0_r9_c0_rr4;
  wire [15:0] t0_r9_c0_rr5;
  wire [15:0] t0_r9_c0_rr6;
  wire [15:0] t0_r9_c0_rr7;
  wire [15:0] t0_r9_c0_rr8;
  wire [15:0] t0_r9_c0_rr9;
  wire [15:0] t1_r9_c0_rr0;
  wire [15:0] t1_r9_c0_rr1;
  wire [15:0] t1_r9_c0_rr2;
  wire [15:0] t1_r9_c0_rr3;
  wire [15:0] t1_r9_c0_rr4;
  wire [15:0] t2_r9_c0_rr0;
  wire [15:0] t2_r9_c0_rr1;
  wire [15:0] t2_r9_c0_rr2;
  wire [15:0] t3_r9_c0_rr0;
  wire [15:0] t3_r9_c0_rr1;
  wire [15:0] t4_r9_c0_rr0;
  wire [15:0] t0_r9_c1_rr0;
  wire [15:0] t0_r9_c1_rr1;
  wire [15:0] t0_r9_c1_rr2;
  wire [15:0] t0_r9_c1_rr3;
  wire [15:0] t0_r9_c1_rr4;
  wire [15:0] t0_r9_c1_rr5;
  wire [15:0] t0_r9_c1_rr6;
  wire [15:0] t0_r9_c1_rr7;
  wire [15:0] t0_r9_c1_rr8;
  wire [15:0] t0_r9_c1_rr9;
  wire [15:0] t1_r9_c1_rr0;
  wire [15:0] t1_r9_c1_rr1;
  wire [15:0] t1_r9_c1_rr2;
  wire [15:0] t1_r9_c1_rr3;
  wire [15:0] t1_r9_c1_rr4;
  wire [15:0] t2_r9_c1_rr0;
  wire [15:0] t2_r9_c1_rr1;
  wire [15:0] t2_r9_c1_rr2;
  wire [15:0] t3_r9_c1_rr0;
  wire [15:0] t3_r9_c1_rr1;
  wire [15:0] t4_r9_c1_rr0;
  wire [15:0] t0_r9_c2_rr0;
  wire [15:0] t0_r9_c2_rr1;
  wire [15:0] t0_r9_c2_rr2;
  wire [15:0] t0_r9_c2_rr3;
  wire [15:0] t0_r9_c2_rr4;
  wire [15:0] t0_r9_c2_rr5;
  wire [15:0] t0_r9_c2_rr6;
  wire [15:0] t0_r9_c2_rr7;
  wire [15:0] t0_r9_c2_rr8;
  wire [15:0] t0_r9_c2_rr9;
  wire [15:0] t1_r9_c2_rr0;
  wire [15:0] t1_r9_c2_rr1;
  wire [15:0] t1_r9_c2_rr2;
  wire [15:0] t1_r9_c2_rr3;
  wire [15:0] t1_r9_c2_rr4;
  wire [15:0] t2_r9_c2_rr0;
  wire [15:0] t2_r9_c2_rr1;
  wire [15:0] t2_r9_c2_rr2;
  wire [15:0] t3_r9_c2_rr0;
  wire [15:0] t3_r9_c2_rr1;
  wire [15:0] t4_r9_c2_rr0;
  wire [15:0] t0_r9_c3_rr0;
  wire [15:0] t0_r9_c3_rr1;
  wire [15:0] t0_r9_c3_rr2;
  wire [15:0] t0_r9_c3_rr3;
  wire [15:0] t0_r9_c3_rr4;
  wire [15:0] t0_r9_c3_rr5;
  wire [15:0] t0_r9_c3_rr6;
  wire [15:0] t0_r9_c3_rr7;
  wire [15:0] t0_r9_c3_rr8;
  wire [15:0] t0_r9_c3_rr9;
  wire [15:0] t1_r9_c3_rr0;
  wire [15:0] t1_r9_c3_rr1;
  wire [15:0] t1_r9_c3_rr2;
  wire [15:0] t1_r9_c3_rr3;
  wire [15:0] t1_r9_c3_rr4;
  wire [15:0] t2_r9_c3_rr0;
  wire [15:0] t2_r9_c3_rr1;
  wire [15:0] t2_r9_c3_rr2;
  wire [15:0] t3_r9_c3_rr0;
  wire [15:0] t3_r9_c3_rr1;
  wire [15:0] t4_r9_c3_rr0;
  wire [15:0] t0_r9_c4_rr0;
  wire [15:0] t0_r9_c4_rr1;
  wire [15:0] t0_r9_c4_rr2;
  wire [15:0] t0_r9_c4_rr3;
  wire [15:0] t0_r9_c4_rr4;
  wire [15:0] t0_r9_c4_rr5;
  wire [15:0] t0_r9_c4_rr6;
  wire [15:0] t0_r9_c4_rr7;
  wire [15:0] t0_r9_c4_rr8;
  wire [15:0] t0_r9_c4_rr9;
  wire [15:0] t1_r9_c4_rr0;
  wire [15:0] t1_r9_c4_rr1;
  wire [15:0] t1_r9_c4_rr2;
  wire [15:0] t1_r9_c4_rr3;
  wire [15:0] t1_r9_c4_rr4;
  wire [15:0] t2_r9_c4_rr0;
  wire [15:0] t2_r9_c4_rr1;
  wire [15:0] t2_r9_c4_rr2;
  wire [15:0] t3_r9_c4_rr0;
  wire [15:0] t3_r9_c4_rr1;
  wire [15:0] t4_r9_c4_rr0;
  wire [15:0] t0_r9_c5_rr0;
  wire [15:0] t0_r9_c5_rr1;
  wire [15:0] t0_r9_c5_rr2;
  wire [15:0] t0_r9_c5_rr3;
  wire [15:0] t0_r9_c5_rr4;
  wire [15:0] t0_r9_c5_rr5;
  wire [15:0] t0_r9_c5_rr6;
  wire [15:0] t0_r9_c5_rr7;
  wire [15:0] t0_r9_c5_rr8;
  wire [15:0] t0_r9_c5_rr9;
  wire [15:0] t1_r9_c5_rr0;
  wire [15:0] t1_r9_c5_rr1;
  wire [15:0] t1_r9_c5_rr2;
  wire [15:0] t1_r9_c5_rr3;
  wire [15:0] t1_r9_c5_rr4;
  wire [15:0] t2_r9_c5_rr0;
  wire [15:0] t2_r9_c5_rr1;
  wire [15:0] t2_r9_c5_rr2;
  wire [15:0] t3_r9_c5_rr0;
  wire [15:0] t3_r9_c5_rr1;
  wire [15:0] t4_r9_c5_rr0;
  wire [15:0] t0_r9_c6_rr0;
  wire [15:0] t0_r9_c6_rr1;
  wire [15:0] t0_r9_c6_rr2;
  wire [15:0] t0_r9_c6_rr3;
  wire [15:0] t0_r9_c6_rr4;
  wire [15:0] t0_r9_c6_rr5;
  wire [15:0] t0_r9_c6_rr6;
  wire [15:0] t0_r9_c6_rr7;
  wire [15:0] t0_r9_c6_rr8;
  wire [15:0] t0_r9_c6_rr9;
  wire [15:0] t1_r9_c6_rr0;
  wire [15:0] t1_r9_c6_rr1;
  wire [15:0] t1_r9_c6_rr2;
  wire [15:0] t1_r9_c6_rr3;
  wire [15:0] t1_r9_c6_rr4;
  wire [15:0] t2_r9_c6_rr0;
  wire [15:0] t2_r9_c6_rr1;
  wire [15:0] t2_r9_c6_rr2;
  wire [15:0] t3_r9_c6_rr0;
  wire [15:0] t3_r9_c6_rr1;
  wire [15:0] t4_r9_c6_rr0;
  wire [15:0] t0_r9_c7_rr0;
  wire [15:0] t0_r9_c7_rr1;
  wire [15:0] t0_r9_c7_rr2;
  wire [15:0] t0_r9_c7_rr3;
  wire [15:0] t0_r9_c7_rr4;
  wire [15:0] t0_r9_c7_rr5;
  wire [15:0] t0_r9_c7_rr6;
  wire [15:0] t0_r9_c7_rr7;
  wire [15:0] t0_r9_c7_rr8;
  wire [15:0] t0_r9_c7_rr9;
  wire [15:0] t1_r9_c7_rr0;
  wire [15:0] t1_r9_c7_rr1;
  wire [15:0] t1_r9_c7_rr2;
  wire [15:0] t1_r9_c7_rr3;
  wire [15:0] t1_r9_c7_rr4;
  wire [15:0] t2_r9_c7_rr0;
  wire [15:0] t2_r9_c7_rr1;
  wire [15:0] t2_r9_c7_rr2;
  wire [15:0] t3_r9_c7_rr0;
  wire [15:0] t3_r9_c7_rr1;
  wire [15:0] t4_r9_c7_rr0;
  wire [15:0] t0_r9_c8_rr0;
  wire [15:0] t0_r9_c8_rr1;
  wire [15:0] t0_r9_c8_rr2;
  wire [15:0] t0_r9_c8_rr3;
  wire [15:0] t0_r9_c8_rr4;
  wire [15:0] t0_r9_c8_rr5;
  wire [15:0] t0_r9_c8_rr6;
  wire [15:0] t0_r9_c8_rr7;
  wire [15:0] t0_r9_c8_rr8;
  wire [15:0] t0_r9_c8_rr9;
  wire [15:0] t1_r9_c8_rr0;
  wire [15:0] t1_r9_c8_rr1;
  wire [15:0] t1_r9_c8_rr2;
  wire [15:0] t1_r9_c8_rr3;
  wire [15:0] t1_r9_c8_rr4;
  wire [15:0] t2_r9_c8_rr0;
  wire [15:0] t2_r9_c8_rr1;
  wire [15:0] t2_r9_c8_rr2;
  wire [15:0] t3_r9_c8_rr0;
  wire [15:0] t3_r9_c8_rr1;
  wire [15:0] t4_r9_c8_rr0;
  wire [15:0] t0_r9_c9_rr0;
  wire [15:0] t0_r9_c9_rr1;
  wire [15:0] t0_r9_c9_rr2;
  wire [15:0] t0_r9_c9_rr3;
  wire [15:0] t0_r9_c9_rr4;
  wire [15:0] t0_r9_c9_rr5;
  wire [15:0] t0_r9_c9_rr6;
  wire [15:0] t0_r9_c9_rr7;
  wire [15:0] t0_r9_c9_rr8;
  wire [15:0] t0_r9_c9_rr9;
  wire [15:0] t1_r9_c9_rr0;
  wire [15:0] t1_r9_c9_rr1;
  wire [15:0] t1_r9_c9_rr2;
  wire [15:0] t1_r9_c9_rr3;
  wire [15:0] t1_r9_c9_rr4;
  wire [15:0] t2_r9_c9_rr0;
  wire [15:0] t2_r9_c9_rr1;
  wire [15:0] t2_r9_c9_rr2;
  wire [15:0] t3_r9_c9_rr0;
  wire [15:0] t3_r9_c9_rr1;
  wire [15:0] t4_r9_c9_rr0;

  assign t0_r0_c0_rr0 = a_0_0 * b_0_0;
  assign t0_r0_c0_rr1 = a_0_1 * b_1_0;
  assign t0_r0_c0_rr2 = a_0_2 * b_2_0;
  assign t0_r0_c0_rr3 = a_0_3 * b_3_0;
  assign t0_r0_c0_rr4 = a_0_4 * b_4_0;
  assign t0_r0_c0_rr5 = a_0_5 * b_5_0;
  assign t0_r0_c0_rr6 = a_0_6 * b_6_0;
  assign t0_r0_c0_rr7 = a_0_7 * b_7_0;
  assign t0_r0_c0_rr8 = a_0_8 * b_8_0;
  assign t0_r0_c0_rr9 = a_0_9 * b_9_0;
  assign t1_r0_c0_rr0 = t0_r0_c0_rr0 + t0_r0_c0_rr1;
  assign t1_r0_c0_rr1 = t0_r0_c0_rr2 + t0_r0_c0_rr3;
  assign t1_r0_c0_rr2 = t0_r0_c0_rr4 + t0_r0_c0_rr5;
  assign t1_r0_c0_rr3 = t0_r0_c0_rr6 + t0_r0_c0_rr7;
  assign t1_r0_c0_rr4 = t0_r0_c0_rr8 + t0_r0_c0_rr9;

  assign t2_r0_c0_rr0 = t1_r0_c0_rr0 + t1_r0_c0_rr1;
  assign t2_r0_c0_rr1 = t1_r0_c0_rr2 + t1_r0_c0_rr3;
  assign t2_r0_c0_rr2 = t1_r0_c0_rr4;

  assign t3_r0_c0_rr0 = t2_r0_c0_rr0 + t2_r0_c0_rr1;
  assign t3_r0_c0_rr1 = t2_r0_c0_rr2;

  assign t4_r0_c0_rr0 = t3_r0_c0_rr0 + t3_r0_c0_rr1;

  assign c_0_0 = t4_r0_c0_rr0;
  assign t0_r0_c1_rr0 = a_0_0 * b_0_1;
  assign t0_r0_c1_rr1 = a_0_1 * b_1_1;
  assign t0_r0_c1_rr2 = a_0_2 * b_2_1;
  assign t0_r0_c1_rr3 = a_0_3 * b_3_1;
  assign t0_r0_c1_rr4 = a_0_4 * b_4_1;
  assign t0_r0_c1_rr5 = a_0_5 * b_5_1;
  assign t0_r0_c1_rr6 = a_0_6 * b_6_1;
  assign t0_r0_c1_rr7 = a_0_7 * b_7_1;
  assign t0_r0_c1_rr8 = a_0_8 * b_8_1;
  assign t0_r0_c1_rr9 = a_0_9 * b_9_1;
  assign t1_r0_c1_rr0 = t0_r0_c1_rr0 + t0_r0_c1_rr1;
  assign t1_r0_c1_rr1 = t0_r0_c1_rr2 + t0_r0_c1_rr3;
  assign t1_r0_c1_rr2 = t0_r0_c1_rr4 + t0_r0_c1_rr5;
  assign t1_r0_c1_rr3 = t0_r0_c1_rr6 + t0_r0_c1_rr7;
  assign t1_r0_c1_rr4 = t0_r0_c1_rr8 + t0_r0_c1_rr9;

  assign t2_r0_c1_rr0 = t1_r0_c1_rr0 + t1_r0_c1_rr1;
  assign t2_r0_c1_rr1 = t1_r0_c1_rr2 + t1_r0_c1_rr3;
  assign t2_r0_c1_rr2 = t1_r0_c1_rr4;

  assign t3_r0_c1_rr0 = t2_r0_c1_rr0 + t2_r0_c1_rr1;
  assign t3_r0_c1_rr1 = t2_r0_c1_rr2;

  assign t4_r0_c1_rr0 = t3_r0_c1_rr0 + t3_r0_c1_rr1;

  assign c_0_1 = t4_r0_c1_rr0;
  assign t0_r0_c2_rr0 = a_0_0 * b_0_2;
  assign t0_r0_c2_rr1 = a_0_1 * b_1_2;
  assign t0_r0_c2_rr2 = a_0_2 * b_2_2;
  assign t0_r0_c2_rr3 = a_0_3 * b_3_2;
  assign t0_r0_c2_rr4 = a_0_4 * b_4_2;
  assign t0_r0_c2_rr5 = a_0_5 * b_5_2;
  assign t0_r0_c2_rr6 = a_0_6 * b_6_2;
  assign t0_r0_c2_rr7 = a_0_7 * b_7_2;
  assign t0_r0_c2_rr8 = a_0_8 * b_8_2;
  assign t0_r0_c2_rr9 = a_0_9 * b_9_2;
  assign t1_r0_c2_rr0 = t0_r0_c2_rr0 + t0_r0_c2_rr1;
  assign t1_r0_c2_rr1 = t0_r0_c2_rr2 + t0_r0_c2_rr3;
  assign t1_r0_c2_rr2 = t0_r0_c2_rr4 + t0_r0_c2_rr5;
  assign t1_r0_c2_rr3 = t0_r0_c2_rr6 + t0_r0_c2_rr7;
  assign t1_r0_c2_rr4 = t0_r0_c2_rr8 + t0_r0_c2_rr9;

  assign t2_r0_c2_rr0 = t1_r0_c2_rr0 + t1_r0_c2_rr1;
  assign t2_r0_c2_rr1 = t1_r0_c2_rr2 + t1_r0_c2_rr3;
  assign t2_r0_c2_rr2 = t1_r0_c2_rr4;

  assign t3_r0_c2_rr0 = t2_r0_c2_rr0 + t2_r0_c2_rr1;
  assign t3_r0_c2_rr1 = t2_r0_c2_rr2;

  assign t4_r0_c2_rr0 = t3_r0_c2_rr0 + t3_r0_c2_rr1;

  assign c_0_2 = t4_r0_c2_rr0;
  assign t0_r0_c3_rr0 = a_0_0 * b_0_3;
  assign t0_r0_c3_rr1 = a_0_1 * b_1_3;
  assign t0_r0_c3_rr2 = a_0_2 * b_2_3;
  assign t0_r0_c3_rr3 = a_0_3 * b_3_3;
  assign t0_r0_c3_rr4 = a_0_4 * b_4_3;
  assign t0_r0_c3_rr5 = a_0_5 * b_5_3;
  assign t0_r0_c3_rr6 = a_0_6 * b_6_3;
  assign t0_r0_c3_rr7 = a_0_7 * b_7_3;
  assign t0_r0_c3_rr8 = a_0_8 * b_8_3;
  assign t0_r0_c3_rr9 = a_0_9 * b_9_3;
  assign t1_r0_c3_rr0 = t0_r0_c3_rr0 + t0_r0_c3_rr1;
  assign t1_r0_c3_rr1 = t0_r0_c3_rr2 + t0_r0_c3_rr3;
  assign t1_r0_c3_rr2 = t0_r0_c3_rr4 + t0_r0_c3_rr5;
  assign t1_r0_c3_rr3 = t0_r0_c3_rr6 + t0_r0_c3_rr7;
  assign t1_r0_c3_rr4 = t0_r0_c3_rr8 + t0_r0_c3_rr9;

  assign t2_r0_c3_rr0 = t1_r0_c3_rr0 + t1_r0_c3_rr1;
  assign t2_r0_c3_rr1 = t1_r0_c3_rr2 + t1_r0_c3_rr3;
  assign t2_r0_c3_rr2 = t1_r0_c3_rr4;

  assign t3_r0_c3_rr0 = t2_r0_c3_rr0 + t2_r0_c3_rr1;
  assign t3_r0_c3_rr1 = t2_r0_c3_rr2;

  assign t4_r0_c3_rr0 = t3_r0_c3_rr0 + t3_r0_c3_rr1;

  assign c_0_3 = t4_r0_c3_rr0;
  assign t0_r0_c4_rr0 = a_0_0 * b_0_4;
  assign t0_r0_c4_rr1 = a_0_1 * b_1_4;
  assign t0_r0_c4_rr2 = a_0_2 * b_2_4;
  assign t0_r0_c4_rr3 = a_0_3 * b_3_4;
  assign t0_r0_c4_rr4 = a_0_4 * b_4_4;
  assign t0_r0_c4_rr5 = a_0_5 * b_5_4;
  assign t0_r0_c4_rr6 = a_0_6 * b_6_4;
  assign t0_r0_c4_rr7 = a_0_7 * b_7_4;
  assign t0_r0_c4_rr8 = a_0_8 * b_8_4;
  assign t0_r0_c4_rr9 = a_0_9 * b_9_4;
  assign t1_r0_c4_rr0 = t0_r0_c4_rr0 + t0_r0_c4_rr1;
  assign t1_r0_c4_rr1 = t0_r0_c4_rr2 + t0_r0_c4_rr3;
  assign t1_r0_c4_rr2 = t0_r0_c4_rr4 + t0_r0_c4_rr5;
  assign t1_r0_c4_rr3 = t0_r0_c4_rr6 + t0_r0_c4_rr7;
  assign t1_r0_c4_rr4 = t0_r0_c4_rr8 + t0_r0_c4_rr9;

  assign t2_r0_c4_rr0 = t1_r0_c4_rr0 + t1_r0_c4_rr1;
  assign t2_r0_c4_rr1 = t1_r0_c4_rr2 + t1_r0_c4_rr3;
  assign t2_r0_c4_rr2 = t1_r0_c4_rr4;

  assign t3_r0_c4_rr0 = t2_r0_c4_rr0 + t2_r0_c4_rr1;
  assign t3_r0_c4_rr1 = t2_r0_c4_rr2;

  assign t4_r0_c4_rr0 = t3_r0_c4_rr0 + t3_r0_c4_rr1;

  assign c_0_4 = t4_r0_c4_rr0;
  assign t0_r0_c5_rr0 = a_0_0 * b_0_5;
  assign t0_r0_c5_rr1 = a_0_1 * b_1_5;
  assign t0_r0_c5_rr2 = a_0_2 * b_2_5;
  assign t0_r0_c5_rr3 = a_0_3 * b_3_5;
  assign t0_r0_c5_rr4 = a_0_4 * b_4_5;
  assign t0_r0_c5_rr5 = a_0_5 * b_5_5;
  assign t0_r0_c5_rr6 = a_0_6 * b_6_5;
  assign t0_r0_c5_rr7 = a_0_7 * b_7_5;
  assign t0_r0_c5_rr8 = a_0_8 * b_8_5;
  assign t0_r0_c5_rr9 = a_0_9 * b_9_5;
  assign t1_r0_c5_rr0 = t0_r0_c5_rr0 + t0_r0_c5_rr1;
  assign t1_r0_c5_rr1 = t0_r0_c5_rr2 + t0_r0_c5_rr3;
  assign t1_r0_c5_rr2 = t0_r0_c5_rr4 + t0_r0_c5_rr5;
  assign t1_r0_c5_rr3 = t0_r0_c5_rr6 + t0_r0_c5_rr7;
  assign t1_r0_c5_rr4 = t0_r0_c5_rr8 + t0_r0_c5_rr9;

  assign t2_r0_c5_rr0 = t1_r0_c5_rr0 + t1_r0_c5_rr1;
  assign t2_r0_c5_rr1 = t1_r0_c5_rr2 + t1_r0_c5_rr3;
  assign t2_r0_c5_rr2 = t1_r0_c5_rr4;

  assign t3_r0_c5_rr0 = t2_r0_c5_rr0 + t2_r0_c5_rr1;
  assign t3_r0_c5_rr1 = t2_r0_c5_rr2;

  assign t4_r0_c5_rr0 = t3_r0_c5_rr0 + t3_r0_c5_rr1;

  assign c_0_5 = t4_r0_c5_rr0;
  assign t0_r0_c6_rr0 = a_0_0 * b_0_6;
  assign t0_r0_c6_rr1 = a_0_1 * b_1_6;
  assign t0_r0_c6_rr2 = a_0_2 * b_2_6;
  assign t0_r0_c6_rr3 = a_0_3 * b_3_6;
  assign t0_r0_c6_rr4 = a_0_4 * b_4_6;
  assign t0_r0_c6_rr5 = a_0_5 * b_5_6;
  assign t0_r0_c6_rr6 = a_0_6 * b_6_6;
  assign t0_r0_c6_rr7 = a_0_7 * b_7_6;
  assign t0_r0_c6_rr8 = a_0_8 * b_8_6;
  assign t0_r0_c6_rr9 = a_0_9 * b_9_6;
  assign t1_r0_c6_rr0 = t0_r0_c6_rr0 + t0_r0_c6_rr1;
  assign t1_r0_c6_rr1 = t0_r0_c6_rr2 + t0_r0_c6_rr3;
  assign t1_r0_c6_rr2 = t0_r0_c6_rr4 + t0_r0_c6_rr5;
  assign t1_r0_c6_rr3 = t0_r0_c6_rr6 + t0_r0_c6_rr7;
  assign t1_r0_c6_rr4 = t0_r0_c6_rr8 + t0_r0_c6_rr9;

  assign t2_r0_c6_rr0 = t1_r0_c6_rr0 + t1_r0_c6_rr1;
  assign t2_r0_c6_rr1 = t1_r0_c6_rr2 + t1_r0_c6_rr3;
  assign t2_r0_c6_rr2 = t1_r0_c6_rr4;

  assign t3_r0_c6_rr0 = t2_r0_c6_rr0 + t2_r0_c6_rr1;
  assign t3_r0_c6_rr1 = t2_r0_c6_rr2;

  assign t4_r0_c6_rr0 = t3_r0_c6_rr0 + t3_r0_c6_rr1;

  assign c_0_6 = t4_r0_c6_rr0;
  assign t0_r0_c7_rr0 = a_0_0 * b_0_7;
  assign t0_r0_c7_rr1 = a_0_1 * b_1_7;
  assign t0_r0_c7_rr2 = a_0_2 * b_2_7;
  assign t0_r0_c7_rr3 = a_0_3 * b_3_7;
  assign t0_r0_c7_rr4 = a_0_4 * b_4_7;
  assign t0_r0_c7_rr5 = a_0_5 * b_5_7;
  assign t0_r0_c7_rr6 = a_0_6 * b_6_7;
  assign t0_r0_c7_rr7 = a_0_7 * b_7_7;
  assign t0_r0_c7_rr8 = a_0_8 * b_8_7;
  assign t0_r0_c7_rr9 = a_0_9 * b_9_7;
  assign t1_r0_c7_rr0 = t0_r0_c7_rr0 + t0_r0_c7_rr1;
  assign t1_r0_c7_rr1 = t0_r0_c7_rr2 + t0_r0_c7_rr3;
  assign t1_r0_c7_rr2 = t0_r0_c7_rr4 + t0_r0_c7_rr5;
  assign t1_r0_c7_rr3 = t0_r0_c7_rr6 + t0_r0_c7_rr7;
  assign t1_r0_c7_rr4 = t0_r0_c7_rr8 + t0_r0_c7_rr9;

  assign t2_r0_c7_rr0 = t1_r0_c7_rr0 + t1_r0_c7_rr1;
  assign t2_r0_c7_rr1 = t1_r0_c7_rr2 + t1_r0_c7_rr3;
  assign t2_r0_c7_rr2 = t1_r0_c7_rr4;

  assign t3_r0_c7_rr0 = t2_r0_c7_rr0 + t2_r0_c7_rr1;
  assign t3_r0_c7_rr1 = t2_r0_c7_rr2;

  assign t4_r0_c7_rr0 = t3_r0_c7_rr0 + t3_r0_c7_rr1;

  assign c_0_7 = t4_r0_c7_rr0;
  assign t0_r0_c8_rr0 = a_0_0 * b_0_8;
  assign t0_r0_c8_rr1 = a_0_1 * b_1_8;
  assign t0_r0_c8_rr2 = a_0_2 * b_2_8;
  assign t0_r0_c8_rr3 = a_0_3 * b_3_8;
  assign t0_r0_c8_rr4 = a_0_4 * b_4_8;
  assign t0_r0_c8_rr5 = a_0_5 * b_5_8;
  assign t0_r0_c8_rr6 = a_0_6 * b_6_8;
  assign t0_r0_c8_rr7 = a_0_7 * b_7_8;
  assign t0_r0_c8_rr8 = a_0_8 * b_8_8;
  assign t0_r0_c8_rr9 = a_0_9 * b_9_8;
  assign t1_r0_c8_rr0 = t0_r0_c8_rr0 + t0_r0_c8_rr1;
  assign t1_r0_c8_rr1 = t0_r0_c8_rr2 + t0_r0_c8_rr3;
  assign t1_r0_c8_rr2 = t0_r0_c8_rr4 + t0_r0_c8_rr5;
  assign t1_r0_c8_rr3 = t0_r0_c8_rr6 + t0_r0_c8_rr7;
  assign t1_r0_c8_rr4 = t0_r0_c8_rr8 + t0_r0_c8_rr9;

  assign t2_r0_c8_rr0 = t1_r0_c8_rr0 + t1_r0_c8_rr1;
  assign t2_r0_c8_rr1 = t1_r0_c8_rr2 + t1_r0_c8_rr3;
  assign t2_r0_c8_rr2 = t1_r0_c8_rr4;

  assign t3_r0_c8_rr0 = t2_r0_c8_rr0 + t2_r0_c8_rr1;
  assign t3_r0_c8_rr1 = t2_r0_c8_rr2;

  assign t4_r0_c8_rr0 = t3_r0_c8_rr0 + t3_r0_c8_rr1;

  assign c_0_8 = t4_r0_c8_rr0;
  assign t0_r0_c9_rr0 = a_0_0 * b_0_9;
  assign t0_r0_c9_rr1 = a_0_1 * b_1_9;
  assign t0_r0_c9_rr2 = a_0_2 * b_2_9;
  assign t0_r0_c9_rr3 = a_0_3 * b_3_9;
  assign t0_r0_c9_rr4 = a_0_4 * b_4_9;
  assign t0_r0_c9_rr5 = a_0_5 * b_5_9;
  assign t0_r0_c9_rr6 = a_0_6 * b_6_9;
  assign t0_r0_c9_rr7 = a_0_7 * b_7_9;
  assign t0_r0_c9_rr8 = a_0_8 * b_8_9;
  assign t0_r0_c9_rr9 = a_0_9 * b_9_9;
  assign t1_r0_c9_rr0 = t0_r0_c9_rr0 + t0_r0_c9_rr1;
  assign t1_r0_c9_rr1 = t0_r0_c9_rr2 + t0_r0_c9_rr3;
  assign t1_r0_c9_rr2 = t0_r0_c9_rr4 + t0_r0_c9_rr5;
  assign t1_r0_c9_rr3 = t0_r0_c9_rr6 + t0_r0_c9_rr7;
  assign t1_r0_c9_rr4 = t0_r0_c9_rr8 + t0_r0_c9_rr9;

  assign t2_r0_c9_rr0 = t1_r0_c9_rr0 + t1_r0_c9_rr1;
  assign t2_r0_c9_rr1 = t1_r0_c9_rr2 + t1_r0_c9_rr3;
  assign t2_r0_c9_rr2 = t1_r0_c9_rr4;

  assign t3_r0_c9_rr0 = t2_r0_c9_rr0 + t2_r0_c9_rr1;
  assign t3_r0_c9_rr1 = t2_r0_c9_rr2;

  assign t4_r0_c9_rr0 = t3_r0_c9_rr0 + t3_r0_c9_rr1;

  assign c_0_9 = t4_r0_c9_rr0;
  assign t0_r1_c0_rr0 = a_1_0 * b_0_0;
  assign t0_r1_c0_rr1 = a_1_1 * b_1_0;
  assign t0_r1_c0_rr2 = a_1_2 * b_2_0;
  assign t0_r1_c0_rr3 = a_1_3 * b_3_0;
  assign t0_r1_c0_rr4 = a_1_4 * b_4_0;
  assign t0_r1_c0_rr5 = a_1_5 * b_5_0;
  assign t0_r1_c0_rr6 = a_1_6 * b_6_0;
  assign t0_r1_c0_rr7 = a_1_7 * b_7_0;
  assign t0_r1_c0_rr8 = a_1_8 * b_8_0;
  assign t0_r1_c0_rr9 = a_1_9 * b_9_0;
  assign t1_r1_c0_rr0 = t0_r1_c0_rr0 + t0_r1_c0_rr1;
  assign t1_r1_c0_rr1 = t0_r1_c0_rr2 + t0_r1_c0_rr3;
  assign t1_r1_c0_rr2 = t0_r1_c0_rr4 + t0_r1_c0_rr5;
  assign t1_r1_c0_rr3 = t0_r1_c0_rr6 + t0_r1_c0_rr7;
  assign t1_r1_c0_rr4 = t0_r1_c0_rr8 + t0_r1_c0_rr9;

  assign t2_r1_c0_rr0 = t1_r1_c0_rr0 + t1_r1_c0_rr1;
  assign t2_r1_c0_rr1 = t1_r1_c0_rr2 + t1_r1_c0_rr3;
  assign t2_r1_c0_rr2 = t1_r1_c0_rr4;

  assign t3_r1_c0_rr0 = t2_r1_c0_rr0 + t2_r1_c0_rr1;
  assign t3_r1_c0_rr1 = t2_r1_c0_rr2;

  assign t4_r1_c0_rr0 = t3_r1_c0_rr0 + t3_r1_c0_rr1;

  assign c_1_0 = t4_r1_c0_rr0;
  assign t0_r1_c1_rr0 = a_1_0 * b_0_1;
  assign t0_r1_c1_rr1 = a_1_1 * b_1_1;
  assign t0_r1_c1_rr2 = a_1_2 * b_2_1;
  assign t0_r1_c1_rr3 = a_1_3 * b_3_1;
  assign t0_r1_c1_rr4 = a_1_4 * b_4_1;
  assign t0_r1_c1_rr5 = a_1_5 * b_5_1;
  assign t0_r1_c1_rr6 = a_1_6 * b_6_1;
  assign t0_r1_c1_rr7 = a_1_7 * b_7_1;
  assign t0_r1_c1_rr8 = a_1_8 * b_8_1;
  assign t0_r1_c1_rr9 = a_1_9 * b_9_1;
  assign t1_r1_c1_rr0 = t0_r1_c1_rr0 + t0_r1_c1_rr1;
  assign t1_r1_c1_rr1 = t0_r1_c1_rr2 + t0_r1_c1_rr3;
  assign t1_r1_c1_rr2 = t0_r1_c1_rr4 + t0_r1_c1_rr5;
  assign t1_r1_c1_rr3 = t0_r1_c1_rr6 + t0_r1_c1_rr7;
  assign t1_r1_c1_rr4 = t0_r1_c1_rr8 + t0_r1_c1_rr9;

  assign t2_r1_c1_rr0 = t1_r1_c1_rr0 + t1_r1_c1_rr1;
  assign t2_r1_c1_rr1 = t1_r1_c1_rr2 + t1_r1_c1_rr3;
  assign t2_r1_c1_rr2 = t1_r1_c1_rr4;

  assign t3_r1_c1_rr0 = t2_r1_c1_rr0 + t2_r1_c1_rr1;
  assign t3_r1_c1_rr1 = t2_r1_c1_rr2;

  assign t4_r1_c1_rr0 = t3_r1_c1_rr0 + t3_r1_c1_rr1;

  assign c_1_1 = t4_r1_c1_rr0;
  assign t0_r1_c2_rr0 = a_1_0 * b_0_2;
  assign t0_r1_c2_rr1 = a_1_1 * b_1_2;
  assign t0_r1_c2_rr2 = a_1_2 * b_2_2;
  assign t0_r1_c2_rr3 = a_1_3 * b_3_2;
  assign t0_r1_c2_rr4 = a_1_4 * b_4_2;
  assign t0_r1_c2_rr5 = a_1_5 * b_5_2;
  assign t0_r1_c2_rr6 = a_1_6 * b_6_2;
  assign t0_r1_c2_rr7 = a_1_7 * b_7_2;
  assign t0_r1_c2_rr8 = a_1_8 * b_8_2;
  assign t0_r1_c2_rr9 = a_1_9 * b_9_2;
  assign t1_r1_c2_rr0 = t0_r1_c2_rr0 + t0_r1_c2_rr1;
  assign t1_r1_c2_rr1 = t0_r1_c2_rr2 + t0_r1_c2_rr3;
  assign t1_r1_c2_rr2 = t0_r1_c2_rr4 + t0_r1_c2_rr5;
  assign t1_r1_c2_rr3 = t0_r1_c2_rr6 + t0_r1_c2_rr7;
  assign t1_r1_c2_rr4 = t0_r1_c2_rr8 + t0_r1_c2_rr9;

  assign t2_r1_c2_rr0 = t1_r1_c2_rr0 + t1_r1_c2_rr1;
  assign t2_r1_c2_rr1 = t1_r1_c2_rr2 + t1_r1_c2_rr3;
  assign t2_r1_c2_rr2 = t1_r1_c2_rr4;

  assign t3_r1_c2_rr0 = t2_r1_c2_rr0 + t2_r1_c2_rr1;
  assign t3_r1_c2_rr1 = t2_r1_c2_rr2;

  assign t4_r1_c2_rr0 = t3_r1_c2_rr0 + t3_r1_c2_rr1;

  assign c_1_2 = t4_r1_c2_rr0;
  assign t0_r1_c3_rr0 = a_1_0 * b_0_3;
  assign t0_r1_c3_rr1 = a_1_1 * b_1_3;
  assign t0_r1_c3_rr2 = a_1_2 * b_2_3;
  assign t0_r1_c3_rr3 = a_1_3 * b_3_3;
  assign t0_r1_c3_rr4 = a_1_4 * b_4_3;
  assign t0_r1_c3_rr5 = a_1_5 * b_5_3;
  assign t0_r1_c3_rr6 = a_1_6 * b_6_3;
  assign t0_r1_c3_rr7 = a_1_7 * b_7_3;
  assign t0_r1_c3_rr8 = a_1_8 * b_8_3;
  assign t0_r1_c3_rr9 = a_1_9 * b_9_3;
  assign t1_r1_c3_rr0 = t0_r1_c3_rr0 + t0_r1_c3_rr1;
  assign t1_r1_c3_rr1 = t0_r1_c3_rr2 + t0_r1_c3_rr3;
  assign t1_r1_c3_rr2 = t0_r1_c3_rr4 + t0_r1_c3_rr5;
  assign t1_r1_c3_rr3 = t0_r1_c3_rr6 + t0_r1_c3_rr7;
  assign t1_r1_c3_rr4 = t0_r1_c3_rr8 + t0_r1_c3_rr9;

  assign t2_r1_c3_rr0 = t1_r1_c3_rr0 + t1_r1_c3_rr1;
  assign t2_r1_c3_rr1 = t1_r1_c3_rr2 + t1_r1_c3_rr3;
  assign t2_r1_c3_rr2 = t1_r1_c3_rr4;

  assign t3_r1_c3_rr0 = t2_r1_c3_rr0 + t2_r1_c3_rr1;
  assign t3_r1_c3_rr1 = t2_r1_c3_rr2;

  assign t4_r1_c3_rr0 = t3_r1_c3_rr0 + t3_r1_c3_rr1;

  assign c_1_3 = t4_r1_c3_rr0;
  assign t0_r1_c4_rr0 = a_1_0 * b_0_4;
  assign t0_r1_c4_rr1 = a_1_1 * b_1_4;
  assign t0_r1_c4_rr2 = a_1_2 * b_2_4;
  assign t0_r1_c4_rr3 = a_1_3 * b_3_4;
  assign t0_r1_c4_rr4 = a_1_4 * b_4_4;
  assign t0_r1_c4_rr5 = a_1_5 * b_5_4;
  assign t0_r1_c4_rr6 = a_1_6 * b_6_4;
  assign t0_r1_c4_rr7 = a_1_7 * b_7_4;
  assign t0_r1_c4_rr8 = a_1_8 * b_8_4;
  assign t0_r1_c4_rr9 = a_1_9 * b_9_4;
  assign t1_r1_c4_rr0 = t0_r1_c4_rr0 + t0_r1_c4_rr1;
  assign t1_r1_c4_rr1 = t0_r1_c4_rr2 + t0_r1_c4_rr3;
  assign t1_r1_c4_rr2 = t0_r1_c4_rr4 + t0_r1_c4_rr5;
  assign t1_r1_c4_rr3 = t0_r1_c4_rr6 + t0_r1_c4_rr7;
  assign t1_r1_c4_rr4 = t0_r1_c4_rr8 + t0_r1_c4_rr9;

  assign t2_r1_c4_rr0 = t1_r1_c4_rr0 + t1_r1_c4_rr1;
  assign t2_r1_c4_rr1 = t1_r1_c4_rr2 + t1_r1_c4_rr3;
  assign t2_r1_c4_rr2 = t1_r1_c4_rr4;

  assign t3_r1_c4_rr0 = t2_r1_c4_rr0 + t2_r1_c4_rr1;
  assign t3_r1_c4_rr1 = t2_r1_c4_rr2;

  assign t4_r1_c4_rr0 = t3_r1_c4_rr0 + t3_r1_c4_rr1;

  assign c_1_4 = t4_r1_c4_rr0;
  assign t0_r1_c5_rr0 = a_1_0 * b_0_5;
  assign t0_r1_c5_rr1 = a_1_1 * b_1_5;
  assign t0_r1_c5_rr2 = a_1_2 * b_2_5;
  assign t0_r1_c5_rr3 = a_1_3 * b_3_5;
  assign t0_r1_c5_rr4 = a_1_4 * b_4_5;
  assign t0_r1_c5_rr5 = a_1_5 * b_5_5;
  assign t0_r1_c5_rr6 = a_1_6 * b_6_5;
  assign t0_r1_c5_rr7 = a_1_7 * b_7_5;
  assign t0_r1_c5_rr8 = a_1_8 * b_8_5;
  assign t0_r1_c5_rr9 = a_1_9 * b_9_5;
  assign t1_r1_c5_rr0 = t0_r1_c5_rr0 + t0_r1_c5_rr1;
  assign t1_r1_c5_rr1 = t0_r1_c5_rr2 + t0_r1_c5_rr3;
  assign t1_r1_c5_rr2 = t0_r1_c5_rr4 + t0_r1_c5_rr5;
  assign t1_r1_c5_rr3 = t0_r1_c5_rr6 + t0_r1_c5_rr7;
  assign t1_r1_c5_rr4 = t0_r1_c5_rr8 + t0_r1_c5_rr9;

  assign t2_r1_c5_rr0 = t1_r1_c5_rr0 + t1_r1_c5_rr1;
  assign t2_r1_c5_rr1 = t1_r1_c5_rr2 + t1_r1_c5_rr3;
  assign t2_r1_c5_rr2 = t1_r1_c5_rr4;

  assign t3_r1_c5_rr0 = t2_r1_c5_rr0 + t2_r1_c5_rr1;
  assign t3_r1_c5_rr1 = t2_r1_c5_rr2;

  assign t4_r1_c5_rr0 = t3_r1_c5_rr0 + t3_r1_c5_rr1;

  assign c_1_5 = t4_r1_c5_rr0;
  assign t0_r1_c6_rr0 = a_1_0 * b_0_6;
  assign t0_r1_c6_rr1 = a_1_1 * b_1_6;
  assign t0_r1_c6_rr2 = a_1_2 * b_2_6;
  assign t0_r1_c6_rr3 = a_1_3 * b_3_6;
  assign t0_r1_c6_rr4 = a_1_4 * b_4_6;
  assign t0_r1_c6_rr5 = a_1_5 * b_5_6;
  assign t0_r1_c6_rr6 = a_1_6 * b_6_6;
  assign t0_r1_c6_rr7 = a_1_7 * b_7_6;
  assign t0_r1_c6_rr8 = a_1_8 * b_8_6;
  assign t0_r1_c6_rr9 = a_1_9 * b_9_6;
  assign t1_r1_c6_rr0 = t0_r1_c6_rr0 + t0_r1_c6_rr1;
  assign t1_r1_c6_rr1 = t0_r1_c6_rr2 + t0_r1_c6_rr3;
  assign t1_r1_c6_rr2 = t0_r1_c6_rr4 + t0_r1_c6_rr5;
  assign t1_r1_c6_rr3 = t0_r1_c6_rr6 + t0_r1_c6_rr7;
  assign t1_r1_c6_rr4 = t0_r1_c6_rr8 + t0_r1_c6_rr9;

  assign t2_r1_c6_rr0 = t1_r1_c6_rr0 + t1_r1_c6_rr1;
  assign t2_r1_c6_rr1 = t1_r1_c6_rr2 + t1_r1_c6_rr3;
  assign t2_r1_c6_rr2 = t1_r1_c6_rr4;

  assign t3_r1_c6_rr0 = t2_r1_c6_rr0 + t2_r1_c6_rr1;
  assign t3_r1_c6_rr1 = t2_r1_c6_rr2;

  assign t4_r1_c6_rr0 = t3_r1_c6_rr0 + t3_r1_c6_rr1;

  assign c_1_6 = t4_r1_c6_rr0;
  assign t0_r1_c7_rr0 = a_1_0 * b_0_7;
  assign t0_r1_c7_rr1 = a_1_1 * b_1_7;
  assign t0_r1_c7_rr2 = a_1_2 * b_2_7;
  assign t0_r1_c7_rr3 = a_1_3 * b_3_7;
  assign t0_r1_c7_rr4 = a_1_4 * b_4_7;
  assign t0_r1_c7_rr5 = a_1_5 * b_5_7;
  assign t0_r1_c7_rr6 = a_1_6 * b_6_7;
  assign t0_r1_c7_rr7 = a_1_7 * b_7_7;
  assign t0_r1_c7_rr8 = a_1_8 * b_8_7;
  assign t0_r1_c7_rr9 = a_1_9 * b_9_7;
  assign t1_r1_c7_rr0 = t0_r1_c7_rr0 + t0_r1_c7_rr1;
  assign t1_r1_c7_rr1 = t0_r1_c7_rr2 + t0_r1_c7_rr3;
  assign t1_r1_c7_rr2 = t0_r1_c7_rr4 + t0_r1_c7_rr5;
  assign t1_r1_c7_rr3 = t0_r1_c7_rr6 + t0_r1_c7_rr7;
  assign t1_r1_c7_rr4 = t0_r1_c7_rr8 + t0_r1_c7_rr9;

  assign t2_r1_c7_rr0 = t1_r1_c7_rr0 + t1_r1_c7_rr1;
  assign t2_r1_c7_rr1 = t1_r1_c7_rr2 + t1_r1_c7_rr3;
  assign t2_r1_c7_rr2 = t1_r1_c7_rr4;

  assign t3_r1_c7_rr0 = t2_r1_c7_rr0 + t2_r1_c7_rr1;
  assign t3_r1_c7_rr1 = t2_r1_c7_rr2;

  assign t4_r1_c7_rr0 = t3_r1_c7_rr0 + t3_r1_c7_rr1;

  assign c_1_7 = t4_r1_c7_rr0;
  assign t0_r1_c8_rr0 = a_1_0 * b_0_8;
  assign t0_r1_c8_rr1 = a_1_1 * b_1_8;
  assign t0_r1_c8_rr2 = a_1_2 * b_2_8;
  assign t0_r1_c8_rr3 = a_1_3 * b_3_8;
  assign t0_r1_c8_rr4 = a_1_4 * b_4_8;
  assign t0_r1_c8_rr5 = a_1_5 * b_5_8;
  assign t0_r1_c8_rr6 = a_1_6 * b_6_8;
  assign t0_r1_c8_rr7 = a_1_7 * b_7_8;
  assign t0_r1_c8_rr8 = a_1_8 * b_8_8;
  assign t0_r1_c8_rr9 = a_1_9 * b_9_8;
  assign t1_r1_c8_rr0 = t0_r1_c8_rr0 + t0_r1_c8_rr1;
  assign t1_r1_c8_rr1 = t0_r1_c8_rr2 + t0_r1_c8_rr3;
  assign t1_r1_c8_rr2 = t0_r1_c8_rr4 + t0_r1_c8_rr5;
  assign t1_r1_c8_rr3 = t0_r1_c8_rr6 + t0_r1_c8_rr7;
  assign t1_r1_c8_rr4 = t0_r1_c8_rr8 + t0_r1_c8_rr9;

  assign t2_r1_c8_rr0 = t1_r1_c8_rr0 + t1_r1_c8_rr1;
  assign t2_r1_c8_rr1 = t1_r1_c8_rr2 + t1_r1_c8_rr3;
  assign t2_r1_c8_rr2 = t1_r1_c8_rr4;

  assign t3_r1_c8_rr0 = t2_r1_c8_rr0 + t2_r1_c8_rr1;
  assign t3_r1_c8_rr1 = t2_r1_c8_rr2;

  assign t4_r1_c8_rr0 = t3_r1_c8_rr0 + t3_r1_c8_rr1;

  assign c_1_8 = t4_r1_c8_rr0;
  assign t0_r1_c9_rr0 = a_1_0 * b_0_9;
  assign t0_r1_c9_rr1 = a_1_1 * b_1_9;
  assign t0_r1_c9_rr2 = a_1_2 * b_2_9;
  assign t0_r1_c9_rr3 = a_1_3 * b_3_9;
  assign t0_r1_c9_rr4 = a_1_4 * b_4_9;
  assign t0_r1_c9_rr5 = a_1_5 * b_5_9;
  assign t0_r1_c9_rr6 = a_1_6 * b_6_9;
  assign t0_r1_c9_rr7 = a_1_7 * b_7_9;
  assign t0_r1_c9_rr8 = a_1_8 * b_8_9;
  assign t0_r1_c9_rr9 = a_1_9 * b_9_9;
  assign t1_r1_c9_rr0 = t0_r1_c9_rr0 + t0_r1_c9_rr1;
  assign t1_r1_c9_rr1 = t0_r1_c9_rr2 + t0_r1_c9_rr3;
  assign t1_r1_c9_rr2 = t0_r1_c9_rr4 + t0_r1_c9_rr5;
  assign t1_r1_c9_rr3 = t0_r1_c9_rr6 + t0_r1_c9_rr7;
  assign t1_r1_c9_rr4 = t0_r1_c9_rr8 + t0_r1_c9_rr9;

  assign t2_r1_c9_rr0 = t1_r1_c9_rr0 + t1_r1_c9_rr1;
  assign t2_r1_c9_rr1 = t1_r1_c9_rr2 + t1_r1_c9_rr3;
  assign t2_r1_c9_rr2 = t1_r1_c9_rr4;

  assign t3_r1_c9_rr0 = t2_r1_c9_rr0 + t2_r1_c9_rr1;
  assign t3_r1_c9_rr1 = t2_r1_c9_rr2;

  assign t4_r1_c9_rr0 = t3_r1_c9_rr0 + t3_r1_c9_rr1;

  assign c_1_9 = t4_r1_c9_rr0;
  assign t0_r2_c0_rr0 = a_2_0 * b_0_0;
  assign t0_r2_c0_rr1 = a_2_1 * b_1_0;
  assign t0_r2_c0_rr2 = a_2_2 * b_2_0;
  assign t0_r2_c0_rr3 = a_2_3 * b_3_0;
  assign t0_r2_c0_rr4 = a_2_4 * b_4_0;
  assign t0_r2_c0_rr5 = a_2_5 * b_5_0;
  assign t0_r2_c0_rr6 = a_2_6 * b_6_0;
  assign t0_r2_c0_rr7 = a_2_7 * b_7_0;
  assign t0_r2_c0_rr8 = a_2_8 * b_8_0;
  assign t0_r2_c0_rr9 = a_2_9 * b_9_0;
  assign t1_r2_c0_rr0 = t0_r2_c0_rr0 + t0_r2_c0_rr1;
  assign t1_r2_c0_rr1 = t0_r2_c0_rr2 + t0_r2_c0_rr3;
  assign t1_r2_c0_rr2 = t0_r2_c0_rr4 + t0_r2_c0_rr5;
  assign t1_r2_c0_rr3 = t0_r2_c0_rr6 + t0_r2_c0_rr7;
  assign t1_r2_c0_rr4 = t0_r2_c0_rr8 + t0_r2_c0_rr9;

  assign t2_r2_c0_rr0 = t1_r2_c0_rr0 + t1_r2_c0_rr1;
  assign t2_r2_c0_rr1 = t1_r2_c0_rr2 + t1_r2_c0_rr3;
  assign t2_r2_c0_rr2 = t1_r2_c0_rr4;

  assign t3_r2_c0_rr0 = t2_r2_c0_rr0 + t2_r2_c0_rr1;
  assign t3_r2_c0_rr1 = t2_r2_c0_rr2;

  assign t4_r2_c0_rr0 = t3_r2_c0_rr0 + t3_r2_c0_rr1;

  assign c_2_0 = t4_r2_c0_rr0;
  assign t0_r2_c1_rr0 = a_2_0 * b_0_1;
  assign t0_r2_c1_rr1 = a_2_1 * b_1_1;
  assign t0_r2_c1_rr2 = a_2_2 * b_2_1;
  assign t0_r2_c1_rr3 = a_2_3 * b_3_1;
  assign t0_r2_c1_rr4 = a_2_4 * b_4_1;
  assign t0_r2_c1_rr5 = a_2_5 * b_5_1;
  assign t0_r2_c1_rr6 = a_2_6 * b_6_1;
  assign t0_r2_c1_rr7 = a_2_7 * b_7_1;
  assign t0_r2_c1_rr8 = a_2_8 * b_8_1;
  assign t0_r2_c1_rr9 = a_2_9 * b_9_1;
  assign t1_r2_c1_rr0 = t0_r2_c1_rr0 + t0_r2_c1_rr1;
  assign t1_r2_c1_rr1 = t0_r2_c1_rr2 + t0_r2_c1_rr3;
  assign t1_r2_c1_rr2 = t0_r2_c1_rr4 + t0_r2_c1_rr5;
  assign t1_r2_c1_rr3 = t0_r2_c1_rr6 + t0_r2_c1_rr7;
  assign t1_r2_c1_rr4 = t0_r2_c1_rr8 + t0_r2_c1_rr9;

  assign t2_r2_c1_rr0 = t1_r2_c1_rr0 + t1_r2_c1_rr1;
  assign t2_r2_c1_rr1 = t1_r2_c1_rr2 + t1_r2_c1_rr3;
  assign t2_r2_c1_rr2 = t1_r2_c1_rr4;

  assign t3_r2_c1_rr0 = t2_r2_c1_rr0 + t2_r2_c1_rr1;
  assign t3_r2_c1_rr1 = t2_r2_c1_rr2;

  assign t4_r2_c1_rr0 = t3_r2_c1_rr0 + t3_r2_c1_rr1;

  assign c_2_1 = t4_r2_c1_rr0;
  assign t0_r2_c2_rr0 = a_2_0 * b_0_2;
  assign t0_r2_c2_rr1 = a_2_1 * b_1_2;
  assign t0_r2_c2_rr2 = a_2_2 * b_2_2;
  assign t0_r2_c2_rr3 = a_2_3 * b_3_2;
  assign t0_r2_c2_rr4 = a_2_4 * b_4_2;
  assign t0_r2_c2_rr5 = a_2_5 * b_5_2;
  assign t0_r2_c2_rr6 = a_2_6 * b_6_2;
  assign t0_r2_c2_rr7 = a_2_7 * b_7_2;
  assign t0_r2_c2_rr8 = a_2_8 * b_8_2;
  assign t0_r2_c2_rr9 = a_2_9 * b_9_2;
  assign t1_r2_c2_rr0 = t0_r2_c2_rr0 + t0_r2_c2_rr1;
  assign t1_r2_c2_rr1 = t0_r2_c2_rr2 + t0_r2_c2_rr3;
  assign t1_r2_c2_rr2 = t0_r2_c2_rr4 + t0_r2_c2_rr5;
  assign t1_r2_c2_rr3 = t0_r2_c2_rr6 + t0_r2_c2_rr7;
  assign t1_r2_c2_rr4 = t0_r2_c2_rr8 + t0_r2_c2_rr9;

  assign t2_r2_c2_rr0 = t1_r2_c2_rr0 + t1_r2_c2_rr1;
  assign t2_r2_c2_rr1 = t1_r2_c2_rr2 + t1_r2_c2_rr3;
  assign t2_r2_c2_rr2 = t1_r2_c2_rr4;

  assign t3_r2_c2_rr0 = t2_r2_c2_rr0 + t2_r2_c2_rr1;
  assign t3_r2_c2_rr1 = t2_r2_c2_rr2;

  assign t4_r2_c2_rr0 = t3_r2_c2_rr0 + t3_r2_c2_rr1;

  assign c_2_2 = t4_r2_c2_rr0;
  assign t0_r2_c3_rr0 = a_2_0 * b_0_3;
  assign t0_r2_c3_rr1 = a_2_1 * b_1_3;
  assign t0_r2_c3_rr2 = a_2_2 * b_2_3;
  assign t0_r2_c3_rr3 = a_2_3 * b_3_3;
  assign t0_r2_c3_rr4 = a_2_4 * b_4_3;
  assign t0_r2_c3_rr5 = a_2_5 * b_5_3;
  assign t0_r2_c3_rr6 = a_2_6 * b_6_3;
  assign t0_r2_c3_rr7 = a_2_7 * b_7_3;
  assign t0_r2_c3_rr8 = a_2_8 * b_8_3;
  assign t0_r2_c3_rr9 = a_2_9 * b_9_3;
  assign t1_r2_c3_rr0 = t0_r2_c3_rr0 + t0_r2_c3_rr1;
  assign t1_r2_c3_rr1 = t0_r2_c3_rr2 + t0_r2_c3_rr3;
  assign t1_r2_c3_rr2 = t0_r2_c3_rr4 + t0_r2_c3_rr5;
  assign t1_r2_c3_rr3 = t0_r2_c3_rr6 + t0_r2_c3_rr7;
  assign t1_r2_c3_rr4 = t0_r2_c3_rr8 + t0_r2_c3_rr9;

  assign t2_r2_c3_rr0 = t1_r2_c3_rr0 + t1_r2_c3_rr1;
  assign t2_r2_c3_rr1 = t1_r2_c3_rr2 + t1_r2_c3_rr3;
  assign t2_r2_c3_rr2 = t1_r2_c3_rr4;

  assign t3_r2_c3_rr0 = t2_r2_c3_rr0 + t2_r2_c3_rr1;
  assign t3_r2_c3_rr1 = t2_r2_c3_rr2;

  assign t4_r2_c3_rr0 = t3_r2_c3_rr0 + t3_r2_c3_rr1;

  assign c_2_3 = t4_r2_c3_rr0;
  assign t0_r2_c4_rr0 = a_2_0 * b_0_4;
  assign t0_r2_c4_rr1 = a_2_1 * b_1_4;
  assign t0_r2_c4_rr2 = a_2_2 * b_2_4;
  assign t0_r2_c4_rr3 = a_2_3 * b_3_4;
  assign t0_r2_c4_rr4 = a_2_4 * b_4_4;
  assign t0_r2_c4_rr5 = a_2_5 * b_5_4;
  assign t0_r2_c4_rr6 = a_2_6 * b_6_4;
  assign t0_r2_c4_rr7 = a_2_7 * b_7_4;
  assign t0_r2_c4_rr8 = a_2_8 * b_8_4;
  assign t0_r2_c4_rr9 = a_2_9 * b_9_4;
  assign t1_r2_c4_rr0 = t0_r2_c4_rr0 + t0_r2_c4_rr1;
  assign t1_r2_c4_rr1 = t0_r2_c4_rr2 + t0_r2_c4_rr3;
  assign t1_r2_c4_rr2 = t0_r2_c4_rr4 + t0_r2_c4_rr5;
  assign t1_r2_c4_rr3 = t0_r2_c4_rr6 + t0_r2_c4_rr7;
  assign t1_r2_c4_rr4 = t0_r2_c4_rr8 + t0_r2_c4_rr9;

  assign t2_r2_c4_rr0 = t1_r2_c4_rr0 + t1_r2_c4_rr1;
  assign t2_r2_c4_rr1 = t1_r2_c4_rr2 + t1_r2_c4_rr3;
  assign t2_r2_c4_rr2 = t1_r2_c4_rr4;

  assign t3_r2_c4_rr0 = t2_r2_c4_rr0 + t2_r2_c4_rr1;
  assign t3_r2_c4_rr1 = t2_r2_c4_rr2;

  assign t4_r2_c4_rr0 = t3_r2_c4_rr0 + t3_r2_c4_rr1;

  assign c_2_4 = t4_r2_c4_rr0;
  assign t0_r2_c5_rr0 = a_2_0 * b_0_5;
  assign t0_r2_c5_rr1 = a_2_1 * b_1_5;
  assign t0_r2_c5_rr2 = a_2_2 * b_2_5;
  assign t0_r2_c5_rr3 = a_2_3 * b_3_5;
  assign t0_r2_c5_rr4 = a_2_4 * b_4_5;
  assign t0_r2_c5_rr5 = a_2_5 * b_5_5;
  assign t0_r2_c5_rr6 = a_2_6 * b_6_5;
  assign t0_r2_c5_rr7 = a_2_7 * b_7_5;
  assign t0_r2_c5_rr8 = a_2_8 * b_8_5;
  assign t0_r2_c5_rr9 = a_2_9 * b_9_5;
  assign t1_r2_c5_rr0 = t0_r2_c5_rr0 + t0_r2_c5_rr1;
  assign t1_r2_c5_rr1 = t0_r2_c5_rr2 + t0_r2_c5_rr3;
  assign t1_r2_c5_rr2 = t0_r2_c5_rr4 + t0_r2_c5_rr5;
  assign t1_r2_c5_rr3 = t0_r2_c5_rr6 + t0_r2_c5_rr7;
  assign t1_r2_c5_rr4 = t0_r2_c5_rr8 + t0_r2_c5_rr9;

  assign t2_r2_c5_rr0 = t1_r2_c5_rr0 + t1_r2_c5_rr1;
  assign t2_r2_c5_rr1 = t1_r2_c5_rr2 + t1_r2_c5_rr3;
  assign t2_r2_c5_rr2 = t1_r2_c5_rr4;

  assign t3_r2_c5_rr0 = t2_r2_c5_rr0 + t2_r2_c5_rr1;
  assign t3_r2_c5_rr1 = t2_r2_c5_rr2;

  assign t4_r2_c5_rr0 = t3_r2_c5_rr0 + t3_r2_c5_rr1;

  assign c_2_5 = t4_r2_c5_rr0;
  assign t0_r2_c6_rr0 = a_2_0 * b_0_6;
  assign t0_r2_c6_rr1 = a_2_1 * b_1_6;
  assign t0_r2_c6_rr2 = a_2_2 * b_2_6;
  assign t0_r2_c6_rr3 = a_2_3 * b_3_6;
  assign t0_r2_c6_rr4 = a_2_4 * b_4_6;
  assign t0_r2_c6_rr5 = a_2_5 * b_5_6;
  assign t0_r2_c6_rr6 = a_2_6 * b_6_6;
  assign t0_r2_c6_rr7 = a_2_7 * b_7_6;
  assign t0_r2_c6_rr8 = a_2_8 * b_8_6;
  assign t0_r2_c6_rr9 = a_2_9 * b_9_6;
  assign t1_r2_c6_rr0 = t0_r2_c6_rr0 + t0_r2_c6_rr1;
  assign t1_r2_c6_rr1 = t0_r2_c6_rr2 + t0_r2_c6_rr3;
  assign t1_r2_c6_rr2 = t0_r2_c6_rr4 + t0_r2_c6_rr5;
  assign t1_r2_c6_rr3 = t0_r2_c6_rr6 + t0_r2_c6_rr7;
  assign t1_r2_c6_rr4 = t0_r2_c6_rr8 + t0_r2_c6_rr9;

  assign t2_r2_c6_rr0 = t1_r2_c6_rr0 + t1_r2_c6_rr1;
  assign t2_r2_c6_rr1 = t1_r2_c6_rr2 + t1_r2_c6_rr3;
  assign t2_r2_c6_rr2 = t1_r2_c6_rr4;

  assign t3_r2_c6_rr0 = t2_r2_c6_rr0 + t2_r2_c6_rr1;
  assign t3_r2_c6_rr1 = t2_r2_c6_rr2;

  assign t4_r2_c6_rr0 = t3_r2_c6_rr0 + t3_r2_c6_rr1;

  assign c_2_6 = t4_r2_c6_rr0;
  assign t0_r2_c7_rr0 = a_2_0 * b_0_7;
  assign t0_r2_c7_rr1 = a_2_1 * b_1_7;
  assign t0_r2_c7_rr2 = a_2_2 * b_2_7;
  assign t0_r2_c7_rr3 = a_2_3 * b_3_7;
  assign t0_r2_c7_rr4 = a_2_4 * b_4_7;
  assign t0_r2_c7_rr5 = a_2_5 * b_5_7;
  assign t0_r2_c7_rr6 = a_2_6 * b_6_7;
  assign t0_r2_c7_rr7 = a_2_7 * b_7_7;
  assign t0_r2_c7_rr8 = a_2_8 * b_8_7;
  assign t0_r2_c7_rr9 = a_2_9 * b_9_7;
  assign t1_r2_c7_rr0 = t0_r2_c7_rr0 + t0_r2_c7_rr1;
  assign t1_r2_c7_rr1 = t0_r2_c7_rr2 + t0_r2_c7_rr3;
  assign t1_r2_c7_rr2 = t0_r2_c7_rr4 + t0_r2_c7_rr5;
  assign t1_r2_c7_rr3 = t0_r2_c7_rr6 + t0_r2_c7_rr7;
  assign t1_r2_c7_rr4 = t0_r2_c7_rr8 + t0_r2_c7_rr9;

  assign t2_r2_c7_rr0 = t1_r2_c7_rr0 + t1_r2_c7_rr1;
  assign t2_r2_c7_rr1 = t1_r2_c7_rr2 + t1_r2_c7_rr3;
  assign t2_r2_c7_rr2 = t1_r2_c7_rr4;

  assign t3_r2_c7_rr0 = t2_r2_c7_rr0 + t2_r2_c7_rr1;
  assign t3_r2_c7_rr1 = t2_r2_c7_rr2;

  assign t4_r2_c7_rr0 = t3_r2_c7_rr0 + t3_r2_c7_rr1;

  assign c_2_7 = t4_r2_c7_rr0;
  assign t0_r2_c8_rr0 = a_2_0 * b_0_8;
  assign t0_r2_c8_rr1 = a_2_1 * b_1_8;
  assign t0_r2_c8_rr2 = a_2_2 * b_2_8;
  assign t0_r2_c8_rr3 = a_2_3 * b_3_8;
  assign t0_r2_c8_rr4 = a_2_4 * b_4_8;
  assign t0_r2_c8_rr5 = a_2_5 * b_5_8;
  assign t0_r2_c8_rr6 = a_2_6 * b_6_8;
  assign t0_r2_c8_rr7 = a_2_7 * b_7_8;
  assign t0_r2_c8_rr8 = a_2_8 * b_8_8;
  assign t0_r2_c8_rr9 = a_2_9 * b_9_8;
  assign t1_r2_c8_rr0 = t0_r2_c8_rr0 + t0_r2_c8_rr1;
  assign t1_r2_c8_rr1 = t0_r2_c8_rr2 + t0_r2_c8_rr3;
  assign t1_r2_c8_rr2 = t0_r2_c8_rr4 + t0_r2_c8_rr5;
  assign t1_r2_c8_rr3 = t0_r2_c8_rr6 + t0_r2_c8_rr7;
  assign t1_r2_c8_rr4 = t0_r2_c8_rr8 + t0_r2_c8_rr9;

  assign t2_r2_c8_rr0 = t1_r2_c8_rr0 + t1_r2_c8_rr1;
  assign t2_r2_c8_rr1 = t1_r2_c8_rr2 + t1_r2_c8_rr3;
  assign t2_r2_c8_rr2 = t1_r2_c8_rr4;

  assign t3_r2_c8_rr0 = t2_r2_c8_rr0 + t2_r2_c8_rr1;
  assign t3_r2_c8_rr1 = t2_r2_c8_rr2;

  assign t4_r2_c8_rr0 = t3_r2_c8_rr0 + t3_r2_c8_rr1;

  assign c_2_8 = t4_r2_c8_rr0;
  assign t0_r2_c9_rr0 = a_2_0 * b_0_9;
  assign t0_r2_c9_rr1 = a_2_1 * b_1_9;
  assign t0_r2_c9_rr2 = a_2_2 * b_2_9;
  assign t0_r2_c9_rr3 = a_2_3 * b_3_9;
  assign t0_r2_c9_rr4 = a_2_4 * b_4_9;
  assign t0_r2_c9_rr5 = a_2_5 * b_5_9;
  assign t0_r2_c9_rr6 = a_2_6 * b_6_9;
  assign t0_r2_c9_rr7 = a_2_7 * b_7_9;
  assign t0_r2_c9_rr8 = a_2_8 * b_8_9;
  assign t0_r2_c9_rr9 = a_2_9 * b_9_9;
  assign t1_r2_c9_rr0 = t0_r2_c9_rr0 + t0_r2_c9_rr1;
  assign t1_r2_c9_rr1 = t0_r2_c9_rr2 + t0_r2_c9_rr3;
  assign t1_r2_c9_rr2 = t0_r2_c9_rr4 + t0_r2_c9_rr5;
  assign t1_r2_c9_rr3 = t0_r2_c9_rr6 + t0_r2_c9_rr7;
  assign t1_r2_c9_rr4 = t0_r2_c9_rr8 + t0_r2_c9_rr9;

  assign t2_r2_c9_rr0 = t1_r2_c9_rr0 + t1_r2_c9_rr1;
  assign t2_r2_c9_rr1 = t1_r2_c9_rr2 + t1_r2_c9_rr3;
  assign t2_r2_c9_rr2 = t1_r2_c9_rr4;

  assign t3_r2_c9_rr0 = t2_r2_c9_rr0 + t2_r2_c9_rr1;
  assign t3_r2_c9_rr1 = t2_r2_c9_rr2;

  assign t4_r2_c9_rr0 = t3_r2_c9_rr0 + t3_r2_c9_rr1;

  assign c_2_9 = t4_r2_c9_rr0;
  assign t0_r3_c0_rr0 = a_3_0 * b_0_0;
  assign t0_r3_c0_rr1 = a_3_1 * b_1_0;
  assign t0_r3_c0_rr2 = a_3_2 * b_2_0;
  assign t0_r3_c0_rr3 = a_3_3 * b_3_0;
  assign t0_r3_c0_rr4 = a_3_4 * b_4_0;
  assign t0_r3_c0_rr5 = a_3_5 * b_5_0;
  assign t0_r3_c0_rr6 = a_3_6 * b_6_0;
  assign t0_r3_c0_rr7 = a_3_7 * b_7_0;
  assign t0_r3_c0_rr8 = a_3_8 * b_8_0;
  assign t0_r3_c0_rr9 = a_3_9 * b_9_0;
  assign t1_r3_c0_rr0 = t0_r3_c0_rr0 + t0_r3_c0_rr1;
  assign t1_r3_c0_rr1 = t0_r3_c0_rr2 + t0_r3_c0_rr3;
  assign t1_r3_c0_rr2 = t0_r3_c0_rr4 + t0_r3_c0_rr5;
  assign t1_r3_c0_rr3 = t0_r3_c0_rr6 + t0_r3_c0_rr7;
  assign t1_r3_c0_rr4 = t0_r3_c0_rr8 + t0_r3_c0_rr9;

  assign t2_r3_c0_rr0 = t1_r3_c0_rr0 + t1_r3_c0_rr1;
  assign t2_r3_c0_rr1 = t1_r3_c0_rr2 + t1_r3_c0_rr3;
  assign t2_r3_c0_rr2 = t1_r3_c0_rr4;

  assign t3_r3_c0_rr0 = t2_r3_c0_rr0 + t2_r3_c0_rr1;
  assign t3_r3_c0_rr1 = t2_r3_c0_rr2;

  assign t4_r3_c0_rr0 = t3_r3_c0_rr0 + t3_r3_c0_rr1;

  assign c_3_0 = t4_r3_c0_rr0;
  assign t0_r3_c1_rr0 = a_3_0 * b_0_1;
  assign t0_r3_c1_rr1 = a_3_1 * b_1_1;
  assign t0_r3_c1_rr2 = a_3_2 * b_2_1;
  assign t0_r3_c1_rr3 = a_3_3 * b_3_1;
  assign t0_r3_c1_rr4 = a_3_4 * b_4_1;
  assign t0_r3_c1_rr5 = a_3_5 * b_5_1;
  assign t0_r3_c1_rr6 = a_3_6 * b_6_1;
  assign t0_r3_c1_rr7 = a_3_7 * b_7_1;
  assign t0_r3_c1_rr8 = a_3_8 * b_8_1;
  assign t0_r3_c1_rr9 = a_3_9 * b_9_1;
  assign t1_r3_c1_rr0 = t0_r3_c1_rr0 + t0_r3_c1_rr1;
  assign t1_r3_c1_rr1 = t0_r3_c1_rr2 + t0_r3_c1_rr3;
  assign t1_r3_c1_rr2 = t0_r3_c1_rr4 + t0_r3_c1_rr5;
  assign t1_r3_c1_rr3 = t0_r3_c1_rr6 + t0_r3_c1_rr7;
  assign t1_r3_c1_rr4 = t0_r3_c1_rr8 + t0_r3_c1_rr9;

  assign t2_r3_c1_rr0 = t1_r3_c1_rr0 + t1_r3_c1_rr1;
  assign t2_r3_c1_rr1 = t1_r3_c1_rr2 + t1_r3_c1_rr3;
  assign t2_r3_c1_rr2 = t1_r3_c1_rr4;

  assign t3_r3_c1_rr0 = t2_r3_c1_rr0 + t2_r3_c1_rr1;
  assign t3_r3_c1_rr1 = t2_r3_c1_rr2;

  assign t4_r3_c1_rr0 = t3_r3_c1_rr0 + t3_r3_c1_rr1;

  assign c_3_1 = t4_r3_c1_rr0;
  assign t0_r3_c2_rr0 = a_3_0 * b_0_2;
  assign t0_r3_c2_rr1 = a_3_1 * b_1_2;
  assign t0_r3_c2_rr2 = a_3_2 * b_2_2;
  assign t0_r3_c2_rr3 = a_3_3 * b_3_2;
  assign t0_r3_c2_rr4 = a_3_4 * b_4_2;
  assign t0_r3_c2_rr5 = a_3_5 * b_5_2;
  assign t0_r3_c2_rr6 = a_3_6 * b_6_2;
  assign t0_r3_c2_rr7 = a_3_7 * b_7_2;
  assign t0_r3_c2_rr8 = a_3_8 * b_8_2;
  assign t0_r3_c2_rr9 = a_3_9 * b_9_2;
  assign t1_r3_c2_rr0 = t0_r3_c2_rr0 + t0_r3_c2_rr1;
  assign t1_r3_c2_rr1 = t0_r3_c2_rr2 + t0_r3_c2_rr3;
  assign t1_r3_c2_rr2 = t0_r3_c2_rr4 + t0_r3_c2_rr5;
  assign t1_r3_c2_rr3 = t0_r3_c2_rr6 + t0_r3_c2_rr7;
  assign t1_r3_c2_rr4 = t0_r3_c2_rr8 + t0_r3_c2_rr9;

  assign t2_r3_c2_rr0 = t1_r3_c2_rr0 + t1_r3_c2_rr1;
  assign t2_r3_c2_rr1 = t1_r3_c2_rr2 + t1_r3_c2_rr3;
  assign t2_r3_c2_rr2 = t1_r3_c2_rr4;

  assign t3_r3_c2_rr0 = t2_r3_c2_rr0 + t2_r3_c2_rr1;
  assign t3_r3_c2_rr1 = t2_r3_c2_rr2;

  assign t4_r3_c2_rr0 = t3_r3_c2_rr0 + t3_r3_c2_rr1;

  assign c_3_2 = t4_r3_c2_rr0;
  assign t0_r3_c3_rr0 = a_3_0 * b_0_3;
  assign t0_r3_c3_rr1 = a_3_1 * b_1_3;
  assign t0_r3_c3_rr2 = a_3_2 * b_2_3;
  assign t0_r3_c3_rr3 = a_3_3 * b_3_3;
  assign t0_r3_c3_rr4 = a_3_4 * b_4_3;
  assign t0_r3_c3_rr5 = a_3_5 * b_5_3;
  assign t0_r3_c3_rr6 = a_3_6 * b_6_3;
  assign t0_r3_c3_rr7 = a_3_7 * b_7_3;
  assign t0_r3_c3_rr8 = a_3_8 * b_8_3;
  assign t0_r3_c3_rr9 = a_3_9 * b_9_3;
  assign t1_r3_c3_rr0 = t0_r3_c3_rr0 + t0_r3_c3_rr1;
  assign t1_r3_c3_rr1 = t0_r3_c3_rr2 + t0_r3_c3_rr3;
  assign t1_r3_c3_rr2 = t0_r3_c3_rr4 + t0_r3_c3_rr5;
  assign t1_r3_c3_rr3 = t0_r3_c3_rr6 + t0_r3_c3_rr7;
  assign t1_r3_c3_rr4 = t0_r3_c3_rr8 + t0_r3_c3_rr9;

  assign t2_r3_c3_rr0 = t1_r3_c3_rr0 + t1_r3_c3_rr1;
  assign t2_r3_c3_rr1 = t1_r3_c3_rr2 + t1_r3_c3_rr3;
  assign t2_r3_c3_rr2 = t1_r3_c3_rr4;

  assign t3_r3_c3_rr0 = t2_r3_c3_rr0 + t2_r3_c3_rr1;
  assign t3_r3_c3_rr1 = t2_r3_c3_rr2;

  assign t4_r3_c3_rr0 = t3_r3_c3_rr0 + t3_r3_c3_rr1;

  assign c_3_3 = t4_r3_c3_rr0;
  assign t0_r3_c4_rr0 = a_3_0 * b_0_4;
  assign t0_r3_c4_rr1 = a_3_1 * b_1_4;
  assign t0_r3_c4_rr2 = a_3_2 * b_2_4;
  assign t0_r3_c4_rr3 = a_3_3 * b_3_4;
  assign t0_r3_c4_rr4 = a_3_4 * b_4_4;
  assign t0_r3_c4_rr5 = a_3_5 * b_5_4;
  assign t0_r3_c4_rr6 = a_3_6 * b_6_4;
  assign t0_r3_c4_rr7 = a_3_7 * b_7_4;
  assign t0_r3_c4_rr8 = a_3_8 * b_8_4;
  assign t0_r3_c4_rr9 = a_3_9 * b_9_4;
  assign t1_r3_c4_rr0 = t0_r3_c4_rr0 + t0_r3_c4_rr1;
  assign t1_r3_c4_rr1 = t0_r3_c4_rr2 + t0_r3_c4_rr3;
  assign t1_r3_c4_rr2 = t0_r3_c4_rr4 + t0_r3_c4_rr5;
  assign t1_r3_c4_rr3 = t0_r3_c4_rr6 + t0_r3_c4_rr7;
  assign t1_r3_c4_rr4 = t0_r3_c4_rr8 + t0_r3_c4_rr9;

  assign t2_r3_c4_rr0 = t1_r3_c4_rr0 + t1_r3_c4_rr1;
  assign t2_r3_c4_rr1 = t1_r3_c4_rr2 + t1_r3_c4_rr3;
  assign t2_r3_c4_rr2 = t1_r3_c4_rr4;

  assign t3_r3_c4_rr0 = t2_r3_c4_rr0 + t2_r3_c4_rr1;
  assign t3_r3_c4_rr1 = t2_r3_c4_rr2;

  assign t4_r3_c4_rr0 = t3_r3_c4_rr0 + t3_r3_c4_rr1;

  assign c_3_4 = t4_r3_c4_rr0;
  assign t0_r3_c5_rr0 = a_3_0 * b_0_5;
  assign t0_r3_c5_rr1 = a_3_1 * b_1_5;
  assign t0_r3_c5_rr2 = a_3_2 * b_2_5;
  assign t0_r3_c5_rr3 = a_3_3 * b_3_5;
  assign t0_r3_c5_rr4 = a_3_4 * b_4_5;
  assign t0_r3_c5_rr5 = a_3_5 * b_5_5;
  assign t0_r3_c5_rr6 = a_3_6 * b_6_5;
  assign t0_r3_c5_rr7 = a_3_7 * b_7_5;
  assign t0_r3_c5_rr8 = a_3_8 * b_8_5;
  assign t0_r3_c5_rr9 = a_3_9 * b_9_5;
  assign t1_r3_c5_rr0 = t0_r3_c5_rr0 + t0_r3_c5_rr1;
  assign t1_r3_c5_rr1 = t0_r3_c5_rr2 + t0_r3_c5_rr3;
  assign t1_r3_c5_rr2 = t0_r3_c5_rr4 + t0_r3_c5_rr5;
  assign t1_r3_c5_rr3 = t0_r3_c5_rr6 + t0_r3_c5_rr7;
  assign t1_r3_c5_rr4 = t0_r3_c5_rr8 + t0_r3_c5_rr9;

  assign t2_r3_c5_rr0 = t1_r3_c5_rr0 + t1_r3_c5_rr1;
  assign t2_r3_c5_rr1 = t1_r3_c5_rr2 + t1_r3_c5_rr3;
  assign t2_r3_c5_rr2 = t1_r3_c5_rr4;

  assign t3_r3_c5_rr0 = t2_r3_c5_rr0 + t2_r3_c5_rr1;
  assign t3_r3_c5_rr1 = t2_r3_c5_rr2;

  assign t4_r3_c5_rr0 = t3_r3_c5_rr0 + t3_r3_c5_rr1;

  assign c_3_5 = t4_r3_c5_rr0;
  assign t0_r3_c6_rr0 = a_3_0 * b_0_6;
  assign t0_r3_c6_rr1 = a_3_1 * b_1_6;
  assign t0_r3_c6_rr2 = a_3_2 * b_2_6;
  assign t0_r3_c6_rr3 = a_3_3 * b_3_6;
  assign t0_r3_c6_rr4 = a_3_4 * b_4_6;
  assign t0_r3_c6_rr5 = a_3_5 * b_5_6;
  assign t0_r3_c6_rr6 = a_3_6 * b_6_6;
  assign t0_r3_c6_rr7 = a_3_7 * b_7_6;
  assign t0_r3_c6_rr8 = a_3_8 * b_8_6;
  assign t0_r3_c6_rr9 = a_3_9 * b_9_6;
  assign t1_r3_c6_rr0 = t0_r3_c6_rr0 + t0_r3_c6_rr1;
  assign t1_r3_c6_rr1 = t0_r3_c6_rr2 + t0_r3_c6_rr3;
  assign t1_r3_c6_rr2 = t0_r3_c6_rr4 + t0_r3_c6_rr5;
  assign t1_r3_c6_rr3 = t0_r3_c6_rr6 + t0_r3_c6_rr7;
  assign t1_r3_c6_rr4 = t0_r3_c6_rr8 + t0_r3_c6_rr9;

  assign t2_r3_c6_rr0 = t1_r3_c6_rr0 + t1_r3_c6_rr1;
  assign t2_r3_c6_rr1 = t1_r3_c6_rr2 + t1_r3_c6_rr3;
  assign t2_r3_c6_rr2 = t1_r3_c6_rr4;

  assign t3_r3_c6_rr0 = t2_r3_c6_rr0 + t2_r3_c6_rr1;
  assign t3_r3_c6_rr1 = t2_r3_c6_rr2;

  assign t4_r3_c6_rr0 = t3_r3_c6_rr0 + t3_r3_c6_rr1;

  assign c_3_6 = t4_r3_c6_rr0;
  assign t0_r3_c7_rr0 = a_3_0 * b_0_7;
  assign t0_r3_c7_rr1 = a_3_1 * b_1_7;
  assign t0_r3_c7_rr2 = a_3_2 * b_2_7;
  assign t0_r3_c7_rr3 = a_3_3 * b_3_7;
  assign t0_r3_c7_rr4 = a_3_4 * b_4_7;
  assign t0_r3_c7_rr5 = a_3_5 * b_5_7;
  assign t0_r3_c7_rr6 = a_3_6 * b_6_7;
  assign t0_r3_c7_rr7 = a_3_7 * b_7_7;
  assign t0_r3_c7_rr8 = a_3_8 * b_8_7;
  assign t0_r3_c7_rr9 = a_3_9 * b_9_7;
  assign t1_r3_c7_rr0 = t0_r3_c7_rr0 + t0_r3_c7_rr1;
  assign t1_r3_c7_rr1 = t0_r3_c7_rr2 + t0_r3_c7_rr3;
  assign t1_r3_c7_rr2 = t0_r3_c7_rr4 + t0_r3_c7_rr5;
  assign t1_r3_c7_rr3 = t0_r3_c7_rr6 + t0_r3_c7_rr7;
  assign t1_r3_c7_rr4 = t0_r3_c7_rr8 + t0_r3_c7_rr9;

  assign t2_r3_c7_rr0 = t1_r3_c7_rr0 + t1_r3_c7_rr1;
  assign t2_r3_c7_rr1 = t1_r3_c7_rr2 + t1_r3_c7_rr3;
  assign t2_r3_c7_rr2 = t1_r3_c7_rr4;

  assign t3_r3_c7_rr0 = t2_r3_c7_rr0 + t2_r3_c7_rr1;
  assign t3_r3_c7_rr1 = t2_r3_c7_rr2;

  assign t4_r3_c7_rr0 = t3_r3_c7_rr0 + t3_r3_c7_rr1;

  assign c_3_7 = t4_r3_c7_rr0;
  assign t0_r3_c8_rr0 = a_3_0 * b_0_8;
  assign t0_r3_c8_rr1 = a_3_1 * b_1_8;
  assign t0_r3_c8_rr2 = a_3_2 * b_2_8;
  assign t0_r3_c8_rr3 = a_3_3 * b_3_8;
  assign t0_r3_c8_rr4 = a_3_4 * b_4_8;
  assign t0_r3_c8_rr5 = a_3_5 * b_5_8;
  assign t0_r3_c8_rr6 = a_3_6 * b_6_8;
  assign t0_r3_c8_rr7 = a_3_7 * b_7_8;
  assign t0_r3_c8_rr8 = a_3_8 * b_8_8;
  assign t0_r3_c8_rr9 = a_3_9 * b_9_8;
  assign t1_r3_c8_rr0 = t0_r3_c8_rr0 + t0_r3_c8_rr1;
  assign t1_r3_c8_rr1 = t0_r3_c8_rr2 + t0_r3_c8_rr3;
  assign t1_r3_c8_rr2 = t0_r3_c8_rr4 + t0_r3_c8_rr5;
  assign t1_r3_c8_rr3 = t0_r3_c8_rr6 + t0_r3_c8_rr7;
  assign t1_r3_c8_rr4 = t0_r3_c8_rr8 + t0_r3_c8_rr9;

  assign t2_r3_c8_rr0 = t1_r3_c8_rr0 + t1_r3_c8_rr1;
  assign t2_r3_c8_rr1 = t1_r3_c8_rr2 + t1_r3_c8_rr3;
  assign t2_r3_c8_rr2 = t1_r3_c8_rr4;

  assign t3_r3_c8_rr0 = t2_r3_c8_rr0 + t2_r3_c8_rr1;
  assign t3_r3_c8_rr1 = t2_r3_c8_rr2;

  assign t4_r3_c8_rr0 = t3_r3_c8_rr0 + t3_r3_c8_rr1;

  assign c_3_8 = t4_r3_c8_rr0;
  assign t0_r3_c9_rr0 = a_3_0 * b_0_9;
  assign t0_r3_c9_rr1 = a_3_1 * b_1_9;
  assign t0_r3_c9_rr2 = a_3_2 * b_2_9;
  assign t0_r3_c9_rr3 = a_3_3 * b_3_9;
  assign t0_r3_c9_rr4 = a_3_4 * b_4_9;
  assign t0_r3_c9_rr5 = a_3_5 * b_5_9;
  assign t0_r3_c9_rr6 = a_3_6 * b_6_9;
  assign t0_r3_c9_rr7 = a_3_7 * b_7_9;
  assign t0_r3_c9_rr8 = a_3_8 * b_8_9;
  assign t0_r3_c9_rr9 = a_3_9 * b_9_9;
  assign t1_r3_c9_rr0 = t0_r3_c9_rr0 + t0_r3_c9_rr1;
  assign t1_r3_c9_rr1 = t0_r3_c9_rr2 + t0_r3_c9_rr3;
  assign t1_r3_c9_rr2 = t0_r3_c9_rr4 + t0_r3_c9_rr5;
  assign t1_r3_c9_rr3 = t0_r3_c9_rr6 + t0_r3_c9_rr7;
  assign t1_r3_c9_rr4 = t0_r3_c9_rr8 + t0_r3_c9_rr9;

  assign t2_r3_c9_rr0 = t1_r3_c9_rr0 + t1_r3_c9_rr1;
  assign t2_r3_c9_rr1 = t1_r3_c9_rr2 + t1_r3_c9_rr3;
  assign t2_r3_c9_rr2 = t1_r3_c9_rr4;

  assign t3_r3_c9_rr0 = t2_r3_c9_rr0 + t2_r3_c9_rr1;
  assign t3_r3_c9_rr1 = t2_r3_c9_rr2;

  assign t4_r3_c9_rr0 = t3_r3_c9_rr0 + t3_r3_c9_rr1;

  assign c_3_9 = t4_r3_c9_rr0;
  assign t0_r4_c0_rr0 = a_4_0 * b_0_0;
  assign t0_r4_c0_rr1 = a_4_1 * b_1_0;
  assign t0_r4_c0_rr2 = a_4_2 * b_2_0;
  assign t0_r4_c0_rr3 = a_4_3 * b_3_0;
  assign t0_r4_c0_rr4 = a_4_4 * b_4_0;
  assign t0_r4_c0_rr5 = a_4_5 * b_5_0;
  assign t0_r4_c0_rr6 = a_4_6 * b_6_0;
  assign t0_r4_c0_rr7 = a_4_7 * b_7_0;
  assign t0_r4_c0_rr8 = a_4_8 * b_8_0;
  assign t0_r4_c0_rr9 = a_4_9 * b_9_0;
  assign t1_r4_c0_rr0 = t0_r4_c0_rr0 + t0_r4_c0_rr1;
  assign t1_r4_c0_rr1 = t0_r4_c0_rr2 + t0_r4_c0_rr3;
  assign t1_r4_c0_rr2 = t0_r4_c0_rr4 + t0_r4_c0_rr5;
  assign t1_r4_c0_rr3 = t0_r4_c0_rr6 + t0_r4_c0_rr7;
  assign t1_r4_c0_rr4 = t0_r4_c0_rr8 + t0_r4_c0_rr9;

  assign t2_r4_c0_rr0 = t1_r4_c0_rr0 + t1_r4_c0_rr1;
  assign t2_r4_c0_rr1 = t1_r4_c0_rr2 + t1_r4_c0_rr3;
  assign t2_r4_c0_rr2 = t1_r4_c0_rr4;

  assign t3_r4_c0_rr0 = t2_r4_c0_rr0 + t2_r4_c0_rr1;
  assign t3_r4_c0_rr1 = t2_r4_c0_rr2;

  assign t4_r4_c0_rr0 = t3_r4_c0_rr0 + t3_r4_c0_rr1;

  assign c_4_0 = t4_r4_c0_rr0;
  assign t0_r4_c1_rr0 = a_4_0 * b_0_1;
  assign t0_r4_c1_rr1 = a_4_1 * b_1_1;
  assign t0_r4_c1_rr2 = a_4_2 * b_2_1;
  assign t0_r4_c1_rr3 = a_4_3 * b_3_1;
  assign t0_r4_c1_rr4 = a_4_4 * b_4_1;
  assign t0_r4_c1_rr5 = a_4_5 * b_5_1;
  assign t0_r4_c1_rr6 = a_4_6 * b_6_1;
  assign t0_r4_c1_rr7 = a_4_7 * b_7_1;
  assign t0_r4_c1_rr8 = a_4_8 * b_8_1;
  assign t0_r4_c1_rr9 = a_4_9 * b_9_1;
  assign t1_r4_c1_rr0 = t0_r4_c1_rr0 + t0_r4_c1_rr1;
  assign t1_r4_c1_rr1 = t0_r4_c1_rr2 + t0_r4_c1_rr3;
  assign t1_r4_c1_rr2 = t0_r4_c1_rr4 + t0_r4_c1_rr5;
  assign t1_r4_c1_rr3 = t0_r4_c1_rr6 + t0_r4_c1_rr7;
  assign t1_r4_c1_rr4 = t0_r4_c1_rr8 + t0_r4_c1_rr9;

  assign t2_r4_c1_rr0 = t1_r4_c1_rr0 + t1_r4_c1_rr1;
  assign t2_r4_c1_rr1 = t1_r4_c1_rr2 + t1_r4_c1_rr3;
  assign t2_r4_c1_rr2 = t1_r4_c1_rr4;

  assign t3_r4_c1_rr0 = t2_r4_c1_rr0 + t2_r4_c1_rr1;
  assign t3_r4_c1_rr1 = t2_r4_c1_rr2;

  assign t4_r4_c1_rr0 = t3_r4_c1_rr0 + t3_r4_c1_rr1;

  assign c_4_1 = t4_r4_c1_rr0;
  assign t0_r4_c2_rr0 = a_4_0 * b_0_2;
  assign t0_r4_c2_rr1 = a_4_1 * b_1_2;
  assign t0_r4_c2_rr2 = a_4_2 * b_2_2;
  assign t0_r4_c2_rr3 = a_4_3 * b_3_2;
  assign t0_r4_c2_rr4 = a_4_4 * b_4_2;
  assign t0_r4_c2_rr5 = a_4_5 * b_5_2;
  assign t0_r4_c2_rr6 = a_4_6 * b_6_2;
  assign t0_r4_c2_rr7 = a_4_7 * b_7_2;
  assign t0_r4_c2_rr8 = a_4_8 * b_8_2;
  assign t0_r4_c2_rr9 = a_4_9 * b_9_2;
  assign t1_r4_c2_rr0 = t0_r4_c2_rr0 + t0_r4_c2_rr1;
  assign t1_r4_c2_rr1 = t0_r4_c2_rr2 + t0_r4_c2_rr3;
  assign t1_r4_c2_rr2 = t0_r4_c2_rr4 + t0_r4_c2_rr5;
  assign t1_r4_c2_rr3 = t0_r4_c2_rr6 + t0_r4_c2_rr7;
  assign t1_r4_c2_rr4 = t0_r4_c2_rr8 + t0_r4_c2_rr9;

  assign t2_r4_c2_rr0 = t1_r4_c2_rr0 + t1_r4_c2_rr1;
  assign t2_r4_c2_rr1 = t1_r4_c2_rr2 + t1_r4_c2_rr3;
  assign t2_r4_c2_rr2 = t1_r4_c2_rr4;

  assign t3_r4_c2_rr0 = t2_r4_c2_rr0 + t2_r4_c2_rr1;
  assign t3_r4_c2_rr1 = t2_r4_c2_rr2;

  assign t4_r4_c2_rr0 = t3_r4_c2_rr0 + t3_r4_c2_rr1;

  assign c_4_2 = t4_r4_c2_rr0;
  assign t0_r4_c3_rr0 = a_4_0 * b_0_3;
  assign t0_r4_c3_rr1 = a_4_1 * b_1_3;
  assign t0_r4_c3_rr2 = a_4_2 * b_2_3;
  assign t0_r4_c3_rr3 = a_4_3 * b_3_3;
  assign t0_r4_c3_rr4 = a_4_4 * b_4_3;
  assign t0_r4_c3_rr5 = a_4_5 * b_5_3;
  assign t0_r4_c3_rr6 = a_4_6 * b_6_3;
  assign t0_r4_c3_rr7 = a_4_7 * b_7_3;
  assign t0_r4_c3_rr8 = a_4_8 * b_8_3;
  assign t0_r4_c3_rr9 = a_4_9 * b_9_3;
  assign t1_r4_c3_rr0 = t0_r4_c3_rr0 + t0_r4_c3_rr1;
  assign t1_r4_c3_rr1 = t0_r4_c3_rr2 + t0_r4_c3_rr3;
  assign t1_r4_c3_rr2 = t0_r4_c3_rr4 + t0_r4_c3_rr5;
  assign t1_r4_c3_rr3 = t0_r4_c3_rr6 + t0_r4_c3_rr7;
  assign t1_r4_c3_rr4 = t0_r4_c3_rr8 + t0_r4_c3_rr9;

  assign t2_r4_c3_rr0 = t1_r4_c3_rr0 + t1_r4_c3_rr1;
  assign t2_r4_c3_rr1 = t1_r4_c3_rr2 + t1_r4_c3_rr3;
  assign t2_r4_c3_rr2 = t1_r4_c3_rr4;

  assign t3_r4_c3_rr0 = t2_r4_c3_rr0 + t2_r4_c3_rr1;
  assign t3_r4_c3_rr1 = t2_r4_c3_rr2;

  assign t4_r4_c3_rr0 = t3_r4_c3_rr0 + t3_r4_c3_rr1;

  assign c_4_3 = t4_r4_c3_rr0;
  assign t0_r4_c4_rr0 = a_4_0 * b_0_4;
  assign t0_r4_c4_rr1 = a_4_1 * b_1_4;
  assign t0_r4_c4_rr2 = a_4_2 * b_2_4;
  assign t0_r4_c4_rr3 = a_4_3 * b_3_4;
  assign t0_r4_c4_rr4 = a_4_4 * b_4_4;
  assign t0_r4_c4_rr5 = a_4_5 * b_5_4;
  assign t0_r4_c4_rr6 = a_4_6 * b_6_4;
  assign t0_r4_c4_rr7 = a_4_7 * b_7_4;
  assign t0_r4_c4_rr8 = a_4_8 * b_8_4;
  assign t0_r4_c4_rr9 = a_4_9 * b_9_4;
  assign t1_r4_c4_rr0 = t0_r4_c4_rr0 + t0_r4_c4_rr1;
  assign t1_r4_c4_rr1 = t0_r4_c4_rr2 + t0_r4_c4_rr3;
  assign t1_r4_c4_rr2 = t0_r4_c4_rr4 + t0_r4_c4_rr5;
  assign t1_r4_c4_rr3 = t0_r4_c4_rr6 + t0_r4_c4_rr7;
  assign t1_r4_c4_rr4 = t0_r4_c4_rr8 + t0_r4_c4_rr9;

  assign t2_r4_c4_rr0 = t1_r4_c4_rr0 + t1_r4_c4_rr1;
  assign t2_r4_c4_rr1 = t1_r4_c4_rr2 + t1_r4_c4_rr3;
  assign t2_r4_c4_rr2 = t1_r4_c4_rr4;

  assign t3_r4_c4_rr0 = t2_r4_c4_rr0 + t2_r4_c4_rr1;
  assign t3_r4_c4_rr1 = t2_r4_c4_rr2;

  assign t4_r4_c4_rr0 = t3_r4_c4_rr0 + t3_r4_c4_rr1;

  assign c_4_4 = t4_r4_c4_rr0;
  assign t0_r4_c5_rr0 = a_4_0 * b_0_5;
  assign t0_r4_c5_rr1 = a_4_1 * b_1_5;
  assign t0_r4_c5_rr2 = a_4_2 * b_2_5;
  assign t0_r4_c5_rr3 = a_4_3 * b_3_5;
  assign t0_r4_c5_rr4 = a_4_4 * b_4_5;
  assign t0_r4_c5_rr5 = a_4_5 * b_5_5;
  assign t0_r4_c5_rr6 = a_4_6 * b_6_5;
  assign t0_r4_c5_rr7 = a_4_7 * b_7_5;
  assign t0_r4_c5_rr8 = a_4_8 * b_8_5;
  assign t0_r4_c5_rr9 = a_4_9 * b_9_5;
  assign t1_r4_c5_rr0 = t0_r4_c5_rr0 + t0_r4_c5_rr1;
  assign t1_r4_c5_rr1 = t0_r4_c5_rr2 + t0_r4_c5_rr3;
  assign t1_r4_c5_rr2 = t0_r4_c5_rr4 + t0_r4_c5_rr5;
  assign t1_r4_c5_rr3 = t0_r4_c5_rr6 + t0_r4_c5_rr7;
  assign t1_r4_c5_rr4 = t0_r4_c5_rr8 + t0_r4_c5_rr9;

  assign t2_r4_c5_rr0 = t1_r4_c5_rr0 + t1_r4_c5_rr1;
  assign t2_r4_c5_rr1 = t1_r4_c5_rr2 + t1_r4_c5_rr3;
  assign t2_r4_c5_rr2 = t1_r4_c5_rr4;

  assign t3_r4_c5_rr0 = t2_r4_c5_rr0 + t2_r4_c5_rr1;
  assign t3_r4_c5_rr1 = t2_r4_c5_rr2;

  assign t4_r4_c5_rr0 = t3_r4_c5_rr0 + t3_r4_c5_rr1;

  assign c_4_5 = t4_r4_c5_rr0;
  assign t0_r4_c6_rr0 = a_4_0 * b_0_6;
  assign t0_r4_c6_rr1 = a_4_1 * b_1_6;
  assign t0_r4_c6_rr2 = a_4_2 * b_2_6;
  assign t0_r4_c6_rr3 = a_4_3 * b_3_6;
  assign t0_r4_c6_rr4 = a_4_4 * b_4_6;
  assign t0_r4_c6_rr5 = a_4_5 * b_5_6;
  assign t0_r4_c6_rr6 = a_4_6 * b_6_6;
  assign t0_r4_c6_rr7 = a_4_7 * b_7_6;
  assign t0_r4_c6_rr8 = a_4_8 * b_8_6;
  assign t0_r4_c6_rr9 = a_4_9 * b_9_6;
  assign t1_r4_c6_rr0 = t0_r4_c6_rr0 + t0_r4_c6_rr1;
  assign t1_r4_c6_rr1 = t0_r4_c6_rr2 + t0_r4_c6_rr3;
  assign t1_r4_c6_rr2 = t0_r4_c6_rr4 + t0_r4_c6_rr5;
  assign t1_r4_c6_rr3 = t0_r4_c6_rr6 + t0_r4_c6_rr7;
  assign t1_r4_c6_rr4 = t0_r4_c6_rr8 + t0_r4_c6_rr9;

  assign t2_r4_c6_rr0 = t1_r4_c6_rr0 + t1_r4_c6_rr1;
  assign t2_r4_c6_rr1 = t1_r4_c6_rr2 + t1_r4_c6_rr3;
  assign t2_r4_c6_rr2 = t1_r4_c6_rr4;

  assign t3_r4_c6_rr0 = t2_r4_c6_rr0 + t2_r4_c6_rr1;
  assign t3_r4_c6_rr1 = t2_r4_c6_rr2;

  assign t4_r4_c6_rr0 = t3_r4_c6_rr0 + t3_r4_c6_rr1;

  assign c_4_6 = t4_r4_c6_rr0;
  assign t0_r4_c7_rr0 = a_4_0 * b_0_7;
  assign t0_r4_c7_rr1 = a_4_1 * b_1_7;
  assign t0_r4_c7_rr2 = a_4_2 * b_2_7;
  assign t0_r4_c7_rr3 = a_4_3 * b_3_7;
  assign t0_r4_c7_rr4 = a_4_4 * b_4_7;
  assign t0_r4_c7_rr5 = a_4_5 * b_5_7;
  assign t0_r4_c7_rr6 = a_4_6 * b_6_7;
  assign t0_r4_c7_rr7 = a_4_7 * b_7_7;
  assign t0_r4_c7_rr8 = a_4_8 * b_8_7;
  assign t0_r4_c7_rr9 = a_4_9 * b_9_7;
  assign t1_r4_c7_rr0 = t0_r4_c7_rr0 + t0_r4_c7_rr1;
  assign t1_r4_c7_rr1 = t0_r4_c7_rr2 + t0_r4_c7_rr3;
  assign t1_r4_c7_rr2 = t0_r4_c7_rr4 + t0_r4_c7_rr5;
  assign t1_r4_c7_rr3 = t0_r4_c7_rr6 + t0_r4_c7_rr7;
  assign t1_r4_c7_rr4 = t0_r4_c7_rr8 + t0_r4_c7_rr9;

  assign t2_r4_c7_rr0 = t1_r4_c7_rr0 + t1_r4_c7_rr1;
  assign t2_r4_c7_rr1 = t1_r4_c7_rr2 + t1_r4_c7_rr3;
  assign t2_r4_c7_rr2 = t1_r4_c7_rr4;

  assign t3_r4_c7_rr0 = t2_r4_c7_rr0 + t2_r4_c7_rr1;
  assign t3_r4_c7_rr1 = t2_r4_c7_rr2;

  assign t4_r4_c7_rr0 = t3_r4_c7_rr0 + t3_r4_c7_rr1;

  assign c_4_7 = t4_r4_c7_rr0;
  assign t0_r4_c8_rr0 = a_4_0 * b_0_8;
  assign t0_r4_c8_rr1 = a_4_1 * b_1_8;
  assign t0_r4_c8_rr2 = a_4_2 * b_2_8;
  assign t0_r4_c8_rr3 = a_4_3 * b_3_8;
  assign t0_r4_c8_rr4 = a_4_4 * b_4_8;
  assign t0_r4_c8_rr5 = a_4_5 * b_5_8;
  assign t0_r4_c8_rr6 = a_4_6 * b_6_8;
  assign t0_r4_c8_rr7 = a_4_7 * b_7_8;
  assign t0_r4_c8_rr8 = a_4_8 * b_8_8;
  assign t0_r4_c8_rr9 = a_4_9 * b_9_8;
  assign t1_r4_c8_rr0 = t0_r4_c8_rr0 + t0_r4_c8_rr1;
  assign t1_r4_c8_rr1 = t0_r4_c8_rr2 + t0_r4_c8_rr3;
  assign t1_r4_c8_rr2 = t0_r4_c8_rr4 + t0_r4_c8_rr5;
  assign t1_r4_c8_rr3 = t0_r4_c8_rr6 + t0_r4_c8_rr7;
  assign t1_r4_c8_rr4 = t0_r4_c8_rr8 + t0_r4_c8_rr9;

  assign t2_r4_c8_rr0 = t1_r4_c8_rr0 + t1_r4_c8_rr1;
  assign t2_r4_c8_rr1 = t1_r4_c8_rr2 + t1_r4_c8_rr3;
  assign t2_r4_c8_rr2 = t1_r4_c8_rr4;

  assign t3_r4_c8_rr0 = t2_r4_c8_rr0 + t2_r4_c8_rr1;
  assign t3_r4_c8_rr1 = t2_r4_c8_rr2;

  assign t4_r4_c8_rr0 = t3_r4_c8_rr0 + t3_r4_c8_rr1;

  assign c_4_8 = t4_r4_c8_rr0;
  assign t0_r4_c9_rr0 = a_4_0 * b_0_9;
  assign t0_r4_c9_rr1 = a_4_1 * b_1_9;
  assign t0_r4_c9_rr2 = a_4_2 * b_2_9;
  assign t0_r4_c9_rr3 = a_4_3 * b_3_9;
  assign t0_r4_c9_rr4 = a_4_4 * b_4_9;
  assign t0_r4_c9_rr5 = a_4_5 * b_5_9;
  assign t0_r4_c9_rr6 = a_4_6 * b_6_9;
  assign t0_r4_c9_rr7 = a_4_7 * b_7_9;
  assign t0_r4_c9_rr8 = a_4_8 * b_8_9;
  assign t0_r4_c9_rr9 = a_4_9 * b_9_9;
  assign t1_r4_c9_rr0 = t0_r4_c9_rr0 + t0_r4_c9_rr1;
  assign t1_r4_c9_rr1 = t0_r4_c9_rr2 + t0_r4_c9_rr3;
  assign t1_r4_c9_rr2 = t0_r4_c9_rr4 + t0_r4_c9_rr5;
  assign t1_r4_c9_rr3 = t0_r4_c9_rr6 + t0_r4_c9_rr7;
  assign t1_r4_c9_rr4 = t0_r4_c9_rr8 + t0_r4_c9_rr9;

  assign t2_r4_c9_rr0 = t1_r4_c9_rr0 + t1_r4_c9_rr1;
  assign t2_r4_c9_rr1 = t1_r4_c9_rr2 + t1_r4_c9_rr3;
  assign t2_r4_c9_rr2 = t1_r4_c9_rr4;

  assign t3_r4_c9_rr0 = t2_r4_c9_rr0 + t2_r4_c9_rr1;
  assign t3_r4_c9_rr1 = t2_r4_c9_rr2;

  assign t4_r4_c9_rr0 = t3_r4_c9_rr0 + t3_r4_c9_rr1;

  assign c_4_9 = t4_r4_c9_rr0;
  assign t0_r5_c0_rr0 = a_5_0 * b_0_0;
  assign t0_r5_c0_rr1 = a_5_1 * b_1_0;
  assign t0_r5_c0_rr2 = a_5_2 * b_2_0;
  assign t0_r5_c0_rr3 = a_5_3 * b_3_0;
  assign t0_r5_c0_rr4 = a_5_4 * b_4_0;
  assign t0_r5_c0_rr5 = a_5_5 * b_5_0;
  assign t0_r5_c0_rr6 = a_5_6 * b_6_0;
  assign t0_r5_c0_rr7 = a_5_7 * b_7_0;
  assign t0_r5_c0_rr8 = a_5_8 * b_8_0;
  assign t0_r5_c0_rr9 = a_5_9 * b_9_0;
  assign t1_r5_c0_rr0 = t0_r5_c0_rr0 + t0_r5_c0_rr1;
  assign t1_r5_c0_rr1 = t0_r5_c0_rr2 + t0_r5_c0_rr3;
  assign t1_r5_c0_rr2 = t0_r5_c0_rr4 + t0_r5_c0_rr5;
  assign t1_r5_c0_rr3 = t0_r5_c0_rr6 + t0_r5_c0_rr7;
  assign t1_r5_c0_rr4 = t0_r5_c0_rr8 + t0_r5_c0_rr9;

  assign t2_r5_c0_rr0 = t1_r5_c0_rr0 + t1_r5_c0_rr1;
  assign t2_r5_c0_rr1 = t1_r5_c0_rr2 + t1_r5_c0_rr3;
  assign t2_r5_c0_rr2 = t1_r5_c0_rr4;

  assign t3_r5_c0_rr0 = t2_r5_c0_rr0 + t2_r5_c0_rr1;
  assign t3_r5_c0_rr1 = t2_r5_c0_rr2;

  assign t4_r5_c0_rr0 = t3_r5_c0_rr0 + t3_r5_c0_rr1;

  assign c_5_0 = t4_r5_c0_rr0;
  assign t0_r5_c1_rr0 = a_5_0 * b_0_1;
  assign t0_r5_c1_rr1 = a_5_1 * b_1_1;
  assign t0_r5_c1_rr2 = a_5_2 * b_2_1;
  assign t0_r5_c1_rr3 = a_5_3 * b_3_1;
  assign t0_r5_c1_rr4 = a_5_4 * b_4_1;
  assign t0_r5_c1_rr5 = a_5_5 * b_5_1;
  assign t0_r5_c1_rr6 = a_5_6 * b_6_1;
  assign t0_r5_c1_rr7 = a_5_7 * b_7_1;
  assign t0_r5_c1_rr8 = a_5_8 * b_8_1;
  assign t0_r5_c1_rr9 = a_5_9 * b_9_1;
  assign t1_r5_c1_rr0 = t0_r5_c1_rr0 + t0_r5_c1_rr1;
  assign t1_r5_c1_rr1 = t0_r5_c1_rr2 + t0_r5_c1_rr3;
  assign t1_r5_c1_rr2 = t0_r5_c1_rr4 + t0_r5_c1_rr5;
  assign t1_r5_c1_rr3 = t0_r5_c1_rr6 + t0_r5_c1_rr7;
  assign t1_r5_c1_rr4 = t0_r5_c1_rr8 + t0_r5_c1_rr9;

  assign t2_r5_c1_rr0 = t1_r5_c1_rr0 + t1_r5_c1_rr1;
  assign t2_r5_c1_rr1 = t1_r5_c1_rr2 + t1_r5_c1_rr3;
  assign t2_r5_c1_rr2 = t1_r5_c1_rr4;

  assign t3_r5_c1_rr0 = t2_r5_c1_rr0 + t2_r5_c1_rr1;
  assign t3_r5_c1_rr1 = t2_r5_c1_rr2;

  assign t4_r5_c1_rr0 = t3_r5_c1_rr0 + t3_r5_c1_rr1;

  assign c_5_1 = t4_r5_c1_rr0;
  assign t0_r5_c2_rr0 = a_5_0 * b_0_2;
  assign t0_r5_c2_rr1 = a_5_1 * b_1_2;
  assign t0_r5_c2_rr2 = a_5_2 * b_2_2;
  assign t0_r5_c2_rr3 = a_5_3 * b_3_2;
  assign t0_r5_c2_rr4 = a_5_4 * b_4_2;
  assign t0_r5_c2_rr5 = a_5_5 * b_5_2;
  assign t0_r5_c2_rr6 = a_5_6 * b_6_2;
  assign t0_r5_c2_rr7 = a_5_7 * b_7_2;
  assign t0_r5_c2_rr8 = a_5_8 * b_8_2;
  assign t0_r5_c2_rr9 = a_5_9 * b_9_2;
  assign t1_r5_c2_rr0 = t0_r5_c2_rr0 + t0_r5_c2_rr1;
  assign t1_r5_c2_rr1 = t0_r5_c2_rr2 + t0_r5_c2_rr3;
  assign t1_r5_c2_rr2 = t0_r5_c2_rr4 + t0_r5_c2_rr5;
  assign t1_r5_c2_rr3 = t0_r5_c2_rr6 + t0_r5_c2_rr7;
  assign t1_r5_c2_rr4 = t0_r5_c2_rr8 + t0_r5_c2_rr9;

  assign t2_r5_c2_rr0 = t1_r5_c2_rr0 + t1_r5_c2_rr1;
  assign t2_r5_c2_rr1 = t1_r5_c2_rr2 + t1_r5_c2_rr3;
  assign t2_r5_c2_rr2 = t1_r5_c2_rr4;

  assign t3_r5_c2_rr0 = t2_r5_c2_rr0 + t2_r5_c2_rr1;
  assign t3_r5_c2_rr1 = t2_r5_c2_rr2;

  assign t4_r5_c2_rr0 = t3_r5_c2_rr0 + t3_r5_c2_rr1;

  assign c_5_2 = t4_r5_c2_rr0;
  assign t0_r5_c3_rr0 = a_5_0 * b_0_3;
  assign t0_r5_c3_rr1 = a_5_1 * b_1_3;
  assign t0_r5_c3_rr2 = a_5_2 * b_2_3;
  assign t0_r5_c3_rr3 = a_5_3 * b_3_3;
  assign t0_r5_c3_rr4 = a_5_4 * b_4_3;
  assign t0_r5_c3_rr5 = a_5_5 * b_5_3;
  assign t0_r5_c3_rr6 = a_5_6 * b_6_3;
  assign t0_r5_c3_rr7 = a_5_7 * b_7_3;
  assign t0_r5_c3_rr8 = a_5_8 * b_8_3;
  assign t0_r5_c3_rr9 = a_5_9 * b_9_3;
  assign t1_r5_c3_rr0 = t0_r5_c3_rr0 + t0_r5_c3_rr1;
  assign t1_r5_c3_rr1 = t0_r5_c3_rr2 + t0_r5_c3_rr3;
  assign t1_r5_c3_rr2 = t0_r5_c3_rr4 + t0_r5_c3_rr5;
  assign t1_r5_c3_rr3 = t0_r5_c3_rr6 + t0_r5_c3_rr7;
  assign t1_r5_c3_rr4 = t0_r5_c3_rr8 + t0_r5_c3_rr9;

  assign t2_r5_c3_rr0 = t1_r5_c3_rr0 + t1_r5_c3_rr1;
  assign t2_r5_c3_rr1 = t1_r5_c3_rr2 + t1_r5_c3_rr3;
  assign t2_r5_c3_rr2 = t1_r5_c3_rr4;

  assign t3_r5_c3_rr0 = t2_r5_c3_rr0 + t2_r5_c3_rr1;
  assign t3_r5_c3_rr1 = t2_r5_c3_rr2;

  assign t4_r5_c3_rr0 = t3_r5_c3_rr0 + t3_r5_c3_rr1;

  assign c_5_3 = t4_r5_c3_rr0;
  assign t0_r5_c4_rr0 = a_5_0 * b_0_4;
  assign t0_r5_c4_rr1 = a_5_1 * b_1_4;
  assign t0_r5_c4_rr2 = a_5_2 * b_2_4;
  assign t0_r5_c4_rr3 = a_5_3 * b_3_4;
  assign t0_r5_c4_rr4 = a_5_4 * b_4_4;
  assign t0_r5_c4_rr5 = a_5_5 * b_5_4;
  assign t0_r5_c4_rr6 = a_5_6 * b_6_4;
  assign t0_r5_c4_rr7 = a_5_7 * b_7_4;
  assign t0_r5_c4_rr8 = a_5_8 * b_8_4;
  assign t0_r5_c4_rr9 = a_5_9 * b_9_4;
  assign t1_r5_c4_rr0 = t0_r5_c4_rr0 + t0_r5_c4_rr1;
  assign t1_r5_c4_rr1 = t0_r5_c4_rr2 + t0_r5_c4_rr3;
  assign t1_r5_c4_rr2 = t0_r5_c4_rr4 + t0_r5_c4_rr5;
  assign t1_r5_c4_rr3 = t0_r5_c4_rr6 + t0_r5_c4_rr7;
  assign t1_r5_c4_rr4 = t0_r5_c4_rr8 + t0_r5_c4_rr9;

  assign t2_r5_c4_rr0 = t1_r5_c4_rr0 + t1_r5_c4_rr1;
  assign t2_r5_c4_rr1 = t1_r5_c4_rr2 + t1_r5_c4_rr3;
  assign t2_r5_c4_rr2 = t1_r5_c4_rr4;

  assign t3_r5_c4_rr0 = t2_r5_c4_rr0 + t2_r5_c4_rr1;
  assign t3_r5_c4_rr1 = t2_r5_c4_rr2;

  assign t4_r5_c4_rr0 = t3_r5_c4_rr0 + t3_r5_c4_rr1;

  assign c_5_4 = t4_r5_c4_rr0;
  assign t0_r5_c5_rr0 = a_5_0 * b_0_5;
  assign t0_r5_c5_rr1 = a_5_1 * b_1_5;
  assign t0_r5_c5_rr2 = a_5_2 * b_2_5;
  assign t0_r5_c5_rr3 = a_5_3 * b_3_5;
  assign t0_r5_c5_rr4 = a_5_4 * b_4_5;
  assign t0_r5_c5_rr5 = a_5_5 * b_5_5;
  assign t0_r5_c5_rr6 = a_5_6 * b_6_5;
  assign t0_r5_c5_rr7 = a_5_7 * b_7_5;
  assign t0_r5_c5_rr8 = a_5_8 * b_8_5;
  assign t0_r5_c5_rr9 = a_5_9 * b_9_5;
  assign t1_r5_c5_rr0 = t0_r5_c5_rr0 + t0_r5_c5_rr1;
  assign t1_r5_c5_rr1 = t0_r5_c5_rr2 + t0_r5_c5_rr3;
  assign t1_r5_c5_rr2 = t0_r5_c5_rr4 + t0_r5_c5_rr5;
  assign t1_r5_c5_rr3 = t0_r5_c5_rr6 + t0_r5_c5_rr7;
  assign t1_r5_c5_rr4 = t0_r5_c5_rr8 + t0_r5_c5_rr9;

  assign t2_r5_c5_rr0 = t1_r5_c5_rr0 + t1_r5_c5_rr1;
  assign t2_r5_c5_rr1 = t1_r5_c5_rr2 + t1_r5_c5_rr3;
  assign t2_r5_c5_rr2 = t1_r5_c5_rr4;

  assign t3_r5_c5_rr0 = t2_r5_c5_rr0 + t2_r5_c5_rr1;
  assign t3_r5_c5_rr1 = t2_r5_c5_rr2;

  assign t4_r5_c5_rr0 = t3_r5_c5_rr0 + t3_r5_c5_rr1;

  assign c_5_5 = t4_r5_c5_rr0;
  assign t0_r5_c6_rr0 = a_5_0 * b_0_6;
  assign t0_r5_c6_rr1 = a_5_1 * b_1_6;
  assign t0_r5_c6_rr2 = a_5_2 * b_2_6;
  assign t0_r5_c6_rr3 = a_5_3 * b_3_6;
  assign t0_r5_c6_rr4 = a_5_4 * b_4_6;
  assign t0_r5_c6_rr5 = a_5_5 * b_5_6;
  assign t0_r5_c6_rr6 = a_5_6 * b_6_6;
  assign t0_r5_c6_rr7 = a_5_7 * b_7_6;
  assign t0_r5_c6_rr8 = a_5_8 * b_8_6;
  assign t0_r5_c6_rr9 = a_5_9 * b_9_6;
  assign t1_r5_c6_rr0 = t0_r5_c6_rr0 + t0_r5_c6_rr1;
  assign t1_r5_c6_rr1 = t0_r5_c6_rr2 + t0_r5_c6_rr3;
  assign t1_r5_c6_rr2 = t0_r5_c6_rr4 + t0_r5_c6_rr5;
  assign t1_r5_c6_rr3 = t0_r5_c6_rr6 + t0_r5_c6_rr7;
  assign t1_r5_c6_rr4 = t0_r5_c6_rr8 + t0_r5_c6_rr9;

  assign t2_r5_c6_rr0 = t1_r5_c6_rr0 + t1_r5_c6_rr1;
  assign t2_r5_c6_rr1 = t1_r5_c6_rr2 + t1_r5_c6_rr3;
  assign t2_r5_c6_rr2 = t1_r5_c6_rr4;

  assign t3_r5_c6_rr0 = t2_r5_c6_rr0 + t2_r5_c6_rr1;
  assign t3_r5_c6_rr1 = t2_r5_c6_rr2;

  assign t4_r5_c6_rr0 = t3_r5_c6_rr0 + t3_r5_c6_rr1;

  assign c_5_6 = t4_r5_c6_rr0;
  assign t0_r5_c7_rr0 = a_5_0 * b_0_7;
  assign t0_r5_c7_rr1 = a_5_1 * b_1_7;
  assign t0_r5_c7_rr2 = a_5_2 * b_2_7;
  assign t0_r5_c7_rr3 = a_5_3 * b_3_7;
  assign t0_r5_c7_rr4 = a_5_4 * b_4_7;
  assign t0_r5_c7_rr5 = a_5_5 * b_5_7;
  assign t0_r5_c7_rr6 = a_5_6 * b_6_7;
  assign t0_r5_c7_rr7 = a_5_7 * b_7_7;
  assign t0_r5_c7_rr8 = a_5_8 * b_8_7;
  assign t0_r5_c7_rr9 = a_5_9 * b_9_7;
  assign t1_r5_c7_rr0 = t0_r5_c7_rr0 + t0_r5_c7_rr1;
  assign t1_r5_c7_rr1 = t0_r5_c7_rr2 + t0_r5_c7_rr3;
  assign t1_r5_c7_rr2 = t0_r5_c7_rr4 + t0_r5_c7_rr5;
  assign t1_r5_c7_rr3 = t0_r5_c7_rr6 + t0_r5_c7_rr7;
  assign t1_r5_c7_rr4 = t0_r5_c7_rr8 + t0_r5_c7_rr9;

  assign t2_r5_c7_rr0 = t1_r5_c7_rr0 + t1_r5_c7_rr1;
  assign t2_r5_c7_rr1 = t1_r5_c7_rr2 + t1_r5_c7_rr3;
  assign t2_r5_c7_rr2 = t1_r5_c7_rr4;

  assign t3_r5_c7_rr0 = t2_r5_c7_rr0 + t2_r5_c7_rr1;
  assign t3_r5_c7_rr1 = t2_r5_c7_rr2;

  assign t4_r5_c7_rr0 = t3_r5_c7_rr0 + t3_r5_c7_rr1;

  assign c_5_7 = t4_r5_c7_rr0;
  assign t0_r5_c8_rr0 = a_5_0 * b_0_8;
  assign t0_r5_c8_rr1 = a_5_1 * b_1_8;
  assign t0_r5_c8_rr2 = a_5_2 * b_2_8;
  assign t0_r5_c8_rr3 = a_5_3 * b_3_8;
  assign t0_r5_c8_rr4 = a_5_4 * b_4_8;
  assign t0_r5_c8_rr5 = a_5_5 * b_5_8;
  assign t0_r5_c8_rr6 = a_5_6 * b_6_8;
  assign t0_r5_c8_rr7 = a_5_7 * b_7_8;
  assign t0_r5_c8_rr8 = a_5_8 * b_8_8;
  assign t0_r5_c8_rr9 = a_5_9 * b_9_8;
  assign t1_r5_c8_rr0 = t0_r5_c8_rr0 + t0_r5_c8_rr1;
  assign t1_r5_c8_rr1 = t0_r5_c8_rr2 + t0_r5_c8_rr3;
  assign t1_r5_c8_rr2 = t0_r5_c8_rr4 + t0_r5_c8_rr5;
  assign t1_r5_c8_rr3 = t0_r5_c8_rr6 + t0_r5_c8_rr7;
  assign t1_r5_c8_rr4 = t0_r5_c8_rr8 + t0_r5_c8_rr9;

  assign t2_r5_c8_rr0 = t1_r5_c8_rr0 + t1_r5_c8_rr1;
  assign t2_r5_c8_rr1 = t1_r5_c8_rr2 + t1_r5_c8_rr3;
  assign t2_r5_c8_rr2 = t1_r5_c8_rr4;

  assign t3_r5_c8_rr0 = t2_r5_c8_rr0 + t2_r5_c8_rr1;
  assign t3_r5_c8_rr1 = t2_r5_c8_rr2;

  assign t4_r5_c8_rr0 = t3_r5_c8_rr0 + t3_r5_c8_rr1;

  assign c_5_8 = t4_r5_c8_rr0;
  assign t0_r5_c9_rr0 = a_5_0 * b_0_9;
  assign t0_r5_c9_rr1 = a_5_1 * b_1_9;
  assign t0_r5_c9_rr2 = a_5_2 * b_2_9;
  assign t0_r5_c9_rr3 = a_5_3 * b_3_9;
  assign t0_r5_c9_rr4 = a_5_4 * b_4_9;
  assign t0_r5_c9_rr5 = a_5_5 * b_5_9;
  assign t0_r5_c9_rr6 = a_5_6 * b_6_9;
  assign t0_r5_c9_rr7 = a_5_7 * b_7_9;
  assign t0_r5_c9_rr8 = a_5_8 * b_8_9;
  assign t0_r5_c9_rr9 = a_5_9 * b_9_9;
  assign t1_r5_c9_rr0 = t0_r5_c9_rr0 + t0_r5_c9_rr1;
  assign t1_r5_c9_rr1 = t0_r5_c9_rr2 + t0_r5_c9_rr3;
  assign t1_r5_c9_rr2 = t0_r5_c9_rr4 + t0_r5_c9_rr5;
  assign t1_r5_c9_rr3 = t0_r5_c9_rr6 + t0_r5_c9_rr7;
  assign t1_r5_c9_rr4 = t0_r5_c9_rr8 + t0_r5_c9_rr9;

  assign t2_r5_c9_rr0 = t1_r5_c9_rr0 + t1_r5_c9_rr1;
  assign t2_r5_c9_rr1 = t1_r5_c9_rr2 + t1_r5_c9_rr3;
  assign t2_r5_c9_rr2 = t1_r5_c9_rr4;

  assign t3_r5_c9_rr0 = t2_r5_c9_rr0 + t2_r5_c9_rr1;
  assign t3_r5_c9_rr1 = t2_r5_c9_rr2;

  assign t4_r5_c9_rr0 = t3_r5_c9_rr0 + t3_r5_c9_rr1;

  assign c_5_9 = t4_r5_c9_rr0;
  assign t0_r6_c0_rr0 = a_6_0 * b_0_0;
  assign t0_r6_c0_rr1 = a_6_1 * b_1_0;
  assign t0_r6_c0_rr2 = a_6_2 * b_2_0;
  assign t0_r6_c0_rr3 = a_6_3 * b_3_0;
  assign t0_r6_c0_rr4 = a_6_4 * b_4_0;
  assign t0_r6_c0_rr5 = a_6_5 * b_5_0;
  assign t0_r6_c0_rr6 = a_6_6 * b_6_0;
  assign t0_r6_c0_rr7 = a_6_7 * b_7_0;
  assign t0_r6_c0_rr8 = a_6_8 * b_8_0;
  assign t0_r6_c0_rr9 = a_6_9 * b_9_0;
  assign t1_r6_c0_rr0 = t0_r6_c0_rr0 + t0_r6_c0_rr1;
  assign t1_r6_c0_rr1 = t0_r6_c0_rr2 + t0_r6_c0_rr3;
  assign t1_r6_c0_rr2 = t0_r6_c0_rr4 + t0_r6_c0_rr5;
  assign t1_r6_c0_rr3 = t0_r6_c0_rr6 + t0_r6_c0_rr7;
  assign t1_r6_c0_rr4 = t0_r6_c0_rr8 + t0_r6_c0_rr9;

  assign t2_r6_c0_rr0 = t1_r6_c0_rr0 + t1_r6_c0_rr1;
  assign t2_r6_c0_rr1 = t1_r6_c0_rr2 + t1_r6_c0_rr3;
  assign t2_r6_c0_rr2 = t1_r6_c0_rr4;

  assign t3_r6_c0_rr0 = t2_r6_c0_rr0 + t2_r6_c0_rr1;
  assign t3_r6_c0_rr1 = t2_r6_c0_rr2;

  assign t4_r6_c0_rr0 = t3_r6_c0_rr0 + t3_r6_c0_rr1;

  assign c_6_0 = t4_r6_c0_rr0;
  assign t0_r6_c1_rr0 = a_6_0 * b_0_1;
  assign t0_r6_c1_rr1 = a_6_1 * b_1_1;
  assign t0_r6_c1_rr2 = a_6_2 * b_2_1;
  assign t0_r6_c1_rr3 = a_6_3 * b_3_1;
  assign t0_r6_c1_rr4 = a_6_4 * b_4_1;
  assign t0_r6_c1_rr5 = a_6_5 * b_5_1;
  assign t0_r6_c1_rr6 = a_6_6 * b_6_1;
  assign t0_r6_c1_rr7 = a_6_7 * b_7_1;
  assign t0_r6_c1_rr8 = a_6_8 * b_8_1;
  assign t0_r6_c1_rr9 = a_6_9 * b_9_1;
  assign t1_r6_c1_rr0 = t0_r6_c1_rr0 + t0_r6_c1_rr1;
  assign t1_r6_c1_rr1 = t0_r6_c1_rr2 + t0_r6_c1_rr3;
  assign t1_r6_c1_rr2 = t0_r6_c1_rr4 + t0_r6_c1_rr5;
  assign t1_r6_c1_rr3 = t0_r6_c1_rr6 + t0_r6_c1_rr7;
  assign t1_r6_c1_rr4 = t0_r6_c1_rr8 + t0_r6_c1_rr9;

  assign t2_r6_c1_rr0 = t1_r6_c1_rr0 + t1_r6_c1_rr1;
  assign t2_r6_c1_rr1 = t1_r6_c1_rr2 + t1_r6_c1_rr3;
  assign t2_r6_c1_rr2 = t1_r6_c1_rr4;

  assign t3_r6_c1_rr0 = t2_r6_c1_rr0 + t2_r6_c1_rr1;
  assign t3_r6_c1_rr1 = t2_r6_c1_rr2;

  assign t4_r6_c1_rr0 = t3_r6_c1_rr0 + t3_r6_c1_rr1;

  assign c_6_1 = t4_r6_c1_rr0;
  assign t0_r6_c2_rr0 = a_6_0 * b_0_2;
  assign t0_r6_c2_rr1 = a_6_1 * b_1_2;
  assign t0_r6_c2_rr2 = a_6_2 * b_2_2;
  assign t0_r6_c2_rr3 = a_6_3 * b_3_2;
  assign t0_r6_c2_rr4 = a_6_4 * b_4_2;
  assign t0_r6_c2_rr5 = a_6_5 * b_5_2;
  assign t0_r6_c2_rr6 = a_6_6 * b_6_2;
  assign t0_r6_c2_rr7 = a_6_7 * b_7_2;
  assign t0_r6_c2_rr8 = a_6_8 * b_8_2;
  assign t0_r6_c2_rr9 = a_6_9 * b_9_2;
  assign t1_r6_c2_rr0 = t0_r6_c2_rr0 + t0_r6_c2_rr1;
  assign t1_r6_c2_rr1 = t0_r6_c2_rr2 + t0_r6_c2_rr3;
  assign t1_r6_c2_rr2 = t0_r6_c2_rr4 + t0_r6_c2_rr5;
  assign t1_r6_c2_rr3 = t0_r6_c2_rr6 + t0_r6_c2_rr7;
  assign t1_r6_c2_rr4 = t0_r6_c2_rr8 + t0_r6_c2_rr9;

  assign t2_r6_c2_rr0 = t1_r6_c2_rr0 + t1_r6_c2_rr1;
  assign t2_r6_c2_rr1 = t1_r6_c2_rr2 + t1_r6_c2_rr3;
  assign t2_r6_c2_rr2 = t1_r6_c2_rr4;

  assign t3_r6_c2_rr0 = t2_r6_c2_rr0 + t2_r6_c2_rr1;
  assign t3_r6_c2_rr1 = t2_r6_c2_rr2;

  assign t4_r6_c2_rr0 = t3_r6_c2_rr0 + t3_r6_c2_rr1;

  assign c_6_2 = t4_r6_c2_rr0;
  assign t0_r6_c3_rr0 = a_6_0 * b_0_3;
  assign t0_r6_c3_rr1 = a_6_1 * b_1_3;
  assign t0_r6_c3_rr2 = a_6_2 * b_2_3;
  assign t0_r6_c3_rr3 = a_6_3 * b_3_3;
  assign t0_r6_c3_rr4 = a_6_4 * b_4_3;
  assign t0_r6_c3_rr5 = a_6_5 * b_5_3;
  assign t0_r6_c3_rr6 = a_6_6 * b_6_3;
  assign t0_r6_c3_rr7 = a_6_7 * b_7_3;
  assign t0_r6_c3_rr8 = a_6_8 * b_8_3;
  assign t0_r6_c3_rr9 = a_6_9 * b_9_3;
  assign t1_r6_c3_rr0 = t0_r6_c3_rr0 + t0_r6_c3_rr1;
  assign t1_r6_c3_rr1 = t0_r6_c3_rr2 + t0_r6_c3_rr3;
  assign t1_r6_c3_rr2 = t0_r6_c3_rr4 + t0_r6_c3_rr5;
  assign t1_r6_c3_rr3 = t0_r6_c3_rr6 + t0_r6_c3_rr7;
  assign t1_r6_c3_rr4 = t0_r6_c3_rr8 + t0_r6_c3_rr9;

  assign t2_r6_c3_rr0 = t1_r6_c3_rr0 + t1_r6_c3_rr1;
  assign t2_r6_c3_rr1 = t1_r6_c3_rr2 + t1_r6_c3_rr3;
  assign t2_r6_c3_rr2 = t1_r6_c3_rr4;

  assign t3_r6_c3_rr0 = t2_r6_c3_rr0 + t2_r6_c3_rr1;
  assign t3_r6_c3_rr1 = t2_r6_c3_rr2;

  assign t4_r6_c3_rr0 = t3_r6_c3_rr0 + t3_r6_c3_rr1;

  assign c_6_3 = t4_r6_c3_rr0;
  assign t0_r6_c4_rr0 = a_6_0 * b_0_4;
  assign t0_r6_c4_rr1 = a_6_1 * b_1_4;
  assign t0_r6_c4_rr2 = a_6_2 * b_2_4;
  assign t0_r6_c4_rr3 = a_6_3 * b_3_4;
  assign t0_r6_c4_rr4 = a_6_4 * b_4_4;
  assign t0_r6_c4_rr5 = a_6_5 * b_5_4;
  assign t0_r6_c4_rr6 = a_6_6 * b_6_4;
  assign t0_r6_c4_rr7 = a_6_7 * b_7_4;
  assign t0_r6_c4_rr8 = a_6_8 * b_8_4;
  assign t0_r6_c4_rr9 = a_6_9 * b_9_4;
  assign t1_r6_c4_rr0 = t0_r6_c4_rr0 + t0_r6_c4_rr1;
  assign t1_r6_c4_rr1 = t0_r6_c4_rr2 + t0_r6_c4_rr3;
  assign t1_r6_c4_rr2 = t0_r6_c4_rr4 + t0_r6_c4_rr5;
  assign t1_r6_c4_rr3 = t0_r6_c4_rr6 + t0_r6_c4_rr7;
  assign t1_r6_c4_rr4 = t0_r6_c4_rr8 + t0_r6_c4_rr9;

  assign t2_r6_c4_rr0 = t1_r6_c4_rr0 + t1_r6_c4_rr1;
  assign t2_r6_c4_rr1 = t1_r6_c4_rr2 + t1_r6_c4_rr3;
  assign t2_r6_c4_rr2 = t1_r6_c4_rr4;

  assign t3_r6_c4_rr0 = t2_r6_c4_rr0 + t2_r6_c4_rr1;
  assign t3_r6_c4_rr1 = t2_r6_c4_rr2;

  assign t4_r6_c4_rr0 = t3_r6_c4_rr0 + t3_r6_c4_rr1;

  assign c_6_4 = t4_r6_c4_rr0;
  assign t0_r6_c5_rr0 = a_6_0 * b_0_5;
  assign t0_r6_c5_rr1 = a_6_1 * b_1_5;
  assign t0_r6_c5_rr2 = a_6_2 * b_2_5;
  assign t0_r6_c5_rr3 = a_6_3 * b_3_5;
  assign t0_r6_c5_rr4 = a_6_4 * b_4_5;
  assign t0_r6_c5_rr5 = a_6_5 * b_5_5;
  assign t0_r6_c5_rr6 = a_6_6 * b_6_5;
  assign t0_r6_c5_rr7 = a_6_7 * b_7_5;
  assign t0_r6_c5_rr8 = a_6_8 * b_8_5;
  assign t0_r6_c5_rr9 = a_6_9 * b_9_5;
  assign t1_r6_c5_rr0 = t0_r6_c5_rr0 + t0_r6_c5_rr1;
  assign t1_r6_c5_rr1 = t0_r6_c5_rr2 + t0_r6_c5_rr3;
  assign t1_r6_c5_rr2 = t0_r6_c5_rr4 + t0_r6_c5_rr5;
  assign t1_r6_c5_rr3 = t0_r6_c5_rr6 + t0_r6_c5_rr7;
  assign t1_r6_c5_rr4 = t0_r6_c5_rr8 + t0_r6_c5_rr9;

  assign t2_r6_c5_rr0 = t1_r6_c5_rr0 + t1_r6_c5_rr1;
  assign t2_r6_c5_rr1 = t1_r6_c5_rr2 + t1_r6_c5_rr3;
  assign t2_r6_c5_rr2 = t1_r6_c5_rr4;

  assign t3_r6_c5_rr0 = t2_r6_c5_rr0 + t2_r6_c5_rr1;
  assign t3_r6_c5_rr1 = t2_r6_c5_rr2;

  assign t4_r6_c5_rr0 = t3_r6_c5_rr0 + t3_r6_c5_rr1;

  assign c_6_5 = t4_r6_c5_rr0;
  assign t0_r6_c6_rr0 = a_6_0 * b_0_6;
  assign t0_r6_c6_rr1 = a_6_1 * b_1_6;
  assign t0_r6_c6_rr2 = a_6_2 * b_2_6;
  assign t0_r6_c6_rr3 = a_6_3 * b_3_6;
  assign t0_r6_c6_rr4 = a_6_4 * b_4_6;
  assign t0_r6_c6_rr5 = a_6_5 * b_5_6;
  assign t0_r6_c6_rr6 = a_6_6 * b_6_6;
  assign t0_r6_c6_rr7 = a_6_7 * b_7_6;
  assign t0_r6_c6_rr8 = a_6_8 * b_8_6;
  assign t0_r6_c6_rr9 = a_6_9 * b_9_6;
  assign t1_r6_c6_rr0 = t0_r6_c6_rr0 + t0_r6_c6_rr1;
  assign t1_r6_c6_rr1 = t0_r6_c6_rr2 + t0_r6_c6_rr3;
  assign t1_r6_c6_rr2 = t0_r6_c6_rr4 + t0_r6_c6_rr5;
  assign t1_r6_c6_rr3 = t0_r6_c6_rr6 + t0_r6_c6_rr7;
  assign t1_r6_c6_rr4 = t0_r6_c6_rr8 + t0_r6_c6_rr9;

  assign t2_r6_c6_rr0 = t1_r6_c6_rr0 + t1_r6_c6_rr1;
  assign t2_r6_c6_rr1 = t1_r6_c6_rr2 + t1_r6_c6_rr3;
  assign t2_r6_c6_rr2 = t1_r6_c6_rr4;

  assign t3_r6_c6_rr0 = t2_r6_c6_rr0 + t2_r6_c6_rr1;
  assign t3_r6_c6_rr1 = t2_r6_c6_rr2;

  assign t4_r6_c6_rr0 = t3_r6_c6_rr0 + t3_r6_c6_rr1;

  assign c_6_6 = t4_r6_c6_rr0;
  assign t0_r6_c7_rr0 = a_6_0 * b_0_7;
  assign t0_r6_c7_rr1 = a_6_1 * b_1_7;
  assign t0_r6_c7_rr2 = a_6_2 * b_2_7;
  assign t0_r6_c7_rr3 = a_6_3 * b_3_7;
  assign t0_r6_c7_rr4 = a_6_4 * b_4_7;
  assign t0_r6_c7_rr5 = a_6_5 * b_5_7;
  assign t0_r6_c7_rr6 = a_6_6 * b_6_7;
  assign t0_r6_c7_rr7 = a_6_7 * b_7_7;
  assign t0_r6_c7_rr8 = a_6_8 * b_8_7;
  assign t0_r6_c7_rr9 = a_6_9 * b_9_7;
  assign t1_r6_c7_rr0 = t0_r6_c7_rr0 + t0_r6_c7_rr1;
  assign t1_r6_c7_rr1 = t0_r6_c7_rr2 + t0_r6_c7_rr3;
  assign t1_r6_c7_rr2 = t0_r6_c7_rr4 + t0_r6_c7_rr5;
  assign t1_r6_c7_rr3 = t0_r6_c7_rr6 + t0_r6_c7_rr7;
  assign t1_r6_c7_rr4 = t0_r6_c7_rr8 + t0_r6_c7_rr9;

  assign t2_r6_c7_rr0 = t1_r6_c7_rr0 + t1_r6_c7_rr1;
  assign t2_r6_c7_rr1 = t1_r6_c7_rr2 + t1_r6_c7_rr3;
  assign t2_r6_c7_rr2 = t1_r6_c7_rr4;

  assign t3_r6_c7_rr0 = t2_r6_c7_rr0 + t2_r6_c7_rr1;
  assign t3_r6_c7_rr1 = t2_r6_c7_rr2;

  assign t4_r6_c7_rr0 = t3_r6_c7_rr0 + t3_r6_c7_rr1;

  assign c_6_7 = t4_r6_c7_rr0;
  assign t0_r6_c8_rr0 = a_6_0 * b_0_8;
  assign t0_r6_c8_rr1 = a_6_1 * b_1_8;
  assign t0_r6_c8_rr2 = a_6_2 * b_2_8;
  assign t0_r6_c8_rr3 = a_6_3 * b_3_8;
  assign t0_r6_c8_rr4 = a_6_4 * b_4_8;
  assign t0_r6_c8_rr5 = a_6_5 * b_5_8;
  assign t0_r6_c8_rr6 = a_6_6 * b_6_8;
  assign t0_r6_c8_rr7 = a_6_7 * b_7_8;
  assign t0_r6_c8_rr8 = a_6_8 * b_8_8;
  assign t0_r6_c8_rr9 = a_6_9 * b_9_8;
  assign t1_r6_c8_rr0 = t0_r6_c8_rr0 + t0_r6_c8_rr1;
  assign t1_r6_c8_rr1 = t0_r6_c8_rr2 + t0_r6_c8_rr3;
  assign t1_r6_c8_rr2 = t0_r6_c8_rr4 + t0_r6_c8_rr5;
  assign t1_r6_c8_rr3 = t0_r6_c8_rr6 + t0_r6_c8_rr7;
  assign t1_r6_c8_rr4 = t0_r6_c8_rr8 + t0_r6_c8_rr9;

  assign t2_r6_c8_rr0 = t1_r6_c8_rr0 + t1_r6_c8_rr1;
  assign t2_r6_c8_rr1 = t1_r6_c8_rr2 + t1_r6_c8_rr3;
  assign t2_r6_c8_rr2 = t1_r6_c8_rr4;

  assign t3_r6_c8_rr0 = t2_r6_c8_rr0 + t2_r6_c8_rr1;
  assign t3_r6_c8_rr1 = t2_r6_c8_rr2;

  assign t4_r6_c8_rr0 = t3_r6_c8_rr0 + t3_r6_c8_rr1;

  assign c_6_8 = t4_r6_c8_rr0;
  assign t0_r6_c9_rr0 = a_6_0 * b_0_9;
  assign t0_r6_c9_rr1 = a_6_1 * b_1_9;
  assign t0_r6_c9_rr2 = a_6_2 * b_2_9;
  assign t0_r6_c9_rr3 = a_6_3 * b_3_9;
  assign t0_r6_c9_rr4 = a_6_4 * b_4_9;
  assign t0_r6_c9_rr5 = a_6_5 * b_5_9;
  assign t0_r6_c9_rr6 = a_6_6 * b_6_9;
  assign t0_r6_c9_rr7 = a_6_7 * b_7_9;
  assign t0_r6_c9_rr8 = a_6_8 * b_8_9;
  assign t0_r6_c9_rr9 = a_6_9 * b_9_9;
  assign t1_r6_c9_rr0 = t0_r6_c9_rr0 + t0_r6_c9_rr1;
  assign t1_r6_c9_rr1 = t0_r6_c9_rr2 + t0_r6_c9_rr3;
  assign t1_r6_c9_rr2 = t0_r6_c9_rr4 + t0_r6_c9_rr5;
  assign t1_r6_c9_rr3 = t0_r6_c9_rr6 + t0_r6_c9_rr7;
  assign t1_r6_c9_rr4 = t0_r6_c9_rr8 + t0_r6_c9_rr9;

  assign t2_r6_c9_rr0 = t1_r6_c9_rr0 + t1_r6_c9_rr1;
  assign t2_r6_c9_rr1 = t1_r6_c9_rr2 + t1_r6_c9_rr3;
  assign t2_r6_c9_rr2 = t1_r6_c9_rr4;

  assign t3_r6_c9_rr0 = t2_r6_c9_rr0 + t2_r6_c9_rr1;
  assign t3_r6_c9_rr1 = t2_r6_c9_rr2;

  assign t4_r6_c9_rr0 = t3_r6_c9_rr0 + t3_r6_c9_rr1;

  assign c_6_9 = t4_r6_c9_rr0;
  assign t0_r7_c0_rr0 = a_7_0 * b_0_0;
  assign t0_r7_c0_rr1 = a_7_1 * b_1_0;
  assign t0_r7_c0_rr2 = a_7_2 * b_2_0;
  assign t0_r7_c0_rr3 = a_7_3 * b_3_0;
  assign t0_r7_c0_rr4 = a_7_4 * b_4_0;
  assign t0_r7_c0_rr5 = a_7_5 * b_5_0;
  assign t0_r7_c0_rr6 = a_7_6 * b_6_0;
  assign t0_r7_c0_rr7 = a_7_7 * b_7_0;
  assign t0_r7_c0_rr8 = a_7_8 * b_8_0;
  assign t0_r7_c0_rr9 = a_7_9 * b_9_0;
  assign t1_r7_c0_rr0 = t0_r7_c0_rr0 + t0_r7_c0_rr1;
  assign t1_r7_c0_rr1 = t0_r7_c0_rr2 + t0_r7_c0_rr3;
  assign t1_r7_c0_rr2 = t0_r7_c0_rr4 + t0_r7_c0_rr5;
  assign t1_r7_c0_rr3 = t0_r7_c0_rr6 + t0_r7_c0_rr7;
  assign t1_r7_c0_rr4 = t0_r7_c0_rr8 + t0_r7_c0_rr9;

  assign t2_r7_c0_rr0 = t1_r7_c0_rr0 + t1_r7_c0_rr1;
  assign t2_r7_c0_rr1 = t1_r7_c0_rr2 + t1_r7_c0_rr3;
  assign t2_r7_c0_rr2 = t1_r7_c0_rr4;

  assign t3_r7_c0_rr0 = t2_r7_c0_rr0 + t2_r7_c0_rr1;
  assign t3_r7_c0_rr1 = t2_r7_c0_rr2;

  assign t4_r7_c0_rr0 = t3_r7_c0_rr0 + t3_r7_c0_rr1;

  assign c_7_0 = t4_r7_c0_rr0;
  assign t0_r7_c1_rr0 = a_7_0 * b_0_1;
  assign t0_r7_c1_rr1 = a_7_1 * b_1_1;
  assign t0_r7_c1_rr2 = a_7_2 * b_2_1;
  assign t0_r7_c1_rr3 = a_7_3 * b_3_1;
  assign t0_r7_c1_rr4 = a_7_4 * b_4_1;
  assign t0_r7_c1_rr5 = a_7_5 * b_5_1;
  assign t0_r7_c1_rr6 = a_7_6 * b_6_1;
  assign t0_r7_c1_rr7 = a_7_7 * b_7_1;
  assign t0_r7_c1_rr8 = a_7_8 * b_8_1;
  assign t0_r7_c1_rr9 = a_7_9 * b_9_1;
  assign t1_r7_c1_rr0 = t0_r7_c1_rr0 + t0_r7_c1_rr1;
  assign t1_r7_c1_rr1 = t0_r7_c1_rr2 + t0_r7_c1_rr3;
  assign t1_r7_c1_rr2 = t0_r7_c1_rr4 + t0_r7_c1_rr5;
  assign t1_r7_c1_rr3 = t0_r7_c1_rr6 + t0_r7_c1_rr7;
  assign t1_r7_c1_rr4 = t0_r7_c1_rr8 + t0_r7_c1_rr9;

  assign t2_r7_c1_rr0 = t1_r7_c1_rr0 + t1_r7_c1_rr1;
  assign t2_r7_c1_rr1 = t1_r7_c1_rr2 + t1_r7_c1_rr3;
  assign t2_r7_c1_rr2 = t1_r7_c1_rr4;

  assign t3_r7_c1_rr0 = t2_r7_c1_rr0 + t2_r7_c1_rr1;
  assign t3_r7_c1_rr1 = t2_r7_c1_rr2;

  assign t4_r7_c1_rr0 = t3_r7_c1_rr0 + t3_r7_c1_rr1;

  assign c_7_1 = t4_r7_c1_rr0;
  assign t0_r7_c2_rr0 = a_7_0 * b_0_2;
  assign t0_r7_c2_rr1 = a_7_1 * b_1_2;
  assign t0_r7_c2_rr2 = a_7_2 * b_2_2;
  assign t0_r7_c2_rr3 = a_7_3 * b_3_2;
  assign t0_r7_c2_rr4 = a_7_4 * b_4_2;
  assign t0_r7_c2_rr5 = a_7_5 * b_5_2;
  assign t0_r7_c2_rr6 = a_7_6 * b_6_2;
  assign t0_r7_c2_rr7 = a_7_7 * b_7_2;
  assign t0_r7_c2_rr8 = a_7_8 * b_8_2;
  assign t0_r7_c2_rr9 = a_7_9 * b_9_2;
  assign t1_r7_c2_rr0 = t0_r7_c2_rr0 + t0_r7_c2_rr1;
  assign t1_r7_c2_rr1 = t0_r7_c2_rr2 + t0_r7_c2_rr3;
  assign t1_r7_c2_rr2 = t0_r7_c2_rr4 + t0_r7_c2_rr5;
  assign t1_r7_c2_rr3 = t0_r7_c2_rr6 + t0_r7_c2_rr7;
  assign t1_r7_c2_rr4 = t0_r7_c2_rr8 + t0_r7_c2_rr9;

  assign t2_r7_c2_rr0 = t1_r7_c2_rr0 + t1_r7_c2_rr1;
  assign t2_r7_c2_rr1 = t1_r7_c2_rr2 + t1_r7_c2_rr3;
  assign t2_r7_c2_rr2 = t1_r7_c2_rr4;

  assign t3_r7_c2_rr0 = t2_r7_c2_rr0 + t2_r7_c2_rr1;
  assign t3_r7_c2_rr1 = t2_r7_c2_rr2;

  assign t4_r7_c2_rr0 = t3_r7_c2_rr0 + t3_r7_c2_rr1;

  assign c_7_2 = t4_r7_c2_rr0;
  assign t0_r7_c3_rr0 = a_7_0 * b_0_3;
  assign t0_r7_c3_rr1 = a_7_1 * b_1_3;
  assign t0_r7_c3_rr2 = a_7_2 * b_2_3;
  assign t0_r7_c3_rr3 = a_7_3 * b_3_3;
  assign t0_r7_c3_rr4 = a_7_4 * b_4_3;
  assign t0_r7_c3_rr5 = a_7_5 * b_5_3;
  assign t0_r7_c3_rr6 = a_7_6 * b_6_3;
  assign t0_r7_c3_rr7 = a_7_7 * b_7_3;
  assign t0_r7_c3_rr8 = a_7_8 * b_8_3;
  assign t0_r7_c3_rr9 = a_7_9 * b_9_3;
  assign t1_r7_c3_rr0 = t0_r7_c3_rr0 + t0_r7_c3_rr1;
  assign t1_r7_c3_rr1 = t0_r7_c3_rr2 + t0_r7_c3_rr3;
  assign t1_r7_c3_rr2 = t0_r7_c3_rr4 + t0_r7_c3_rr5;
  assign t1_r7_c3_rr3 = t0_r7_c3_rr6 + t0_r7_c3_rr7;
  assign t1_r7_c3_rr4 = t0_r7_c3_rr8 + t0_r7_c3_rr9;

  assign t2_r7_c3_rr0 = t1_r7_c3_rr0 + t1_r7_c3_rr1;
  assign t2_r7_c3_rr1 = t1_r7_c3_rr2 + t1_r7_c3_rr3;
  assign t2_r7_c3_rr2 = t1_r7_c3_rr4;

  assign t3_r7_c3_rr0 = t2_r7_c3_rr0 + t2_r7_c3_rr1;
  assign t3_r7_c3_rr1 = t2_r7_c3_rr2;

  assign t4_r7_c3_rr0 = t3_r7_c3_rr0 + t3_r7_c3_rr1;

  assign c_7_3 = t4_r7_c3_rr0;
  assign t0_r7_c4_rr0 = a_7_0 * b_0_4;
  assign t0_r7_c4_rr1 = a_7_1 * b_1_4;
  assign t0_r7_c4_rr2 = a_7_2 * b_2_4;
  assign t0_r7_c4_rr3 = a_7_3 * b_3_4;
  assign t0_r7_c4_rr4 = a_7_4 * b_4_4;
  assign t0_r7_c4_rr5 = a_7_5 * b_5_4;
  assign t0_r7_c4_rr6 = a_7_6 * b_6_4;
  assign t0_r7_c4_rr7 = a_7_7 * b_7_4;
  assign t0_r7_c4_rr8 = a_7_8 * b_8_4;
  assign t0_r7_c4_rr9 = a_7_9 * b_9_4;
  assign t1_r7_c4_rr0 = t0_r7_c4_rr0 + t0_r7_c4_rr1;
  assign t1_r7_c4_rr1 = t0_r7_c4_rr2 + t0_r7_c4_rr3;
  assign t1_r7_c4_rr2 = t0_r7_c4_rr4 + t0_r7_c4_rr5;
  assign t1_r7_c4_rr3 = t0_r7_c4_rr6 + t0_r7_c4_rr7;
  assign t1_r7_c4_rr4 = t0_r7_c4_rr8 + t0_r7_c4_rr9;

  assign t2_r7_c4_rr0 = t1_r7_c4_rr0 + t1_r7_c4_rr1;
  assign t2_r7_c4_rr1 = t1_r7_c4_rr2 + t1_r7_c4_rr3;
  assign t2_r7_c4_rr2 = t1_r7_c4_rr4;

  assign t3_r7_c4_rr0 = t2_r7_c4_rr0 + t2_r7_c4_rr1;
  assign t3_r7_c4_rr1 = t2_r7_c4_rr2;

  assign t4_r7_c4_rr0 = t3_r7_c4_rr0 + t3_r7_c4_rr1;

  assign c_7_4 = t4_r7_c4_rr0;
  assign t0_r7_c5_rr0 = a_7_0 * b_0_5;
  assign t0_r7_c5_rr1 = a_7_1 * b_1_5;
  assign t0_r7_c5_rr2 = a_7_2 * b_2_5;
  assign t0_r7_c5_rr3 = a_7_3 * b_3_5;
  assign t0_r7_c5_rr4 = a_7_4 * b_4_5;
  assign t0_r7_c5_rr5 = a_7_5 * b_5_5;
  assign t0_r7_c5_rr6 = a_7_6 * b_6_5;
  assign t0_r7_c5_rr7 = a_7_7 * b_7_5;
  assign t0_r7_c5_rr8 = a_7_8 * b_8_5;
  assign t0_r7_c5_rr9 = a_7_9 * b_9_5;
  assign t1_r7_c5_rr0 = t0_r7_c5_rr0 + t0_r7_c5_rr1;
  assign t1_r7_c5_rr1 = t0_r7_c5_rr2 + t0_r7_c5_rr3;
  assign t1_r7_c5_rr2 = t0_r7_c5_rr4 + t0_r7_c5_rr5;
  assign t1_r7_c5_rr3 = t0_r7_c5_rr6 + t0_r7_c5_rr7;
  assign t1_r7_c5_rr4 = t0_r7_c5_rr8 + t0_r7_c5_rr9;

  assign t2_r7_c5_rr0 = t1_r7_c5_rr0 + t1_r7_c5_rr1;
  assign t2_r7_c5_rr1 = t1_r7_c5_rr2 + t1_r7_c5_rr3;
  assign t2_r7_c5_rr2 = t1_r7_c5_rr4;

  assign t3_r7_c5_rr0 = t2_r7_c5_rr0 + t2_r7_c5_rr1;
  assign t3_r7_c5_rr1 = t2_r7_c5_rr2;

  assign t4_r7_c5_rr0 = t3_r7_c5_rr0 + t3_r7_c5_rr1;

  assign c_7_5 = t4_r7_c5_rr0;
  assign t0_r7_c6_rr0 = a_7_0 * b_0_6;
  assign t0_r7_c6_rr1 = a_7_1 * b_1_6;
  assign t0_r7_c6_rr2 = a_7_2 * b_2_6;
  assign t0_r7_c6_rr3 = a_7_3 * b_3_6;
  assign t0_r7_c6_rr4 = a_7_4 * b_4_6;
  assign t0_r7_c6_rr5 = a_7_5 * b_5_6;
  assign t0_r7_c6_rr6 = a_7_6 * b_6_6;
  assign t0_r7_c6_rr7 = a_7_7 * b_7_6;
  assign t0_r7_c6_rr8 = a_7_8 * b_8_6;
  assign t0_r7_c6_rr9 = a_7_9 * b_9_6;
  assign t1_r7_c6_rr0 = t0_r7_c6_rr0 + t0_r7_c6_rr1;
  assign t1_r7_c6_rr1 = t0_r7_c6_rr2 + t0_r7_c6_rr3;
  assign t1_r7_c6_rr2 = t0_r7_c6_rr4 + t0_r7_c6_rr5;
  assign t1_r7_c6_rr3 = t0_r7_c6_rr6 + t0_r7_c6_rr7;
  assign t1_r7_c6_rr4 = t0_r7_c6_rr8 + t0_r7_c6_rr9;

  assign t2_r7_c6_rr0 = t1_r7_c6_rr0 + t1_r7_c6_rr1;
  assign t2_r7_c6_rr1 = t1_r7_c6_rr2 + t1_r7_c6_rr3;
  assign t2_r7_c6_rr2 = t1_r7_c6_rr4;

  assign t3_r7_c6_rr0 = t2_r7_c6_rr0 + t2_r7_c6_rr1;
  assign t3_r7_c6_rr1 = t2_r7_c6_rr2;

  assign t4_r7_c6_rr0 = t3_r7_c6_rr0 + t3_r7_c6_rr1;

  assign c_7_6 = t4_r7_c6_rr0;
  assign t0_r7_c7_rr0 = a_7_0 * b_0_7;
  assign t0_r7_c7_rr1 = a_7_1 * b_1_7;
  assign t0_r7_c7_rr2 = a_7_2 * b_2_7;
  assign t0_r7_c7_rr3 = a_7_3 * b_3_7;
  assign t0_r7_c7_rr4 = a_7_4 * b_4_7;
  assign t0_r7_c7_rr5 = a_7_5 * b_5_7;
  assign t0_r7_c7_rr6 = a_7_6 * b_6_7;
  assign t0_r7_c7_rr7 = a_7_7 * b_7_7;
  assign t0_r7_c7_rr8 = a_7_8 * b_8_7;
  assign t0_r7_c7_rr9 = a_7_9 * b_9_7;
  assign t1_r7_c7_rr0 = t0_r7_c7_rr0 + t0_r7_c7_rr1;
  assign t1_r7_c7_rr1 = t0_r7_c7_rr2 + t0_r7_c7_rr3;
  assign t1_r7_c7_rr2 = t0_r7_c7_rr4 + t0_r7_c7_rr5;
  assign t1_r7_c7_rr3 = t0_r7_c7_rr6 + t0_r7_c7_rr7;
  assign t1_r7_c7_rr4 = t0_r7_c7_rr8 + t0_r7_c7_rr9;

  assign t2_r7_c7_rr0 = t1_r7_c7_rr0 + t1_r7_c7_rr1;
  assign t2_r7_c7_rr1 = t1_r7_c7_rr2 + t1_r7_c7_rr3;
  assign t2_r7_c7_rr2 = t1_r7_c7_rr4;

  assign t3_r7_c7_rr0 = t2_r7_c7_rr0 + t2_r7_c7_rr1;
  assign t3_r7_c7_rr1 = t2_r7_c7_rr2;

  assign t4_r7_c7_rr0 = t3_r7_c7_rr0 + t3_r7_c7_rr1;

  assign c_7_7 = t4_r7_c7_rr0;
  assign t0_r7_c8_rr0 = a_7_0 * b_0_8;
  assign t0_r7_c8_rr1 = a_7_1 * b_1_8;
  assign t0_r7_c8_rr2 = a_7_2 * b_2_8;
  assign t0_r7_c8_rr3 = a_7_3 * b_3_8;
  assign t0_r7_c8_rr4 = a_7_4 * b_4_8;
  assign t0_r7_c8_rr5 = a_7_5 * b_5_8;
  assign t0_r7_c8_rr6 = a_7_6 * b_6_8;
  assign t0_r7_c8_rr7 = a_7_7 * b_7_8;
  assign t0_r7_c8_rr8 = a_7_8 * b_8_8;
  assign t0_r7_c8_rr9 = a_7_9 * b_9_8;
  assign t1_r7_c8_rr0 = t0_r7_c8_rr0 + t0_r7_c8_rr1;
  assign t1_r7_c8_rr1 = t0_r7_c8_rr2 + t0_r7_c8_rr3;
  assign t1_r7_c8_rr2 = t0_r7_c8_rr4 + t0_r7_c8_rr5;
  assign t1_r7_c8_rr3 = t0_r7_c8_rr6 + t0_r7_c8_rr7;
  assign t1_r7_c8_rr4 = t0_r7_c8_rr8 + t0_r7_c8_rr9;

  assign t2_r7_c8_rr0 = t1_r7_c8_rr0 + t1_r7_c8_rr1;
  assign t2_r7_c8_rr1 = t1_r7_c8_rr2 + t1_r7_c8_rr3;
  assign t2_r7_c8_rr2 = t1_r7_c8_rr4;

  assign t3_r7_c8_rr0 = t2_r7_c8_rr0 + t2_r7_c8_rr1;
  assign t3_r7_c8_rr1 = t2_r7_c8_rr2;

  assign t4_r7_c8_rr0 = t3_r7_c8_rr0 + t3_r7_c8_rr1;

  assign c_7_8 = t4_r7_c8_rr0;
  assign t0_r7_c9_rr0 = a_7_0 * b_0_9;
  assign t0_r7_c9_rr1 = a_7_1 * b_1_9;
  assign t0_r7_c9_rr2 = a_7_2 * b_2_9;
  assign t0_r7_c9_rr3 = a_7_3 * b_3_9;
  assign t0_r7_c9_rr4 = a_7_4 * b_4_9;
  assign t0_r7_c9_rr5 = a_7_5 * b_5_9;
  assign t0_r7_c9_rr6 = a_7_6 * b_6_9;
  assign t0_r7_c9_rr7 = a_7_7 * b_7_9;
  assign t0_r7_c9_rr8 = a_7_8 * b_8_9;
  assign t0_r7_c9_rr9 = a_7_9 * b_9_9;
  assign t1_r7_c9_rr0 = t0_r7_c9_rr0 + t0_r7_c9_rr1;
  assign t1_r7_c9_rr1 = t0_r7_c9_rr2 + t0_r7_c9_rr3;
  assign t1_r7_c9_rr2 = t0_r7_c9_rr4 + t0_r7_c9_rr5;
  assign t1_r7_c9_rr3 = t0_r7_c9_rr6 + t0_r7_c9_rr7;
  assign t1_r7_c9_rr4 = t0_r7_c9_rr8 + t0_r7_c9_rr9;

  assign t2_r7_c9_rr0 = t1_r7_c9_rr0 + t1_r7_c9_rr1;
  assign t2_r7_c9_rr1 = t1_r7_c9_rr2 + t1_r7_c9_rr3;
  assign t2_r7_c9_rr2 = t1_r7_c9_rr4;

  assign t3_r7_c9_rr0 = t2_r7_c9_rr0 + t2_r7_c9_rr1;
  assign t3_r7_c9_rr1 = t2_r7_c9_rr2;

  assign t4_r7_c9_rr0 = t3_r7_c9_rr0 + t3_r7_c9_rr1;

  assign c_7_9 = t4_r7_c9_rr0;
  assign t0_r8_c0_rr0 = a_8_0 * b_0_0;
  assign t0_r8_c0_rr1 = a_8_1 * b_1_0;
  assign t0_r8_c0_rr2 = a_8_2 * b_2_0;
  assign t0_r8_c0_rr3 = a_8_3 * b_3_0;
  assign t0_r8_c0_rr4 = a_8_4 * b_4_0;
  assign t0_r8_c0_rr5 = a_8_5 * b_5_0;
  assign t0_r8_c0_rr6 = a_8_6 * b_6_0;
  assign t0_r8_c0_rr7 = a_8_7 * b_7_0;
  assign t0_r8_c0_rr8 = a_8_8 * b_8_0;
  assign t0_r8_c0_rr9 = a_8_9 * b_9_0;
  assign t1_r8_c0_rr0 = t0_r8_c0_rr0 + t0_r8_c0_rr1;
  assign t1_r8_c0_rr1 = t0_r8_c0_rr2 + t0_r8_c0_rr3;
  assign t1_r8_c0_rr2 = t0_r8_c0_rr4 + t0_r8_c0_rr5;
  assign t1_r8_c0_rr3 = t0_r8_c0_rr6 + t0_r8_c0_rr7;
  assign t1_r8_c0_rr4 = t0_r8_c0_rr8 + t0_r8_c0_rr9;

  assign t2_r8_c0_rr0 = t1_r8_c0_rr0 + t1_r8_c0_rr1;
  assign t2_r8_c0_rr1 = t1_r8_c0_rr2 + t1_r8_c0_rr3;
  assign t2_r8_c0_rr2 = t1_r8_c0_rr4;

  assign t3_r8_c0_rr0 = t2_r8_c0_rr0 + t2_r8_c0_rr1;
  assign t3_r8_c0_rr1 = t2_r8_c0_rr2;

  assign t4_r8_c0_rr0 = t3_r8_c0_rr0 + t3_r8_c0_rr1;

  assign c_8_0 = t4_r8_c0_rr0;
  assign t0_r8_c1_rr0 = a_8_0 * b_0_1;
  assign t0_r8_c1_rr1 = a_8_1 * b_1_1;
  assign t0_r8_c1_rr2 = a_8_2 * b_2_1;
  assign t0_r8_c1_rr3 = a_8_3 * b_3_1;
  assign t0_r8_c1_rr4 = a_8_4 * b_4_1;
  assign t0_r8_c1_rr5 = a_8_5 * b_5_1;
  assign t0_r8_c1_rr6 = a_8_6 * b_6_1;
  assign t0_r8_c1_rr7 = a_8_7 * b_7_1;
  assign t0_r8_c1_rr8 = a_8_8 * b_8_1;
  assign t0_r8_c1_rr9 = a_8_9 * b_9_1;
  assign t1_r8_c1_rr0 = t0_r8_c1_rr0 + t0_r8_c1_rr1;
  assign t1_r8_c1_rr1 = t0_r8_c1_rr2 + t0_r8_c1_rr3;
  assign t1_r8_c1_rr2 = t0_r8_c1_rr4 + t0_r8_c1_rr5;
  assign t1_r8_c1_rr3 = t0_r8_c1_rr6 + t0_r8_c1_rr7;
  assign t1_r8_c1_rr4 = t0_r8_c1_rr8 + t0_r8_c1_rr9;

  assign t2_r8_c1_rr0 = t1_r8_c1_rr0 + t1_r8_c1_rr1;
  assign t2_r8_c1_rr1 = t1_r8_c1_rr2 + t1_r8_c1_rr3;
  assign t2_r8_c1_rr2 = t1_r8_c1_rr4;

  assign t3_r8_c1_rr0 = t2_r8_c1_rr0 + t2_r8_c1_rr1;
  assign t3_r8_c1_rr1 = t2_r8_c1_rr2;

  assign t4_r8_c1_rr0 = t3_r8_c1_rr0 + t3_r8_c1_rr1;

  assign c_8_1 = t4_r8_c1_rr0;
  assign t0_r8_c2_rr0 = a_8_0 * b_0_2;
  assign t0_r8_c2_rr1 = a_8_1 * b_1_2;
  assign t0_r8_c2_rr2 = a_8_2 * b_2_2;
  assign t0_r8_c2_rr3 = a_8_3 * b_3_2;
  assign t0_r8_c2_rr4 = a_8_4 * b_4_2;
  assign t0_r8_c2_rr5 = a_8_5 * b_5_2;
  assign t0_r8_c2_rr6 = a_8_6 * b_6_2;
  assign t0_r8_c2_rr7 = a_8_7 * b_7_2;
  assign t0_r8_c2_rr8 = a_8_8 * b_8_2;
  assign t0_r8_c2_rr9 = a_8_9 * b_9_2;
  assign t1_r8_c2_rr0 = t0_r8_c2_rr0 + t0_r8_c2_rr1;
  assign t1_r8_c2_rr1 = t0_r8_c2_rr2 + t0_r8_c2_rr3;
  assign t1_r8_c2_rr2 = t0_r8_c2_rr4 + t0_r8_c2_rr5;
  assign t1_r8_c2_rr3 = t0_r8_c2_rr6 + t0_r8_c2_rr7;
  assign t1_r8_c2_rr4 = t0_r8_c2_rr8 + t0_r8_c2_rr9;

  assign t2_r8_c2_rr0 = t1_r8_c2_rr0 + t1_r8_c2_rr1;
  assign t2_r8_c2_rr1 = t1_r8_c2_rr2 + t1_r8_c2_rr3;
  assign t2_r8_c2_rr2 = t1_r8_c2_rr4;

  assign t3_r8_c2_rr0 = t2_r8_c2_rr0 + t2_r8_c2_rr1;
  assign t3_r8_c2_rr1 = t2_r8_c2_rr2;

  assign t4_r8_c2_rr0 = t3_r8_c2_rr0 + t3_r8_c2_rr1;

  assign c_8_2 = t4_r8_c2_rr0;
  assign t0_r8_c3_rr0 = a_8_0 * b_0_3;
  assign t0_r8_c3_rr1 = a_8_1 * b_1_3;
  assign t0_r8_c3_rr2 = a_8_2 * b_2_3;
  assign t0_r8_c3_rr3 = a_8_3 * b_3_3;
  assign t0_r8_c3_rr4 = a_8_4 * b_4_3;
  assign t0_r8_c3_rr5 = a_8_5 * b_5_3;
  assign t0_r8_c3_rr6 = a_8_6 * b_6_3;
  assign t0_r8_c3_rr7 = a_8_7 * b_7_3;
  assign t0_r8_c3_rr8 = a_8_8 * b_8_3;
  assign t0_r8_c3_rr9 = a_8_9 * b_9_3;
  assign t1_r8_c3_rr0 = t0_r8_c3_rr0 + t0_r8_c3_rr1;
  assign t1_r8_c3_rr1 = t0_r8_c3_rr2 + t0_r8_c3_rr3;
  assign t1_r8_c3_rr2 = t0_r8_c3_rr4 + t0_r8_c3_rr5;
  assign t1_r8_c3_rr3 = t0_r8_c3_rr6 + t0_r8_c3_rr7;
  assign t1_r8_c3_rr4 = t0_r8_c3_rr8 + t0_r8_c3_rr9;

  assign t2_r8_c3_rr0 = t1_r8_c3_rr0 + t1_r8_c3_rr1;
  assign t2_r8_c3_rr1 = t1_r8_c3_rr2 + t1_r8_c3_rr3;
  assign t2_r8_c3_rr2 = t1_r8_c3_rr4;

  assign t3_r8_c3_rr0 = t2_r8_c3_rr0 + t2_r8_c3_rr1;
  assign t3_r8_c3_rr1 = t2_r8_c3_rr2;

  assign t4_r8_c3_rr0 = t3_r8_c3_rr0 + t3_r8_c3_rr1;

  assign c_8_3 = t4_r8_c3_rr0;
  assign t0_r8_c4_rr0 = a_8_0 * b_0_4;
  assign t0_r8_c4_rr1 = a_8_1 * b_1_4;
  assign t0_r8_c4_rr2 = a_8_2 * b_2_4;
  assign t0_r8_c4_rr3 = a_8_3 * b_3_4;
  assign t0_r8_c4_rr4 = a_8_4 * b_4_4;
  assign t0_r8_c4_rr5 = a_8_5 * b_5_4;
  assign t0_r8_c4_rr6 = a_8_6 * b_6_4;
  assign t0_r8_c4_rr7 = a_8_7 * b_7_4;
  assign t0_r8_c4_rr8 = a_8_8 * b_8_4;
  assign t0_r8_c4_rr9 = a_8_9 * b_9_4;
  assign t1_r8_c4_rr0 = t0_r8_c4_rr0 + t0_r8_c4_rr1;
  assign t1_r8_c4_rr1 = t0_r8_c4_rr2 + t0_r8_c4_rr3;
  assign t1_r8_c4_rr2 = t0_r8_c4_rr4 + t0_r8_c4_rr5;
  assign t1_r8_c4_rr3 = t0_r8_c4_rr6 + t0_r8_c4_rr7;
  assign t1_r8_c4_rr4 = t0_r8_c4_rr8 + t0_r8_c4_rr9;

  assign t2_r8_c4_rr0 = t1_r8_c4_rr0 + t1_r8_c4_rr1;
  assign t2_r8_c4_rr1 = t1_r8_c4_rr2 + t1_r8_c4_rr3;
  assign t2_r8_c4_rr2 = t1_r8_c4_rr4;

  assign t3_r8_c4_rr0 = t2_r8_c4_rr0 + t2_r8_c4_rr1;
  assign t3_r8_c4_rr1 = t2_r8_c4_rr2;

  assign t4_r8_c4_rr0 = t3_r8_c4_rr0 + t3_r8_c4_rr1;

  assign c_8_4 = t4_r8_c4_rr0;
  assign t0_r8_c5_rr0 = a_8_0 * b_0_5;
  assign t0_r8_c5_rr1 = a_8_1 * b_1_5;
  assign t0_r8_c5_rr2 = a_8_2 * b_2_5;
  assign t0_r8_c5_rr3 = a_8_3 * b_3_5;
  assign t0_r8_c5_rr4 = a_8_4 * b_4_5;
  assign t0_r8_c5_rr5 = a_8_5 * b_5_5;
  assign t0_r8_c5_rr6 = a_8_6 * b_6_5;
  assign t0_r8_c5_rr7 = a_8_7 * b_7_5;
  assign t0_r8_c5_rr8 = a_8_8 * b_8_5;
  assign t0_r8_c5_rr9 = a_8_9 * b_9_5;
  assign t1_r8_c5_rr0 = t0_r8_c5_rr0 + t0_r8_c5_rr1;
  assign t1_r8_c5_rr1 = t0_r8_c5_rr2 + t0_r8_c5_rr3;
  assign t1_r8_c5_rr2 = t0_r8_c5_rr4 + t0_r8_c5_rr5;
  assign t1_r8_c5_rr3 = t0_r8_c5_rr6 + t0_r8_c5_rr7;
  assign t1_r8_c5_rr4 = t0_r8_c5_rr8 + t0_r8_c5_rr9;

  assign t2_r8_c5_rr0 = t1_r8_c5_rr0 + t1_r8_c5_rr1;
  assign t2_r8_c5_rr1 = t1_r8_c5_rr2 + t1_r8_c5_rr3;
  assign t2_r8_c5_rr2 = t1_r8_c5_rr4;

  assign t3_r8_c5_rr0 = t2_r8_c5_rr0 + t2_r8_c5_rr1;
  assign t3_r8_c5_rr1 = t2_r8_c5_rr2;

  assign t4_r8_c5_rr0 = t3_r8_c5_rr0 + t3_r8_c5_rr1;

  assign c_8_5 = t4_r8_c5_rr0;
  assign t0_r8_c6_rr0 = a_8_0 * b_0_6;
  assign t0_r8_c6_rr1 = a_8_1 * b_1_6;
  assign t0_r8_c6_rr2 = a_8_2 * b_2_6;
  assign t0_r8_c6_rr3 = a_8_3 * b_3_6;
  assign t0_r8_c6_rr4 = a_8_4 * b_4_6;
  assign t0_r8_c6_rr5 = a_8_5 * b_5_6;
  assign t0_r8_c6_rr6 = a_8_6 * b_6_6;
  assign t0_r8_c6_rr7 = a_8_7 * b_7_6;
  assign t0_r8_c6_rr8 = a_8_8 * b_8_6;
  assign t0_r8_c6_rr9 = a_8_9 * b_9_6;
  assign t1_r8_c6_rr0 = t0_r8_c6_rr0 + t0_r8_c6_rr1;
  assign t1_r8_c6_rr1 = t0_r8_c6_rr2 + t0_r8_c6_rr3;
  assign t1_r8_c6_rr2 = t0_r8_c6_rr4 + t0_r8_c6_rr5;
  assign t1_r8_c6_rr3 = t0_r8_c6_rr6 + t0_r8_c6_rr7;
  assign t1_r8_c6_rr4 = t0_r8_c6_rr8 + t0_r8_c6_rr9;

  assign t2_r8_c6_rr0 = t1_r8_c6_rr0 + t1_r8_c6_rr1;
  assign t2_r8_c6_rr1 = t1_r8_c6_rr2 + t1_r8_c6_rr3;
  assign t2_r8_c6_rr2 = t1_r8_c6_rr4;

  assign t3_r8_c6_rr0 = t2_r8_c6_rr0 + t2_r8_c6_rr1;
  assign t3_r8_c6_rr1 = t2_r8_c6_rr2;

  assign t4_r8_c6_rr0 = t3_r8_c6_rr0 + t3_r8_c6_rr1;

  assign c_8_6 = t4_r8_c6_rr0;
  assign t0_r8_c7_rr0 = a_8_0 * b_0_7;
  assign t0_r8_c7_rr1 = a_8_1 * b_1_7;
  assign t0_r8_c7_rr2 = a_8_2 * b_2_7;
  assign t0_r8_c7_rr3 = a_8_3 * b_3_7;
  assign t0_r8_c7_rr4 = a_8_4 * b_4_7;
  assign t0_r8_c7_rr5 = a_8_5 * b_5_7;
  assign t0_r8_c7_rr6 = a_8_6 * b_6_7;
  assign t0_r8_c7_rr7 = a_8_7 * b_7_7;
  assign t0_r8_c7_rr8 = a_8_8 * b_8_7;
  assign t0_r8_c7_rr9 = a_8_9 * b_9_7;
  assign t1_r8_c7_rr0 = t0_r8_c7_rr0 + t0_r8_c7_rr1;
  assign t1_r8_c7_rr1 = t0_r8_c7_rr2 + t0_r8_c7_rr3;
  assign t1_r8_c7_rr2 = t0_r8_c7_rr4 + t0_r8_c7_rr5;
  assign t1_r8_c7_rr3 = t0_r8_c7_rr6 + t0_r8_c7_rr7;
  assign t1_r8_c7_rr4 = t0_r8_c7_rr8 + t0_r8_c7_rr9;

  assign t2_r8_c7_rr0 = t1_r8_c7_rr0 + t1_r8_c7_rr1;
  assign t2_r8_c7_rr1 = t1_r8_c7_rr2 + t1_r8_c7_rr3;
  assign t2_r8_c7_rr2 = t1_r8_c7_rr4;

  assign t3_r8_c7_rr0 = t2_r8_c7_rr0 + t2_r8_c7_rr1;
  assign t3_r8_c7_rr1 = t2_r8_c7_rr2;

  assign t4_r8_c7_rr0 = t3_r8_c7_rr0 + t3_r8_c7_rr1;

  assign c_8_7 = t4_r8_c7_rr0;
  assign t0_r8_c8_rr0 = a_8_0 * b_0_8;
  assign t0_r8_c8_rr1 = a_8_1 * b_1_8;
  assign t0_r8_c8_rr2 = a_8_2 * b_2_8;
  assign t0_r8_c8_rr3 = a_8_3 * b_3_8;
  assign t0_r8_c8_rr4 = a_8_4 * b_4_8;
  assign t0_r8_c8_rr5 = a_8_5 * b_5_8;
  assign t0_r8_c8_rr6 = a_8_6 * b_6_8;
  assign t0_r8_c8_rr7 = a_8_7 * b_7_8;
  assign t0_r8_c8_rr8 = a_8_8 * b_8_8;
  assign t0_r8_c8_rr9 = a_8_9 * b_9_8;
  assign t1_r8_c8_rr0 = t0_r8_c8_rr0 + t0_r8_c8_rr1;
  assign t1_r8_c8_rr1 = t0_r8_c8_rr2 + t0_r8_c8_rr3;
  assign t1_r8_c8_rr2 = t0_r8_c8_rr4 + t0_r8_c8_rr5;
  assign t1_r8_c8_rr3 = t0_r8_c8_rr6 + t0_r8_c8_rr7;
  assign t1_r8_c8_rr4 = t0_r8_c8_rr8 + t0_r8_c8_rr9;

  assign t2_r8_c8_rr0 = t1_r8_c8_rr0 + t1_r8_c8_rr1;
  assign t2_r8_c8_rr1 = t1_r8_c8_rr2 + t1_r8_c8_rr3;
  assign t2_r8_c8_rr2 = t1_r8_c8_rr4;

  assign t3_r8_c8_rr0 = t2_r8_c8_rr0 + t2_r8_c8_rr1;
  assign t3_r8_c8_rr1 = t2_r8_c8_rr2;

  assign t4_r8_c8_rr0 = t3_r8_c8_rr0 + t3_r8_c8_rr1;

  assign c_8_8 = t4_r8_c8_rr0;
  assign t0_r8_c9_rr0 = a_8_0 * b_0_9;
  assign t0_r8_c9_rr1 = a_8_1 * b_1_9;
  assign t0_r8_c9_rr2 = a_8_2 * b_2_9;
  assign t0_r8_c9_rr3 = a_8_3 * b_3_9;
  assign t0_r8_c9_rr4 = a_8_4 * b_4_9;
  assign t0_r8_c9_rr5 = a_8_5 * b_5_9;
  assign t0_r8_c9_rr6 = a_8_6 * b_6_9;
  assign t0_r8_c9_rr7 = a_8_7 * b_7_9;
  assign t0_r8_c9_rr8 = a_8_8 * b_8_9;
  assign t0_r8_c9_rr9 = a_8_9 * b_9_9;
  assign t1_r8_c9_rr0 = t0_r8_c9_rr0 + t0_r8_c9_rr1;
  assign t1_r8_c9_rr1 = t0_r8_c9_rr2 + t0_r8_c9_rr3;
  assign t1_r8_c9_rr2 = t0_r8_c9_rr4 + t0_r8_c9_rr5;
  assign t1_r8_c9_rr3 = t0_r8_c9_rr6 + t0_r8_c9_rr7;
  assign t1_r8_c9_rr4 = t0_r8_c9_rr8 + t0_r8_c9_rr9;

  assign t2_r8_c9_rr0 = t1_r8_c9_rr0 + t1_r8_c9_rr1;
  assign t2_r8_c9_rr1 = t1_r8_c9_rr2 + t1_r8_c9_rr3;
  assign t2_r8_c9_rr2 = t1_r8_c9_rr4;

  assign t3_r8_c9_rr0 = t2_r8_c9_rr0 + t2_r8_c9_rr1;
  assign t3_r8_c9_rr1 = t2_r8_c9_rr2;

  assign t4_r8_c9_rr0 = t3_r8_c9_rr0 + t3_r8_c9_rr1;

  assign c_8_9 = t4_r8_c9_rr0;
  assign t0_r9_c0_rr0 = a_9_0 * b_0_0;
  assign t0_r9_c0_rr1 = a_9_1 * b_1_0;
  assign t0_r9_c0_rr2 = a_9_2 * b_2_0;
  assign t0_r9_c0_rr3 = a_9_3 * b_3_0;
  assign t0_r9_c0_rr4 = a_9_4 * b_4_0;
  assign t0_r9_c0_rr5 = a_9_5 * b_5_0;
  assign t0_r9_c0_rr6 = a_9_6 * b_6_0;
  assign t0_r9_c0_rr7 = a_9_7 * b_7_0;
  assign t0_r9_c0_rr8 = a_9_8 * b_8_0;
  assign t0_r9_c0_rr9 = a_9_9 * b_9_0;
  assign t1_r9_c0_rr0 = t0_r9_c0_rr0 + t0_r9_c0_rr1;
  assign t1_r9_c0_rr1 = t0_r9_c0_rr2 + t0_r9_c0_rr3;
  assign t1_r9_c0_rr2 = t0_r9_c0_rr4 + t0_r9_c0_rr5;
  assign t1_r9_c0_rr3 = t0_r9_c0_rr6 + t0_r9_c0_rr7;
  assign t1_r9_c0_rr4 = t0_r9_c0_rr8 + t0_r9_c0_rr9;

  assign t2_r9_c0_rr0 = t1_r9_c0_rr0 + t1_r9_c0_rr1;
  assign t2_r9_c0_rr1 = t1_r9_c0_rr2 + t1_r9_c0_rr3;
  assign t2_r9_c0_rr2 = t1_r9_c0_rr4;

  assign t3_r9_c0_rr0 = t2_r9_c0_rr0 + t2_r9_c0_rr1;
  assign t3_r9_c0_rr1 = t2_r9_c0_rr2;

  assign t4_r9_c0_rr0 = t3_r9_c0_rr0 + t3_r9_c0_rr1;

  assign c_9_0 = t4_r9_c0_rr0;
  assign t0_r9_c1_rr0 = a_9_0 * b_0_1;
  assign t0_r9_c1_rr1 = a_9_1 * b_1_1;
  assign t0_r9_c1_rr2 = a_9_2 * b_2_1;
  assign t0_r9_c1_rr3 = a_9_3 * b_3_1;
  assign t0_r9_c1_rr4 = a_9_4 * b_4_1;
  assign t0_r9_c1_rr5 = a_9_5 * b_5_1;
  assign t0_r9_c1_rr6 = a_9_6 * b_6_1;
  assign t0_r9_c1_rr7 = a_9_7 * b_7_1;
  assign t0_r9_c1_rr8 = a_9_8 * b_8_1;
  assign t0_r9_c1_rr9 = a_9_9 * b_9_1;
  assign t1_r9_c1_rr0 = t0_r9_c1_rr0 + t0_r9_c1_rr1;
  assign t1_r9_c1_rr1 = t0_r9_c1_rr2 + t0_r9_c1_rr3;
  assign t1_r9_c1_rr2 = t0_r9_c1_rr4 + t0_r9_c1_rr5;
  assign t1_r9_c1_rr3 = t0_r9_c1_rr6 + t0_r9_c1_rr7;
  assign t1_r9_c1_rr4 = t0_r9_c1_rr8 + t0_r9_c1_rr9;

  assign t2_r9_c1_rr0 = t1_r9_c1_rr0 + t1_r9_c1_rr1;
  assign t2_r9_c1_rr1 = t1_r9_c1_rr2 + t1_r9_c1_rr3;
  assign t2_r9_c1_rr2 = t1_r9_c1_rr4;

  assign t3_r9_c1_rr0 = t2_r9_c1_rr0 + t2_r9_c1_rr1;
  assign t3_r9_c1_rr1 = t2_r9_c1_rr2;

  assign t4_r9_c1_rr0 = t3_r9_c1_rr0 + t3_r9_c1_rr1;

  assign c_9_1 = t4_r9_c1_rr0;
  assign t0_r9_c2_rr0 = a_9_0 * b_0_2;
  assign t0_r9_c2_rr1 = a_9_1 * b_1_2;
  assign t0_r9_c2_rr2 = a_9_2 * b_2_2;
  assign t0_r9_c2_rr3 = a_9_3 * b_3_2;
  assign t0_r9_c2_rr4 = a_9_4 * b_4_2;
  assign t0_r9_c2_rr5 = a_9_5 * b_5_2;
  assign t0_r9_c2_rr6 = a_9_6 * b_6_2;
  assign t0_r9_c2_rr7 = a_9_7 * b_7_2;
  assign t0_r9_c2_rr8 = a_9_8 * b_8_2;
  assign t0_r9_c2_rr9 = a_9_9 * b_9_2;
  assign t1_r9_c2_rr0 = t0_r9_c2_rr0 + t0_r9_c2_rr1;
  assign t1_r9_c2_rr1 = t0_r9_c2_rr2 + t0_r9_c2_rr3;
  assign t1_r9_c2_rr2 = t0_r9_c2_rr4 + t0_r9_c2_rr5;
  assign t1_r9_c2_rr3 = t0_r9_c2_rr6 + t0_r9_c2_rr7;
  assign t1_r9_c2_rr4 = t0_r9_c2_rr8 + t0_r9_c2_rr9;

  assign t2_r9_c2_rr0 = t1_r9_c2_rr0 + t1_r9_c2_rr1;
  assign t2_r9_c2_rr1 = t1_r9_c2_rr2 + t1_r9_c2_rr3;
  assign t2_r9_c2_rr2 = t1_r9_c2_rr4;

  assign t3_r9_c2_rr0 = t2_r9_c2_rr0 + t2_r9_c2_rr1;
  assign t3_r9_c2_rr1 = t2_r9_c2_rr2;

  assign t4_r9_c2_rr0 = t3_r9_c2_rr0 + t3_r9_c2_rr1;

  assign c_9_2 = t4_r9_c2_rr0;
  assign t0_r9_c3_rr0 = a_9_0 * b_0_3;
  assign t0_r9_c3_rr1 = a_9_1 * b_1_3;
  assign t0_r9_c3_rr2 = a_9_2 * b_2_3;
  assign t0_r9_c3_rr3 = a_9_3 * b_3_3;
  assign t0_r9_c3_rr4 = a_9_4 * b_4_3;
  assign t0_r9_c3_rr5 = a_9_5 * b_5_3;
  assign t0_r9_c3_rr6 = a_9_6 * b_6_3;
  assign t0_r9_c3_rr7 = a_9_7 * b_7_3;
  assign t0_r9_c3_rr8 = a_9_8 * b_8_3;
  assign t0_r9_c3_rr9 = a_9_9 * b_9_3;
  assign t1_r9_c3_rr0 = t0_r9_c3_rr0 + t0_r9_c3_rr1;
  assign t1_r9_c3_rr1 = t0_r9_c3_rr2 + t0_r9_c3_rr3;
  assign t1_r9_c3_rr2 = t0_r9_c3_rr4 + t0_r9_c3_rr5;
  assign t1_r9_c3_rr3 = t0_r9_c3_rr6 + t0_r9_c3_rr7;
  assign t1_r9_c3_rr4 = t0_r9_c3_rr8 + t0_r9_c3_rr9;

  assign t2_r9_c3_rr0 = t1_r9_c3_rr0 + t1_r9_c3_rr1;
  assign t2_r9_c3_rr1 = t1_r9_c3_rr2 + t1_r9_c3_rr3;
  assign t2_r9_c3_rr2 = t1_r9_c3_rr4;

  assign t3_r9_c3_rr0 = t2_r9_c3_rr0 + t2_r9_c3_rr1;
  assign t3_r9_c3_rr1 = t2_r9_c3_rr2;

  assign t4_r9_c3_rr0 = t3_r9_c3_rr0 + t3_r9_c3_rr1;

  assign c_9_3 = t4_r9_c3_rr0;
  assign t0_r9_c4_rr0 = a_9_0 * b_0_4;
  assign t0_r9_c4_rr1 = a_9_1 * b_1_4;
  assign t0_r9_c4_rr2 = a_9_2 * b_2_4;
  assign t0_r9_c4_rr3 = a_9_3 * b_3_4;
  assign t0_r9_c4_rr4 = a_9_4 * b_4_4;
  assign t0_r9_c4_rr5 = a_9_5 * b_5_4;
  assign t0_r9_c4_rr6 = a_9_6 * b_6_4;
  assign t0_r9_c4_rr7 = a_9_7 * b_7_4;
  assign t0_r9_c4_rr8 = a_9_8 * b_8_4;
  assign t0_r9_c4_rr9 = a_9_9 * b_9_4;
  assign t1_r9_c4_rr0 = t0_r9_c4_rr0 + t0_r9_c4_rr1;
  assign t1_r9_c4_rr1 = t0_r9_c4_rr2 + t0_r9_c4_rr3;
  assign t1_r9_c4_rr2 = t0_r9_c4_rr4 + t0_r9_c4_rr5;
  assign t1_r9_c4_rr3 = t0_r9_c4_rr6 + t0_r9_c4_rr7;
  assign t1_r9_c4_rr4 = t0_r9_c4_rr8 + t0_r9_c4_rr9;

  assign t2_r9_c4_rr0 = t1_r9_c4_rr0 + t1_r9_c4_rr1;
  assign t2_r9_c4_rr1 = t1_r9_c4_rr2 + t1_r9_c4_rr3;
  assign t2_r9_c4_rr2 = t1_r9_c4_rr4;

  assign t3_r9_c4_rr0 = t2_r9_c4_rr0 + t2_r9_c4_rr1;
  assign t3_r9_c4_rr1 = t2_r9_c4_rr2;

  assign t4_r9_c4_rr0 = t3_r9_c4_rr0 + t3_r9_c4_rr1;

  assign c_9_4 = t4_r9_c4_rr0;
  assign t0_r9_c5_rr0 = a_9_0 * b_0_5;
  assign t0_r9_c5_rr1 = a_9_1 * b_1_5;
  assign t0_r9_c5_rr2 = a_9_2 * b_2_5;
  assign t0_r9_c5_rr3 = a_9_3 * b_3_5;
  assign t0_r9_c5_rr4 = a_9_4 * b_4_5;
  assign t0_r9_c5_rr5 = a_9_5 * b_5_5;
  assign t0_r9_c5_rr6 = a_9_6 * b_6_5;
  assign t0_r9_c5_rr7 = a_9_7 * b_7_5;
  assign t0_r9_c5_rr8 = a_9_8 * b_8_5;
  assign t0_r9_c5_rr9 = a_9_9 * b_9_5;
  assign t1_r9_c5_rr0 = t0_r9_c5_rr0 + t0_r9_c5_rr1;
  assign t1_r9_c5_rr1 = t0_r9_c5_rr2 + t0_r9_c5_rr3;
  assign t1_r9_c5_rr2 = t0_r9_c5_rr4 + t0_r9_c5_rr5;
  assign t1_r9_c5_rr3 = t0_r9_c5_rr6 + t0_r9_c5_rr7;
  assign t1_r9_c5_rr4 = t0_r9_c5_rr8 + t0_r9_c5_rr9;

  assign t2_r9_c5_rr0 = t1_r9_c5_rr0 + t1_r9_c5_rr1;
  assign t2_r9_c5_rr1 = t1_r9_c5_rr2 + t1_r9_c5_rr3;
  assign t2_r9_c5_rr2 = t1_r9_c5_rr4;

  assign t3_r9_c5_rr0 = t2_r9_c5_rr0 + t2_r9_c5_rr1;
  assign t3_r9_c5_rr1 = t2_r9_c5_rr2;

  assign t4_r9_c5_rr0 = t3_r9_c5_rr0 + t3_r9_c5_rr1;

  assign c_9_5 = t4_r9_c5_rr0;
  assign t0_r9_c6_rr0 = a_9_0 * b_0_6;
  assign t0_r9_c6_rr1 = a_9_1 * b_1_6;
  assign t0_r9_c6_rr2 = a_9_2 * b_2_6;
  assign t0_r9_c6_rr3 = a_9_3 * b_3_6;
  assign t0_r9_c6_rr4 = a_9_4 * b_4_6;
  assign t0_r9_c6_rr5 = a_9_5 * b_5_6;
  assign t0_r9_c6_rr6 = a_9_6 * b_6_6;
  assign t0_r9_c6_rr7 = a_9_7 * b_7_6;
  assign t0_r9_c6_rr8 = a_9_8 * b_8_6;
  assign t0_r9_c6_rr9 = a_9_9 * b_9_6;
  assign t1_r9_c6_rr0 = t0_r9_c6_rr0 + t0_r9_c6_rr1;
  assign t1_r9_c6_rr1 = t0_r9_c6_rr2 + t0_r9_c6_rr3;
  assign t1_r9_c6_rr2 = t0_r9_c6_rr4 + t0_r9_c6_rr5;
  assign t1_r9_c6_rr3 = t0_r9_c6_rr6 + t0_r9_c6_rr7;
  assign t1_r9_c6_rr4 = t0_r9_c6_rr8 + t0_r9_c6_rr9;

  assign t2_r9_c6_rr0 = t1_r9_c6_rr0 + t1_r9_c6_rr1;
  assign t2_r9_c6_rr1 = t1_r9_c6_rr2 + t1_r9_c6_rr3;
  assign t2_r9_c6_rr2 = t1_r9_c6_rr4;

  assign t3_r9_c6_rr0 = t2_r9_c6_rr0 + t2_r9_c6_rr1;
  assign t3_r9_c6_rr1 = t2_r9_c6_rr2;

  assign t4_r9_c6_rr0 = t3_r9_c6_rr0 + t3_r9_c6_rr1;

  assign c_9_6 = t4_r9_c6_rr0;
  assign t0_r9_c7_rr0 = a_9_0 * b_0_7;
  assign t0_r9_c7_rr1 = a_9_1 * b_1_7;
  assign t0_r9_c7_rr2 = a_9_2 * b_2_7;
  assign t0_r9_c7_rr3 = a_9_3 * b_3_7;
  assign t0_r9_c7_rr4 = a_9_4 * b_4_7;
  assign t0_r9_c7_rr5 = a_9_5 * b_5_7;
  assign t0_r9_c7_rr6 = a_9_6 * b_6_7;
  assign t0_r9_c7_rr7 = a_9_7 * b_7_7;
  assign t0_r9_c7_rr8 = a_9_8 * b_8_7;
  assign t0_r9_c7_rr9 = a_9_9 * b_9_7;
  assign t1_r9_c7_rr0 = t0_r9_c7_rr0 + t0_r9_c7_rr1;
  assign t1_r9_c7_rr1 = t0_r9_c7_rr2 + t0_r9_c7_rr3;
  assign t1_r9_c7_rr2 = t0_r9_c7_rr4 + t0_r9_c7_rr5;
  assign t1_r9_c7_rr3 = t0_r9_c7_rr6 + t0_r9_c7_rr7;
  assign t1_r9_c7_rr4 = t0_r9_c7_rr8 + t0_r9_c7_rr9;

  assign t2_r9_c7_rr0 = t1_r9_c7_rr0 + t1_r9_c7_rr1;
  assign t2_r9_c7_rr1 = t1_r9_c7_rr2 + t1_r9_c7_rr3;
  assign t2_r9_c7_rr2 = t1_r9_c7_rr4;

  assign t3_r9_c7_rr0 = t2_r9_c7_rr0 + t2_r9_c7_rr1;
  assign t3_r9_c7_rr1 = t2_r9_c7_rr2;

  assign t4_r9_c7_rr0 = t3_r9_c7_rr0 + t3_r9_c7_rr1;

  assign c_9_7 = t4_r9_c7_rr0;
  assign t0_r9_c8_rr0 = a_9_0 * b_0_8;
  assign t0_r9_c8_rr1 = a_9_1 * b_1_8;
  assign t0_r9_c8_rr2 = a_9_2 * b_2_8;
  assign t0_r9_c8_rr3 = a_9_3 * b_3_8;
  assign t0_r9_c8_rr4 = a_9_4 * b_4_8;
  assign t0_r9_c8_rr5 = a_9_5 * b_5_8;
  assign t0_r9_c8_rr6 = a_9_6 * b_6_8;
  assign t0_r9_c8_rr7 = a_9_7 * b_7_8;
  assign t0_r9_c8_rr8 = a_9_8 * b_8_8;
  assign t0_r9_c8_rr9 = a_9_9 * b_9_8;
  assign t1_r9_c8_rr0 = t0_r9_c8_rr0 + t0_r9_c8_rr1;
  assign t1_r9_c8_rr1 = t0_r9_c8_rr2 + t0_r9_c8_rr3;
  assign t1_r9_c8_rr2 = t0_r9_c8_rr4 + t0_r9_c8_rr5;
  assign t1_r9_c8_rr3 = t0_r9_c8_rr6 + t0_r9_c8_rr7;
  assign t1_r9_c8_rr4 = t0_r9_c8_rr8 + t0_r9_c8_rr9;

  assign t2_r9_c8_rr0 = t1_r9_c8_rr0 + t1_r9_c8_rr1;
  assign t2_r9_c8_rr1 = t1_r9_c8_rr2 + t1_r9_c8_rr3;
  assign t2_r9_c8_rr2 = t1_r9_c8_rr4;

  assign t3_r9_c8_rr0 = t2_r9_c8_rr0 + t2_r9_c8_rr1;
  assign t3_r9_c8_rr1 = t2_r9_c8_rr2;

  assign t4_r9_c8_rr0 = t3_r9_c8_rr0 + t3_r9_c8_rr1;

  assign c_9_8 = t4_r9_c8_rr0;
  assign t0_r9_c9_rr0 = a_9_0 * b_0_9;
  assign t0_r9_c9_rr1 = a_9_1 * b_1_9;
  assign t0_r9_c9_rr2 = a_9_2 * b_2_9;
  assign t0_r9_c9_rr3 = a_9_3 * b_3_9;
  assign t0_r9_c9_rr4 = a_9_4 * b_4_9;
  assign t0_r9_c9_rr5 = a_9_5 * b_5_9;
  assign t0_r9_c9_rr6 = a_9_6 * b_6_9;
  assign t0_r9_c9_rr7 = a_9_7 * b_7_9;
  assign t0_r9_c9_rr8 = a_9_8 * b_8_9;
  assign t0_r9_c9_rr9 = a_9_9 * b_9_9;
  assign t1_r9_c9_rr0 = t0_r9_c9_rr0 + t0_r9_c9_rr1;
  assign t1_r9_c9_rr1 = t0_r9_c9_rr2 + t0_r9_c9_rr3;
  assign t1_r9_c9_rr2 = t0_r9_c9_rr4 + t0_r9_c9_rr5;
  assign t1_r9_c9_rr3 = t0_r9_c9_rr6 + t0_r9_c9_rr7;
  assign t1_r9_c9_rr4 = t0_r9_c9_rr8 + t0_r9_c9_rr9;

  assign t2_r9_c9_rr0 = t1_r9_c9_rr0 + t1_r9_c9_rr1;
  assign t2_r9_c9_rr1 = t1_r9_c9_rr2 + t1_r9_c9_rr3;
  assign t2_r9_c9_rr2 = t1_r9_c9_rr4;

  assign t3_r9_c9_rr0 = t2_r9_c9_rr0 + t2_r9_c9_rr1;
  assign t3_r9_c9_rr1 = t2_r9_c9_rr2;

  assign t4_r9_c9_rr0 = t3_r9_c9_rr0 + t3_r9_c9_rr1;

  assign c_9_9 = t4_r9_c9_rr0;
endmodule
