module multiplier(G11, G12, G14);
  wire _0000_, _0001_, _0002_, _0003_, _0004_, _0005_, _0006_, _0007_, _0008_, _0009_, _0010_, _0011_, _0012_, _0013_, _0014_, _0015_, _0016_, _0017_, _0018_, _0019_, _0020_, _0021_, _0022_, _0023_, _0024_, _0025_, _0026_, _0027_, _0028_, _0029_, _0030_, _0031_, _0032_, _0033_, _0034_, _0035_, _0036_, _0037_, _0038_, _0039_, _0040_, _0041_, _0042_, _0043_, _0044_, _0045_, _0046_, _0047_, _0048_, _0049_, _0050_, _0051_, _0052_, _0053_, _0054_, _0055_, _0056_, _0057_, _0058_, _0059_, _0060_, _0061_, _0062_, _0063_, _0064_, _0065_, _0066_, _0067_, _0068_, _0069_, _0070_, _0071_, _0072_, _0073_, _0074_, _0075_, _0076_, _0077_, _0078_, _0079_, _0080_, _0081_, _0082_, _0083_, _0084_, _0085_, _0086_, _0087_, _0088_, _0089_, _0090_, _0091_, _0092_, _0093_, _0094_, _0095_, _0096_, _0097_, _0098_, _0099_, _0100_, _0101_, _0102_, _0103_, _0104_, _0105_, _0106_, _0107_, _0108_, _0109_, _0110_, _0111_, _0112_, _0113_, _0114_, _0115_, _0116_, _0117_, _0118_, _0119_, _0120_, _0121_, _0122_, _0123_, _0124_, _0125_, _0126_, _0127_, _0128_, _0129_, _0130_, _0131_, _0132_, _0133_, _0134_, _0135_, _0136_, _0137_, _0138_, _0139_, _0140_, _0141_, _0142_, _0143_, _0144_, _0145_, _0146_, _0147_, _0148_, _0149_, _0150_, _0151_, _0152_, _0153_, _0154_, _0155_, _0156_, _0157_, _0158_, _0159_, _0160_, _0161_, _0162_, _0163_, _0164_, _0165_, _0166_, _0167_, _0168_, _0169_, _0170_, _0171_, _0172_, _0173_, _0174_, _0175_, _0176_, _0177_, _0178_, _0179_, _0180_, _0181_, _0182_, _0183_, _0184_, _0185_, _0186_, _0187_, _0188_, _0189_, _0190_, _0191_, _0192_, _0193_, _0194_, _0195_, _0196_, _0197_, _0198_, _0199_, _0200_, _0201_, _0202_, _0203_, _0204_, _0205_, _0206_, _0207_, _0208_, _0209_, _0210_, _0211_, _0212_, _0213_, _0214_, _0215_, _0216_, _0217_, _0218_, _0219_, _0220_, _0221_, _0222_, _0223_, _0224_, _0225_, _0226_, _0227_, _0228_, _0229_, _0230_, _0231_, _0232_, _0233_, _0234_, _0235_, _0236_, _0237_, _0238_, _0239_, _0240_, _0241_, _0242_, _0243_, _0244_, _0245_, _0246_, _0247_, _0248_, _0249_, _0250_, _0251_, _0252_, _0253_, _0254_, _0255_, _0256_, _0257_, _0258_, _0259_, _0260_, _0261_, _0262_, _0263_, _0264_, _0265_, _0266_, _0267_, _0268_, _0269_, _0270_, _0271_, _0272_, _0273_, _0274_, _0275_, _0276_, _0277_, _0278_, _0279_, _0280_, _0281_, _0282_, _0283_, _0284_, _0285_, _0286_, _0287_, _0288_, _0289_, _0290_, _0291_, _0292_, _0293_, _0294_, _0295_, _0296_, _0297_, _0298_, _0299_, _0300_, _0301_, _0302_, _0303_, _0304_, _0305_, _0306_, _0307_, _0308_, _0309_, _0310_, _0311_, _0312_, _0313_, _0314_, _0315_, _0316_, _0317_, _0318_, _0319_, _0320_, _0321_, _0322_, _0323_, _0324_, _0325_, _0326_, _0327_, _0328_, _0329_, _0330_, _0331_, _0332_, _0333_, _0334_, _0335_, _0336_, _0337_, _0338_, _0339_, _0340_, _0341_, _0342_, _0343_, _0344_, _0345_, _0346_, _0347_, _0348_, _0349_, _0350_, _0351_, _0352_, _0353_, _0354_, _0355_, _0356_, _0357_, _0358_, _0359_, _0360_, _0361_, _0362_, _0363_, _0364_, _0365_, _0366_, _0367_, _0368_, _0369_, _0370_, _0371_, _0372_, _0373_, _0374_, _0375_, _0376_, _0377_, _0378_, _0379_, _0380_, _0381_, _0382_, _0383_, _0384_, _0385_, _0386_, _0387_, _0388_, _0389_, _0390_, _0391_, _0392_, _0393_, _0394_, _0395_, _0396_, _0397_, _0398_, _0399_, _0400_, _0401_, _0402_, _0403_, _0404_, _0405_, _0406_, _0407_, _0408_, _0409_, _0410_, _0411_, _0412_, _0413_, _0414_, _0415_, _0416_, _0417_, _0418_, _0419_, _0420_, _0421_, _0422_, _0423_, _0424_, _0425_, _0426_, _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0433_, _0434_, _0435_, _0436_, _0437_, _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_, _0446_, _0447_, _0448_, _0449_, _0450_, _0451_, _0452_, _0453_, _0454_, _0455_, _0456_, _0457_, _0458_, _0459_, _0460_, _0461_, _0462_, _0463_, _0464_, _0465_, _0466_, _0467_, _0468_, _0469_, _0470_, _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_, _0479_, _0480_, _0481_, _0482_, _0483_, _0484_, _0485_, _0486_, _0487_, _0488_, _0489_, _0490_, _0491_, _0492_, _0493_, _0494_, _0495_, _0496_, _0497_, _0498_, _0499_, _0500_, _0501_, _0502_, _0503_, _0504_, _0505_, _0506_, _0507_, _0508_, _0509_, _0510_, _0511_, _0512_, _0513_, _0514_, _0515_, _0516_, _0517_, _0518_, _0519_, _0520_, _0521_, _0522_, _0523_, _0524_, _0525_, _0526_, _0527_, _0528_, _0529_, _0530_, _0531_, _0532_, _0533_, _0534_, _0535_, _0536_, _0537_, _0538_, _0539_, _0540_, _0541_, _0542_, _0543_, _0544_, _0545_, _0546_, _0547_, _0548_, _0549_, _0550_, _0551_, _0552_, _0553_, _0554_, _0555_, _0556_, _0557_, _0558_, _0559_, _0560_, _0561_, _0562_, _0563_, _0564_, _0565_, _0566_, _0567_, _0568_, _0569_, _0570_, _0571_, _0572_, _0573_, _0574_, _0575_, _0576_, _0577_, _0578_, _0579_, _0580_, _0581_, _0582_, _0583_, _0584_, _0585_, _0586_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_, _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0602_, _0603_, _0604_, _0605_, _0606_, _0607_, _0608_, _0609_, _0610_, _0611_, _0612_, _0613_, _0614_, _0615_, _0616_, _0617_, _0618_, _0619_, _0620_, _0621_, _0622_, _0623_, _0624_, _0625_, _0626_, _0627_, _0628_, _0629_, _0630_, _0631_, _0632_, _0633_, _0634_, _0635_, _0636_, _0637_, _0638_, _0639_, _0640_, _0641_, _0642_, _0643_, _0644_, _0645_, _0646_, _0647_, _0648_, _0649_, _0650_, _0651_, _0652_, _0653_, _0654_, _0655_, _0656_, _0657_, _0658_, _0659_, _0660_, _0661_, _0662_, _0663_, _0664_, _0665_, _0666_, _0667_, _0668_, _0669_, _0670_, _0671_, _0672_, _0673_, _0674_, _0675_, _0676_, _0677_, _0678_, _0679_, _0680_, _0681_, _0682_, _0683_, _0684_, _0685_, _0686_, _0687_, _0688_, _0689_, _0690_, _0691_, _0692_, _0693_, _0694_, _0695_, _0696_, _0697_, _0698_, _0699_, _0700_, _0701_, _0702_, _0703_, _0704_, _0705_, _0706_, _0707_, _0708_, _0709_, _0710_, _0711_, _0712_, _0713_, _0714_, _0715_, _0716_, _0717_, _0718_, _0719_, _0720_, _0721_, _0722_, _0723_, _0724_, _0725_, _0726_, _0727_, _0728_, _0729_, _0730_, _0731_, _0732_, _0733_, _0734_, _0735_, _0736_, _0737_, _0738_, _0739_, _0740_, _0741_, _0742_, _0743_, _0744_, _0745_, _0746_, _0747_, _0748_, _0749_, _0750_, _0751_, _0752_, _0753_, _0754_, _0755_, _0756_, _0757_, _0758_, _0759_, _0760_, _0761_, _0762_, _0763_, _0764_, _0765_, _0766_, _0767_, _0768_, _0769_, _0770_, _0771_, _0772_, _0773_, _0774_, _0775_, _0776_, _0777_, _0778_, _0779_, _0780_, _0781_, _0782_, _0783_, _0784_, _0785_, _0786_, _0787_, _0788_, _0789_, _0790_, _0791_, _0792_, _0793_, _0794_, _0795_, _0796_, _0797_, _0798_, _0799_, _0800_, _0801_, _0802_, _0803_, _0804_, _0805_, _0806_, _0807_, _0808_, _0809_, _0810_, _0811_, _0812_, _0813_, _0814_, _0815_, _0816_, _0817_, _0818_, _0819_, _0820_, _0821_, _0822_, _0823_, _0824_, _0825_, _0826_, _0827_, _0828_, _0829_, _0830_, _0831_, _0832_, _0833_, _0834_, _0835_, _0836_, _0837_, _0838_, _0839_, _0840_, _0841_, _0842_, _0843_, _0844_, _0845_, _0846_, _0847_, _0848_, _0849_, _0850_, _0851_, _0852_, _0853_, _0854_, _0855_, _0856_, _0857_, _0858_, _0859_, _0860_, _0861_, _0862_, _0863_, _0864_, _0865_, _0866_, _0867_, _0868_, _0869_, _0870_, _0871_, _0872_, _0873_, _0874_, _0875_, _0876_, _0877_, _0878_, _0879_, _0880_, _0881_, _0882_, _0883_, _0884_, _0885_, _0886_, _0887_, _0888_, _0889_, _0890_, _0891_, _0892_, _0893_, _0894_, _0895_, _0896_, _0897_, _0898_, _0899_, _0900_, _0901_, _0902_, _0903_, _0904_, _0905_, _0906_, _0907_, _0908_, _0909_, _0910_, _0911_, _0912_, _0913_, _0914_, _0915_, _0916_, _0917_, _0918_, _0919_, _0920_, _0921_, _0922_, _0923_, _0924_, _0925_, _0926_, _0927_, _0928_, _0929_, _0930_, _0931_, _0932_, _0933_, _0934_, _0935_, _0936_, _0937_, _0938_, _0939_, _0940_, _0941_, _0942_, _0943_, _0944_, _0945_, _0946_, _0947_, _0948_, _0949_, _0950_, _0951_, _0952_, _0953_, _0954_, _0955_, _0956_, _0957_, _0958_, _0959_, _0960_, _0961_, _0962_, _0963_, _0964_, _0965_, _0966_, _0967_, _0968_, _0969_, _0970_, _0971_, _0972_, _0973_, _0974_, _0975_, _0976_, _0977_, _0978_, _0979_, _0980_, _0981_, _0982_, _0983_, _0984_, _0985_, _0986_, _0987_, _0988_, _0989_, _0990_, _0991_, _0992_, _0993_, _0994_, _0995_, _0996_, _0997_, _0998_, _0999_, _1000_, _1001_, _1002_, _1003_, _1004_, _1005_, _1006_, _1007_, _1008_, _1009_, _1010_, _1011_, _1012_, _1013_, _1014_, _1015_, _1016_, _1017_, _1018_, _1019_, _1020_, _1021_, _1022_, _1023_, _1024_, _1025_, _1026_, _1027_, _1028_, _1029_, _1030_, _1031_, _1032_, _1033_, _1034_, _1035_, _1036_, _1037_, _1038_, _1039_, _1040_, _1041_, _1042_, _1043_, _1044_, _1045_, _1046_, _1047_, _1048_, _1049_, _1050_, _1051_, _1052_, _1053_, _1054_, _1055_, _1056_, _1057_, _1058_, _1059_, _1060_, _1061_, _1062_, _1063_, _1064_, _1065_, _1066_, _1067_, _1068_, _1069_, _1070_, _1071_, _1072_, _1073_, _1074_, _1075_, _1076_, _1077_, _1078_, _1079_, _1080_, _1081_, _1082_, _1083_, _1084_, _1085_, _1086_, _1087_, _1088_, _1089_, _1090_, _1091_, _1092_, _1093_, _1094_, _1095_, _1096_, _1097_, _1098_, _1099_, _1100_, _1101_, _1102_, _1103_, _1104_, _1105_, _1106_, _1107_, _1108_, _1109_, _1110_, _1111_, _1112_, _1113_, _1114_, _1115_, _1116_, _1117_, _1118_, _1119_, _1120_, _1121_, _1122_, _1123_, _1124_, _1125_, _1126_, _1127_, _1128_, _1129_, _1130_, _1131_, _1132_, _1133_, _1134_, _1135_, _1136_, _1137_, _1138_, _1139_, _1140_, _1141_, _1142_, _1143_, _1144_, _1145_, _1146_, _1147_, _1148_, _1149_, _1150_, _1151_, _1152_, _1153_, _1154_, _1155_, _1156_, _1157_, _1158_, _1159_, _1160_, _1161_, _1162_, _1163_, _1164_, _1165_, _1166_, _1167_, _1168_, _1169_, _1170_, _1171_, _1172_, _1173_, _1174_, _1175_, _1176_, _1177_, _1178_, _1179_, _1180_, _1181_, _1182_, _1183_, _1184_, _1185_, _1186_, _1187_, _1188_, _1189_, _1190_, _1191_, _1192_, _1193_, _1194_, _1195_, _1196_, _1197_, _1198_, _1199_, _1200_, _1201_, _1202_, _1203_, _1204_, _1205_, _1206_, _1207_, _1208_, _1209_, _1210_, _1211_, _1212_, _1213_, _1214_, _1215_, _1216_, _1217_, _1218_, _1219_, _1220_, _1221_, _1222_, _1223_, _1224_, _1225_, _1226_, _1227_, _1228_, _1229_, _1230_, _1231_, _1232_, _1233_, _1234_, _1235_, _1236_, _1237_, _1238_, _1239_, _1240_, _1241_, _1242_, _1243_, _1244_, _1245_, _1246_, _1247_, _1248_, _1249_, _1250_, _1251_, _1252_, _1253_, _1254_, _1255_, _1256_, _1257_, _1258_, _1259_, _1260_, _1261_, _1262_, _1263_, _1264_, _1265_, _1266_, _1267_, _1268_, _1269_, _1270_, _1271_, _1272_, _1273_, _1274_, _1275_, _1276_, _1277_, _1278_, _1279_, _1280_, _1281_, _1282_, _1283_, _1284_, _1285_, _1286_, _1287_, _1288_, _1289_, _1290_, _1291_, _1292_, _1293_, _1294_, _1295_, _1296_, _1297_, _1298_, _1299_, _1300_, _1301_, _1302_, _1303_, _1304_, _1305_, _1306_, _1307_, _1308_, _1309_, _1310_, _1311_, _1312_, _1313_, _1314_, _1315_, _1316_, _1317_, _1318_, _1319_, _1320_, _1321_, _1322_, _1323_, _1324_, _1325_, _1326_, _1327_, _1328_, _1329_, _1330_, _1331_, _1332_, _1333_, _1334_, _1335_, _1336_, _1337_, _1338_, _1339_, _1340_, _1341_, _1342_, _1343_, _1344_, _1345_, _1346_, _1347_, _1348_, _1349_, _1350_, _1351_, _1352_, _1353_, _1354_, _1355_, _1356_, _1357_, _1358_, _1359_, _1360_, _1361_, _1362_, _1363_, _1364_, _1365_, _1366_, _1367_, _1368_, _1369_, _1370_, _1371_, _1372_, _1373_, _1374_, _1375_, _1376_, _1377_, _1378_, _1379_, _1380_, _1381_, _1382_, _1383_, _1384_, _1385_, _1386_, _1387_, _1388_, _1389_, _1390_, _1391_, _1392_, _1393_, _1394_, _1395_, _1396_, _1397_, _1398_, _1399_, _1400_, _1401_, _1402_, _1403_, _1404_, _1405_, _1406_, _1407_, _1408_, _1409_, _1410_, _1411_, _1412_, _1413_, _1414_, _1415_, _1416_, _1417_, _1418_, _1419_, _1420_, _1421_, _1422_, _1423_, _1424_, _1425_, _1426_, _1427_, _1428_, _1429_, _1430_, _1431_, _1432_, _1433_, _1434_, _1435_, _1436_, _1437_, _1438_, _1439_, _1440_, _1441_, _1442_, _1443_, _1444_, _1445_, _1446_, _1447_, _1448_, _1449_, _1450_, _1451_, _1452_, _1453_, _1454_, _1455_, _1456_, _1457_, _1458_, _1459_, _1460_, _1461_, _1462_, _1463_, _1464_, _1465_, _1466_, _1467_, _1468_, _1469_, _1470_, _1471_, _1472_, _1473_, _1474_, _1475_, _1476_, _1477_, _1478_, _1479_, _1480_, _1481_, _1482_, _1483_, _1484_, _1485_, _1486_, _1487_, _1488_, _1489_, _1490_, _1491_, _1492_, _1493_, _1494_, _1495_, _1496_, _1497_, _1498_, _1499_, _1500_, _1501_, _1502_, _1503_, _1504_, _1505_, _1506_, _1507_, _1508_, _1509_, _1510_, _1511_, _1512_, _1513_, _1514_, _1515_, _1516_, _1517_, _1518_, _1519_, _1520_, _1521_, _1522_, _1523_, _1524_, _1525_, _1526_, _1527_, _1528_, _1529_, _1530_, _1531_, _1532_, _1533_, _1534_, _1535_, _1536_, _1537_, _1538_, _1539_, _1540_, _1541_, _1542_, _1543_, _1544_, _1545_, _1546_, _1547_, _1548_, _1549_, _1550_, _1551_, _1552_, _1553_, _1554_, _1555_, _1556_, _1557_, _1558_, _1559_, _1560_, _1561_, _1562_, _1563_, _1564_, _1565_, _1566_, _1567_, _1568_, _1569_, _1570_, _1571_, _1572_, _1573_, _1574_, _1575_, _1576_, _1577_, _1578_, _1579_, _1580_, _1581_, _1582_, _1583_, _1584_, _1585_, _1586_, _1587_, _1588_, _1589_, _1590_, _1591_, _1592_, _1593_, _1594_, _1595_, _1596_, _1597_, _1598_, _1599_, _1600_, _1601_, _1602_, _1603_, _1604_, _1605_, _1606_, _1607_, _1608_, _1609_, _1610_, _1611_, _1612_, _1613_, _1614_, _1615_, _1616_, _1617_, _1618_, _1619_, _1620_, _1621_, _1622_, _1623_, _1624_, _1625_, _1626_, _1627_, _1628_, _1629_, _1630_, _1631_, _1632_, _1633_, _1634_, _1635_, _1636_, _1637_, _1638_, _1639_, _1640_, _1641_, _1642_, _1643_, _1644_, _1645_, _1646_, _1647_, _1648_, _1649_, _1650_, _1651_, _1652_, _1653_, _1654_, _1655_, _1656_, _1657_, _1658_, _1659_, _1660_, _1661_, _1662_, _1663_, _1664_, _1665_, _1666_, _1667_, _1668_, _1669_, _1670_, _1671_, _1672_, _1673_, _1674_, _1675_, _1676_, _1677_, _1678_, _1679_, _1680_, _1681_, _1682_, _1683_, _1684_, _1685_, _1686_, _1687_, _1688_, _1689_, _1690_, _1691_, _1692_, _1693_, _1694_, _1695_, _1696_, _1697_, _1698_, _1699_, _1700_, _1701_, _1702_, _1703_, _1704_, _1705_, _1706_, _1707_, _1708_, _1709_, _1710_, _1711_, _1712_, _1713_, _1714_, _1715_, _1716_, _1717_, _1718_, _1719_, _1720_, _1721_, _1722_, _1723_, _1724_, _1725_, _1726_, _1727_, _1728_, _1729_, _1730_, _1731_, _1732_, _1733_, _1734_, _1735_, _1736_, _1737_, _1738_, _1739_, _1740_, _1741_, _1742_, _1743_, _1744_, _1745_, _1746_, _1747_, _1748_, _1749_, _1750_, _1751_, _1752_, _1753_, _1754_, _1755_, _1756_, _1757_, _1758_, _1759_, _1760_, _1761_, _1762_, _1763_, _1764_, _1765_, _1766_, _1767_, _1768_, _1769_, _1770_, _1771_, _1772_, _1773_, _1774_, _1775_, _1776_, _1777_, _1778_, _1779_, _1780_, _1781_, _1782_, _1783_, _1784_, _1785_, _1786_, _1787_, _1788_, _1789_, _1790_, _1791_, _1792_, _1793_, _1794_, _1795_, _1796_, _1797_, _1798_, _1799_, _1800_, _1801_, _1802_, _1803_, _1804_, _1805_, _1806_, _1807_, _1808_, _1809_, _1810_, _1811_, _1812_, _1813_, _1814_, _1815_, _1816_, _1817_, _1818_, _1819_, _1820_, _1821_, _1822_, _1823_, _1824_, _1825_, _1826_, _1827_, _1828_, _1829_, _1830_, _1831_, _1832_, _1833_, _1834_, _1835_, _1836_, _1837_, _1838_, _1839_, _1840_, _1841_, _1842_, _1843_, _1844_, _1845_, _1846_, _1847_, _1848_, _1849_, _1850_, _1851_, _1852_, _1853_, _1854_, _1855_, _1856_, _1857_, _1858_, _1859_, _1860_, _1861_, _1862_, _1863_, _1864_, _1865_, _1866_, _1867_, _1868_, _1869_, _1870_, _1871_, _1872_, _1873_, _1874_, _1875_, _1876_, _1877_, _1878_, _1879_, _1880_, _1881_, _1882_, _1883_, _1884_, _1885_, _1886_, _1887_, _1888_, _1889_, _1890_, _1891_, _1892_, _1893_, _1894_, _1895_, _1896_, _1897_, _1898_, _1899_, _1900_, _1901_, _1902_, _1903_, _1904_, _1905_, _1906_, _1907_, _1908_, _1909_, _1910_, _1911_, _1912_, _1913_, _1914_, _1915_, _1916_, _1917_, _1918_, _1919_, _1920_, _1921_, _1922_, _1923_, _1924_, _1925_, _1926_, _1927_, _1928_, _1929_, _1930_, _1931_, _1932_, _1933_, _1934_, _1935_, _1936_, _1937_, _1938_, _1939_, _1940_, _1941_, _1942_, _1943_, _1944_, _1945_, _1946_, _1947_, _1948_, _1949_, _1950_, _1951_, _1952_, _1953_, _1954_, _1955_, _1956_, _1957_, _1958_, _1959_, _1960_, _1961_, _1962_, _1963_, _1964_, _1965_, _1966_, _1967_, _1968_, _1969_, _1970_, _1971_, _1972_, _1973_, _1974_, _1975_, _1976_, _1977_, _1978_, _1979_, _1980_, _1981_, _1982_, _1983_, _1984_, _1985_, _1986_, _1987_, _1988_, _1989_, _1990_, _1991_, _1992_, _1993_, _1994_, _1995_, _1996_, _1997_, _1998_, _1999_, _2000_, _2001_, _2002_, _2003_, _2004_, _2005_, _2006_, _2007_, _2008_, _2009_, _2010_, _2011_, _2012_, _2013_, _2014_, _2015_, _2016_, _2017_, _2018_, _2019_, _2020_, _2021_, _2022_, _2023_, _2024_, _2025_, _2026_, _2027_, _2028_, _2029_, _2030_, _2031_, _2032_, _2033_, _2034_, _2035_, _2036_, _2037_, _2038_, _2039_, _2040_, _2041_, _2042_, _2043_, _2044_, _2045_, _2046_, _2047_, _2048_, _2049_, _2050_, _2051_, _2052_, _2053_, _2054_, _2055_, _2056_, _2057_, _2058_, _2059_, _2060_, _2061_, _2062_, _2063_, _2064_, _2065_, _2066_, _2067_, _2068_, _2069_, _2070_, _2071_, _2072_, _2073_, _2074_, _2075_, _2076_, _2077_, _2078_, _2079_, _2080_, _2081_, _2082_, _2083_, _2084_, _2085_, _2086_, _2087_, _2088_, _2089_, _2090_, _2091_, _2092_, _2093_, _2094_, _2095_, _2096_, _2097_, _2098_, _2099_, _2100_, _2101_, _2102_, _2103_, _2104_, _2105_, _2106_, _2107_, _2108_, _2109_, _2110_, _2111_, _2112_, _2113_, _2114_, _2115_, _2116_, _2117_, _2118_, _2119_, _2120_, _2121_, _2122_, _2123_, _2124_, _2125_, _2126_, _2127_, _2128_, _2129_, _2130_, _2131_, _2132_, _2133_, _2134_, _2135_, _2136_, _2137_, _2138_, _2139_, _2140_, _2141_, _2142_, _2143_, _2144_, _2145_, _2146_, _2147_, _2148_, _2149_, _2150_, _2151_, _2152_, _2153_, _2154_, _2155_, _2156_, _2157_, _2158_, _2159_, _2160_, _2161_, _2162_, _2163_, _2164_, _2165_, _2166_, _2167_, _2168_, _2169_, _2170_, _2171_, _2172_, _2173_, _2174_, _2175_, _2176_, _2177_, _2178_, _2179_, _2180_, _2181_, _2182_, _2183_, _2184_, _2185_, _2186_, _2187_, _2188_, _2189_, _2190_, _2191_, _2192_, _2193_, _2194_, _2195_, _2196_, _2197_, _2198_, _2199_, _2200_, _2201_, _2202_, _2203_, _2204_, _2205_, _2206_, _2207_, _2208_, _2209_, _2210_, _2211_, _2212_, _2213_, _2214_, _2215_, _2216_, _2217_, _2218_, _2219_, _2220_, _2221_, _2222_, _2223_, _2224_, _2225_, _2226_, _2227_, _2228_, _2229_, _2230_, _2231_, _2232_, _2233_, _2234_, _2235_, _2236_, _2237_, _2238_, _2239_, _2240_, _2241_, _2242_, _2243_, _2244_, _2245_, _2246_, _2247_, _2248_, _2249_, _2250_, _2251_, _2252_, _2253_, _2254_, _2255_, _2256_, _2257_, _2258_, _2259_, _2260_, _2261_, _2262_, _2263_, _2264_, _2265_, _2266_, _2267_, _2268_, _2269_, _2270_, _2271_, _2272_, _2273_, _2274_, _2275_, _2276_, _2277_, _2278_, _2279_, _2280_, _2281_, _2282_, _2283_, _2284_, _2285_, _2286_, _2287_, _2288_, _2289_, _2290_, _2291_, _2292_, _2293_, _2294_, _2295_, _2296_, _2297_, _2298_, _2299_, _2300_, _2301_, _2302_, _2303_, _2304_, _2305_, _2306_, _2307_, _2308_, _2309_, _2310_, _2311_, _2312_, _2313_, _2314_, _2315_, _2316_, _2317_, _2318_, _2319_, _2320_, _2321_, _2322_, _2323_, _2324_, _2325_, _2326_, _2327_, _2328_, _2329_, _2330_, _2331_, _2332_, _2333_, _2334_, _2335_, _2336_, _2337_, _2338_, _2339_, _2340_, _2341_, _2342_, _2343_, _2344_, _2345_, _2346_, _2347_, _2348_, _2349_, _2350_, _2351_, _2352_, _2353_, _2354_, _2355_, _2356_, _2357_, _2358_, _2359_, _2360_, _2361_, _2362_, _2363_, _2364_, _2365_, _2366_, _2367_, _2368_, _2369_, _2370_, _2371_, _2372_, _2373_, _2374_, _2375_, _2376_, _2377_, _2378_, _2379_, _2380_, _2381_, _2382_, _2383_, _2384_, _2385_, _2386_, _2387_, _2388_, _2389_, _2390_, _2391_, _2392_, _2393_, _2394_, _2395_, _2396_, _2397_, _2398_, _2399_, _2400_, _2401_, _2402_, _2403_, _2404_, _2405_, _2406_, _2407_, _2408_, _2409_, _2410_, _2411_, _2412_, _2413_, _2414_, _2415_, _2416_, _2417_, _2418_, _2419_, _2420_, _2421_, _2422_, _2423_, _2424_, _2425_, _2426_, _2427_, _2428_, _2429_, _2430_, _2431_, _2432_, _2433_, _2434_, _2435_, _2436_, _2437_, _2438_, _2439_, _2440_, _2441_, _2442_, _2443_, _2444_, _2445_, _2446_, _2447_, _2448_, _2449_, _2450_, _2451_, _2452_, _2453_, _2454_, _2455_, _2456_, _2457_, _2458_, _2459_, _2460_, _2461_, _2462_, _2463_, _2464_, _2465_, _2466_, _2467_, _2468_, _2469_, _2470_, _2471_, _2472_, _2473_, _2474_, _2475_, _2476_, _2477_, _2478_, _2479_, _2480_, _2481_, _2482_, _2483_, _2484_, _2485_, _2486_, _2487_, _2488_, _2489_, _2490_, _2491_, _2492_, _2493_, _2494_, _2495_, _2496_, _2497_, _2498_, _2499_, _2500_, _2501_, _2502_, _2503_, _2504_, _2505_, _2506_, _2507_, _2508_, _2509_, _2510_, _2511_, _2512_, _2513_, _2514_, _2515_, _2516_, _2517_, _2518_, _2519_, _2520_, _2521_, _2522_, _2523_, _2524_, _2525_, _2526_, _2527_, _2528_, _2529_, _2530_, _2531_, _2532_, _2533_, _2534_, _2535_, _2536_, _2537_, _2538_, _2539_, _2540_, _2541_, _2542_, _2543_, _2544_, _2545_, _2546_, _2547_, _2548_, _2549_, _2550_, _2551_, _2552_, _2553_, _2554_, _2555_, _2556_, _2557_, _2558_, _2559_, _2560_, _2561_, _2562_, _2563_, _2564_, _2565_, _2566_, _2567_, _2568_, _2569_, _2570_, _2571_, _2572_, _2573_, _2574_, _2575_, _2576_, _2577_, _2578_, _2579_, _2580_, _2581_, _2582_, _2583_, _2584_, _2585_, _2586_, _2587_, _2588_, _2589_, _2590_, _2591_, _2592_, _2593_, _2594_, _2595_, _2596_, _2597_, _2598_, _2599_, _2600_, _2601_, _2602_, _2603_, _2604_, _2605_, _2606_, _2607_, _2608_, _2609_, _2610_, _2611_, _2612_, _2613_, _2614_, _2615_, _2616_, _2617_, _2618_, _2619_, _2620_, _2621_, _2622_, _2623_, _2624_, _2625_, _2626_, _2627_, _2628_, _2629_, _2630_, _2631_, _2632_, _2633_, _2634_, _2635_, _2636_, _2637_, _2638_, _2639_, _2640_, _2641_, _2642_, _2643_, _2644_, _2645_, _2646_, _2647_, _2648_, _2649_, _2650_, _2651_, _2652_, _2653_, _2654_, _2655_, _2656_, _2657_, _2658_, _2659_, _2660_, _2661_, _2662_, _2663_, _2664_, _2665_, _2666_, _2667_, _2668_, _2669_, _2670_, _2671_, _2672_, _2673_, _2674_, _2675_, _2676_, _2677_, _2678_, _2679_, _2680_, _2681_, _2682_, _2683_, _2684_, _2685_, _2686_, _2687_, _2688_, _2689_, _2690_, _2691_, _2692_, _2693_, _2694_, _2695_, _2696_, _2697_, _2698_, _2699_, _2700_, _2701_, _2702_, _2703_, _2704_, _2705_, _2706_, _2707_, _2708_, _2709_, _2710_, _2711_, _2712_, _2713_, _2714_, _2715_, _2716_, _2717_, _2718_, _2719_, _2720_, _2721_, _2722_, _2723_, _2724_, _2725_, _2726_, _2727_, _2728_, _2729_, _2730_, _2731_, _2732_, _2733_, _2734_, _2735_, _2736_, _2737_, _2738_, _2739_, _2740_, _2741_, _2742_, _2743_, _2744_, _2745_, _2746_, _2747_, _2748_, _2749_, _2750_, _2751_, _2752_, _2753_, _2754_, _2755_, _2756_, _2757_, _2758_, _2759_, _2760_, _2761_, _2762_, _2763_, _2764_, _2765_, _2766_, _2767_, _2768_, _2769_, _2770_, _2771_, _2772_, _2773_, _2774_, _2775_, _2776_, _2777_, _2778_, _2779_, _2780_, _2781_, _2782_, _2783_, _2784_, _2785_, _2786_, _2787_, _2788_, _2789_, _2790_, _2791_, _2792_, _2793_, _2794_, _2795_, _2796_, _2797_, _2798_, _2799_, _2800_, _2801_, _2802_, _2803_, _2804_, _2805_, _2806_, _2807_, _2808_, _2809_, _2810_, _2811_, _2812_, _2813_, _2814_, _2815_, _2816_, _2817_, _2818_, _2819_, _2820_, _2821_, _2822_, _2823_, _2824_, _2825_, _2826_, _2827_, _2828_, _2829_, _2830_, _2831_, _2832_, _2833_, _2834_, _2835_, _2836_, _2837_, _2838_, _2839_, _2840_, _2841_, _2842_, _2843_, _2844_, _2845_, _2846_, _2847_, _2848_, _2849_, _2850_, _2851_, _2852_, _2853_, _2854_, _2855_, _2856_, _2857_, _2858_, _2859_, _2860_, _2861_, _2862_, _2863_, _2864_, _2865_, _2866_, _2867_, _2868_, _2869_, _2870_, _2871_, _2872_, _2873_, _2874_, _2875_, _2876_, _2877_, _2878_, _2879_, _2880_, _2881_, _2882_, _2883_, _2884_, _2885_, _2886_, _2887_, _2888_, _2889_, _2890_, _2891_, _2892_, _2893_, _2894_, _2895_, _2896_, _2897_, _2898_, _2899_, _2900_, _2901_, _2902_, _2903_, _2904_, _2905_, _2906_, _2907_, _2908_, _2909_, _2910_, _2911_, _2912_, _2913_, _2914_, _2915_, _2916_, _2917_, _2918_, _2919_, _2920_, _2921_, _2922_, _2923_, _2924_, _2925_, _2926_, _2927_, _2928_, _2929_, _2930_, _2931_, _2932_, _2933_, _2934_, _2935_, _2936_, _2937_, _2938_, _2939_, _2940_, _2941_, _2942_, _2943_, _2944_, _2945_, _2946_, _2947_, _2948_, _2949_, _2950_, _2951_, _2952_, _2953_, _2954_, _2955_, _2956_, _2957_, _2958_, _2959_, _2960_, _2961_, _2962_, _2963_, _2964_, _2965_, _2966_, _2967_, _2968_, _2969_, _2970_, _2971_, _2972_, _2973_, _2974_, _2975_, _2976_, _2977_, _2978_, _2979_, _2980_, _2981_, _2982_, _2983_, _2984_, _2985_, _2986_, _2987_, _2988_, _2989_, _2990_, _2991_, _2992_, _2993_, _2994_, _2995_, _2996_, _2997_, _2998_, _2999_, _3000_, _3001_, _3002_, _3003_, _3004_, _3005_, _3006_, _3007_, _3008_, _3009_, _3010_, _3011_, _3012_, _3013_, _3014_, _3015_, _3016_, _3017_, _3018_, _3019_, _3020_, _3021_, _3022_, _3023_, _3024_, _3025_, _3026_, _3027_, _3028_, _3029_, _3030_, _3031_, _3032_, _3033_, _3034_, _3035_, _3036_, _3037_, _3038_, _3039_, _3040_, _3041_, _3042_, _3043_, _3044_, _3045_, _3046_, _3047_, _3048_, _3049_, _3050_, _3051_, _3052_, _3053_, _3054_, _3055_, _3056_, _3057_, _3058_, _3059_, _3060_, _3061_, _3062_, _3063_, _3064_, _3065_, _3066_, _3067_, _3068_, _3069_, _3070_, _3071_, _3072_, _3073_, _3074_, _3075_, _3076_, _3077_, _3078_, _3079_, _3080_, _3081_, _3082_, _3083_, _3084_, _3085_, _3086_, _3087_, _3088_, _3089_, _3090_, _3091_, _3092_, _3093_, _3094_, _3095_, _3096_, _3097_, _3098_, _3099_, _3100_, _3101_, _3102_, _3103_, _3104_, _3105_, _3106_, _3107_, _3108_, _3109_, _3110_, _3111_, _3112_, _3113_, _3114_, _3115_, _3116_, _3117_, _3118_, _3119_, _3120_, _3121_, _3122_, _3123_, _3124_, _3125_, _3126_, _3127_, _3128_, _3129_, _3130_, _3131_, _3132_, _3133_, _3134_, _3135_, _3136_, _3137_, _3138_, _3139_, _3140_, _3141_, _3142_, _3143_, _3144_, _3145_, _3146_, _3147_, _3148_, _3149_, _3150_, _3151_, _3152_, _3153_, _3154_, _3155_, _3156_, _3157_, _3158_, _3159_, _3160_, _3161_, _3162_, _3163_, _3164_, _3165_, _3166_, _3167_, _3168_, _3169_, _3170_, _3171_, _3172_, _3173_, _3174_, _3175_, _3176_, _3177_, _3178_, _3179_, _3180_, _3181_, _3182_, _3183_, _3184_, _3185_, _3186_, _3187_, _3188_, _3189_, _3190_, _3191_, _3192_, _3193_, _3194_, _3195_, _3196_, _3197_, _3198_, _3199_, _3200_, _3201_, _3202_, _3203_, _3204_, _3205_, _3206_, _3207_, _3208_, _3209_, _3210_, _3211_, _3212_, _3213_, _3214_, _3215_, _3216_, _3217_, _3218_, _3219_, _3220_, _3221_, _3222_, _3223_, _3224_, _3225_, _3226_, _3227_, _3228_, _3229_, _3230_, _3231_, _3232_, _3233_, _3234_, _3235_, _3236_, _3237_, _3238_, _3239_, _3240_, _3241_, _3242_, _3243_, _3244_, _3245_, _3246_, _3247_, _3248_, _3249_, _3250_, _3251_, _3252_, _3253_, _3254_, _3255_, _3256_, _3257_, _3258_, _3259_, _3260_, _3261_, _3262_, _3263_, _3264_, _3265_, _3266_, _3267_, _3268_, _3269_, _3270_, _3271_, _3272_, _3273_, _3274_, _3275_, _3276_, _3277_, _3278_, _3279_, _3280_, _3281_, _3282_, _3283_, _3284_, _3285_, _3286_, _3287_, _3288_, _3289_, _3290_, _3291_, _3292_, _3293_, _3294_, _3295_, _3296_, _3297_, _3298_, _3299_, _3300_, _3301_, _3302_, _3303_, _3304_, _3305_, _3306_, _3307_, _3308_, _3309_, _3310_, _3311_, _3312_, _3313_, _3314_, _3315_, _3316_, _3317_, _3318_, _3319_, _3320_, _3321_, _3322_, _3323_, _3324_, _3325_, _3326_, _3327_, _3328_, _3329_, _3330_, _3331_, _3332_, _3333_, _3334_, _3335_, _3336_, _3337_, _3338_, _3339_, _3340_, _3341_, _3342_, _3343_, _3344_, _3345_, _3346_, _3347_, _3348_, _3349_, _3350_, _3351_, _3352_, _3353_, _3354_, _3355_, _3356_, _3357_, _3358_, _3359_, _3360_, _3361_, _3362_, _3363_, _3364_, _3365_, _3366_, _3367_, _3368_, _3369_, _3370_, _3371_, _3372_, _3373_, _3374_, _3375_, _3376_, _3377_, _3378_, _3379_, _3380_, _3381_, _3382_, _3383_, _3384_, _3385_, _3386_, _3387_, _3388_, _3389_, _3390_, _3391_, _3392_, _3393_, _3394_, _3395_, _3396_, _3397_, _3398_, _3399_, _3400_, _3401_, _3402_, _3403_, _3404_, _3405_, _3406_, _3407_, _3408_, _3409_, _3410_, _3411_, _3412_, _3413_, _3414_, _3415_, _3416_, _3417_, _3418_, _3419_, _3420_, _3421_, _3422_, _3423_, _3424_, _3425_, _3426_, _3427_, _3428_, _3429_, _3430_, _3431_, _3432_, _3433_, _3434_, _3435_, _3436_, _3437_, _3438_, _3439_, _3440_, _3441_, _3442_, _3443_, _3444_, _3445_, _3446_, _3447_, _3448_, _3449_, _3450_, _3451_, _3452_, _3453_, _3454_, _3455_, _3456_, _3457_, _3458_, _3459_, _3460_, _3461_, _3462_, _3463_, _3464_, _3465_, _3466_, _3467_, _3468_, _3469_, _3470_, _3471_, _3472_, _3473_, _3474_, _3475_, _3476_, _3477_, _3478_, _3479_, _3480_, _3481_, _3482_, _3483_, _3484_, _3485_, _3486_, _3487_, _3488_, _3489_, _3490_, _3491_, _3492_, _3493_, _3494_, _3495_, _3496_, _3497_, _3498_, _3499_, _3500_, _3501_, _3502_, _3503_, _3504_, _3505_, _3506_, _3507_, _3508_, _3509_, _3510_, _3511_, _3512_, _3513_, _3514_, _3515_, _3516_, _3517_, _3518_, _3519_, _3520_, _3521_, _3522_, _3523_, _3524_, _3525_, _3526_, _3527_, _3528_, _3529_, _3530_, _3531_, _3532_, _3533_, _3534_, _3535_, _3536_, _3537_, _3538_, _3539_, _3540_, _3541_, _3542_, _3543_, _3544_, _3545_, _3546_, _3547_, _3548_, _3549_, _3550_, _3551_, _3552_, _3553_, _3554_, _3555_, _3556_, _3557_, _3558_, _3559_, _3560_, _3561_, _3562_, _3563_, _3564_, _3565_, _3566_, _3567_, _3568_, _3569_, _3570_, _3571_, _3572_, _3573_, _3574_, _3575_, _3576_, _3577_, _3578_, _3579_, _3580_, _3581_, _3582_, _3583_, _3584_, _3585_, _3586_, _3587_, _3588_, _3589_, _3590_, _3591_, _3592_, _3593_, _3594_, _3595_, _3596_, _3597_, _3598_, _3599_, _3600_, _3601_, _3602_, _3603_, _3604_, _3605_, _3606_, _3607_, _3608_, _3609_, _3610_, _3611_, _3612_, _3613_, _3614_, _3615_, _3616_, _3617_, _3618_, _3619_, _3620_, _3621_, _3622_, _3623_, _3624_, _3625_, _3626_, _3627_, _3628_, _3629_, _3630_, _3631_, _3632_, _3633_, _3634_, _3635_, _3636_, _3637_, _3638_, _3639_, _3640_, _3641_, _3642_, _3643_, _3644_, _3645_, _3646_, _3647_, _3648_, _3649_, _3650_, _3651_, _3652_, _3653_, _3654_, _3655_, _3656_, _3657_, _3658_, _3659_, _3660_, _3661_, _3662_, _3663_, _3664_, _3665_, _3666_, _3667_, _3668_, _3669_, _3670_, _3671_, _3672_, _3673_, _3674_, _3675_, _3676_, _3677_, _3678_, _3679_, _3680_, _3681_, _3682_, _3683_, _3684_, _3685_, _3686_, _3687_, _3688_, _3689_, _3690_, _3691_, _3692_, _3693_, _3694_, _3695_, _3696_, _3697_, _3698_, _3699_, _3700_, _3701_, _3702_, _3703_, _3704_, _3705_, _3706_, _3707_, _3708_, _3709_, _3710_, _3711_, _3712_, _3713_, _3714_, _3715_, _3716_, _3717_, _3718_, _3719_, _3720_, _3721_, _3722_, _3723_, _3724_, _3725_, _3726_, _3727_, _3728_, _3729_, _3730_, _3731_, _3732_, _3733_, _3734_, _3735_, _3736_, _3737_, _3738_, _3739_, _3740_, _3741_, _3742_, _3743_, _3744_, _3745_, _3746_, _3747_, _3748_, _3749_, _3750_, _3751_, _3752_, _3753_, _3754_, _3755_, _3756_, _3757_, _3758_, _3759_, _3760_, _3761_, _3762_, _3763_, _3764_, _3765_, _3766_, _3767_, _3768_, _3769_, _3770_, _3771_, _3772_, _3773_, _3774_, _3775_, _3776_, _3777_, _3778_, _3779_, _3780_, _3781_, _3782_, _3783_, _3784_, _3785_, _3786_, _3787_, _3788_, _3789_, _3790_, _3791_, _3792_, _3793_, _3794_, _3795_, _3796_, _3797_, _3798_, _3799_, _3800_, _3801_, _3802_, _3803_, _3804_, _3805_, _3806_, _3807_, _3808_, _3809_, _3810_, _3811_, _3812_, _3813_, _3814_, _3815_, _3816_, _3817_, _3818_, _3819_, _3820_, _3821_, _3822_, _3823_, _3824_, _3825_, _3826_, _3827_, _3828_, _3829_, _3830_, _3831_, _3832_, _3833_, _3834_, _3835_, _3836_, _3837_, _3838_, _3839_, _3840_, _3841_, _3842_, _3843_, _3844_, _3845_, _3846_, _3847_, _3848_, _3849_, _3850_, _3851_, _3852_, _3853_, _3854_, _3855_, _3856_, _3857_, _3858_, _3859_, _3860_, _3861_, _3862_, _3863_, _3864_, _3865_, _3866_, _3867_, _3868_, _3869_, _3870_, _3871_, _3872_, _3873_, _3874_, _3875_, _3876_, _3877_, _3878_, _3879_, _3880_, _3881_, _3882_, _3883_, _3884_, _3885_, _3886_, _3887_, _3888_, _3889_, _3890_, _3891_, _3892_, _3893_, _3894_, _3895_, _3896_, _3897_, _3898_, _3899_, _3900_, _3901_, _3902_, _3903_, _3904_, _3905_, _3906_, _3907_, _3908_, _3909_, _3910_, _3911_, _3912_, _3913_, _3914_, _3915_, _3916_, _3917_, _3918_, _3919_, _3920_, _3921_, _3922_, _3923_, _3924_, _3925_, _3926_, _3927_, _3928_, _3929_, _3930_, _3931_, _3932_, _3933_, _3934_, _3935_, _3936_, _3937_, _3938_, _3939_, _3940_, _3941_, _3942_, _3943_, _3944_, _3945_, _3946_, _3947_, _3948_, _3949_, _3950_, _3951_, _3952_, _3953_, _3954_, _3955_, _3956_, _3957_, _3958_, _3959_, _3960_, _3961_, _3962_, _3963_, _3964_, _3965_, _3966_, _3967_, _3968_, _3969_, _3970_, _3971_, _3972_, _3973_, _3974_, _3975_, _3976_, _3977_, _3978_, _3979_, _3980_, _3981_, _3982_, _3983_, _3984_, _3985_, _3986_, _3987_, _3988_, _3989_, _3990_, _3991_, _3992_, _3993_, _3994_, _3995_, _3996_, _3997_, _3998_, _3999_, _4000_, _4001_, _4002_, _4003_, _4004_, _4005_, _4006_, _4007_, _4008_, _4009_, _4010_, _4011_, _4012_, _4013_, _4014_, _4015_, _4016_, _4017_, _4018_, _4019_, _4020_, _4021_, _4022_, _4023_, _4024_, _4025_, _4026_, _4027_, _4028_, _4029_, _4030_, _4031_, _4032_, _4033_, _4034_, _4035_, _4036_, _4037_, _4038_, _4039_, _4040_, _4041_, _4042_, _4043_, _4044_, _4045_, _4046_, _4047_, _4048_, _4049_, _4050_, _4051_, _4052_, _4053_, _4054_, _4055_, _4056_, _4057_, _4058_, _4059_, _4060_, _4061_, _4062_, _4063_, _4064_, _4065_, _4066_, _4067_, _4068_, _4069_, _4070_, _4071_, _4072_, _4073_, _4074_, _4075_, _4076_, _4077_, _4078_, _4079_, _4080_, _4081_, _4082_, _4083_, _4084_, _4085_, _4086_, _4087_, _4088_, _4089_, _4090_, _4091_, _4092_, _4093_, _4094_, _4095_, _4096_, _4097_, _4098_, _4099_, _4100_, _4101_, _4102_, _4103_, _4104_, _4105_, _4106_, _4107_, _4108_, _4109_, _4110_, _4111_, _4112_, _4113_, _4114_, _4115_, _4116_, _4117_, _4118_, _4119_, _4120_, _4121_, _4122_, _4123_, _4124_, _4125_, _4126_, _4127_, _4128_, _4129_, _4130_, _4131_, _4132_, _4133_, _4134_, _4135_, _4136_, _4137_, _4138_, _4139_, _4140_, _4141_, _4142_, _4143_, _4144_, _4145_, _4146_, _4147_, _4148_, _4149_, _4150_, _4151_, _4152_, _4153_, _4154_, _4155_, _4156_, _4157_, _4158_, _4159_, _4160_, _4161_, _4162_, _4163_, _4164_, _4165_, _4166_, _4167_, _4168_, _4169_, _4170_, _4171_, _4172_, _4173_, _4174_, _4175_, _4176_, _4177_, _4178_, _4179_, _4180_, _4181_, _4182_, _4183_, _4184_, _4185_, _4186_, _4187_, _4188_, _4189_, _4190_, _4191_, _4192_, _4193_, _4194_, _4195_, _4196_, _4197_, _4198_, _4199_, _4200_, _4201_, _4202_, _4203_, _4204_, _4205_, _4206_, _4207_, _4208_, _4209_, _4210_, _4211_, _4212_, _4213_, _4214_, _4215_, _4216_, _4217_, _4218_, _4219_, _4220_, _4221_, _4222_, _4223_, _4224_, _4225_, _4226_, _4227_, _4228_, _4229_, _4230_, _4231_, _4232_, _4233_, _4234_, _4235_, _4236_, _4237_, _4238_, _4239_, _4240_, _4241_, _4242_, _4243_, _4244_, _4245_, _4246_, _4247_, _4248_, _4249_, _4250_, _4251_, _4252_, _4253_, _4254_, _4255_, _4256_, _4257_, _4258_, _4259_, _4260_, _4261_, _4262_, _4263_, _4264_, _4265_, _4266_, _4267_, _4268_, _4269_, _4270_, _4271_, _4272_, _4273_, _4274_, _4275_, _4276_, _4277_, _4278_, _4279_, _4280_, _4281_, _4282_, _4283_, _4284_, _4285_, _4286_, _4287_, _4288_, _4289_, _4290_, _4291_, _4292_, _4293_, _4294_, _4295_, _4296_, _4297_, _4298_, _4299_, _4300_, _4301_, _4302_, _4303_, _4304_, _4305_, _4306_, _4307_, _4308_, _4309_, _4310_, _4311_, _4312_, _4313_, _4314_, _4315_, _4316_, _4317_, _4318_, _4319_, _4320_, _4321_, _4322_, _4323_, _4324_, _4325_, _4326_, _4327_, _4328_, _4329_, _4330_, _4331_, _4332_, _4333_, _4334_, _4335_, _4336_, _4337_, _4338_, _4339_, _4340_, _4341_, _4342_, _4343_, _4344_, _4345_, _4346_, _4347_, _4348_, _4349_, _4350_, _4351_, _4352_, _4353_, _4354_, _4355_, _4356_, _4357_, _4358_, _4359_, _4360_, _4361_, _4362_, _4363_, _4364_, _4365_, _4366_, _4367_, _4368_, _4369_, _4370_, _4371_, _4372_, _4373_, _4374_, _4375_, _4376_, _4377_, _4378_, _4379_, _4380_, _4381_, _4382_, _4383_, _4384_, _4385_, _4386_, _4387_, _4388_, _4389_, _4390_, _4391_, _4392_, _4393_, _4394_, _4395_, _4396_, _4397_, _4398_, _4399_, _4400_, _4401_, _4402_, _4403_, _4404_, _4405_, _4406_, _4407_, _4408_, _4409_, _4410_, _4411_, _4412_, _4413_, _4414_, _4415_, _4416_, _4417_, _4418_, _4419_, _4420_, _4421_, _4422_, _4423_, _4424_, _4425_, _4426_, _4427_, _4428_, _4429_, _4430_, _4431_, _4432_, _4433_, _4434_, _4435_, _4436_, _4437_, _4438_, _4439_, _4440_, _4441_, _4442_, _4443_, _4444_, _4445_, _4446_, _4447_, _4448_, _4449_, _4450_, _4451_, _4452_, _4453_, _4454_, _4455_, _4456_, _4457_, _4458_, _4459_, _4460_, _4461_, _4462_, _4463_, _4464_, _4465_, _4466_, _4467_, _4468_, _4469_, _4470_, _4471_, _4472_, _4473_, _4474_, _4475_, _4476_, _4477_, _4478_, _4479_, _4480_, _4481_, _4482_, _4483_, _4484_, _4485_, _4486_, _4487_, _4488_, _4489_, _4490_, _4491_, _4492_, _4493_, _4494_, _4495_, _4496_, _4497_, _4498_, _4499_, _4500_, _4501_, _4502_, _4503_, _4504_, _4505_, _4506_, _4507_, _4508_, _4509_, _4510_, _4511_, _4512_, _4513_, _4514_, _4515_, _4516_, _4517_, _4518_, _4519_, _4520_, _4521_, _4522_, _4523_, _4524_, _4525_, _4526_, _4527_, _4528_, _4529_, _4530_, _4531_, _4532_, _4533_, _4534_, _4535_, _4536_, _4537_, _4538_, _4539_, _4540_, _4541_, _4542_, _4543_, _4544_, _4545_, _4546_, _4547_, _4548_, _4549_, _4550_, _4551_, _4552_, _4553_, _4554_, _4555_, _4556_, _4557_, _4558_, _4559_, _4560_, _4561_, _4562_, _4563_, _4564_, _4565_, _4566_, _4567_, _4568_, _4569_, _4570_, _4571_, _4572_, _4573_, _4574_, _4575_, _4576_, _4577_, _4578_, _4579_, _4580_, _4581_, _4582_, _4583_, _4584_, _4585_, _4586_, _4587_, _4588_, _4589_, _4590_, _4591_, _4592_, _4593_, _4594_, _4595_, _4596_, _4597_, _4598_, _4599_, _4600_, _4601_, _4602_, _4603_, _4604_, _4605_, _4606_, _4607_, _4608_, _4609_, _4610_, _4611_, _4612_, _4613_, _4614_, _4615_, _4616_, _4617_, _4618_, _4619_, _4620_, _4621_, _4622_, _4623_, _4624_, _4625_, _4626_, _4627_, _4628_, _4629_, _4630_, _4631_, _4632_, _4633_, _4634_, _4635_, _4636_, _4637_, _4638_, _4639_, _4640_, _4641_, _4642_, _4643_, _4644_, _4645_, _4646_, _4647_, _4648_, _4649_, _4650_, _4651_, _4652_, _4653_, _4654_, _4655_, _4656_, _4657_, _4658_, _4659_, _4660_, _4661_, _4662_, _4663_, _4664_, _4665_, _4666_, _4667_, _4668_, _4669_, _4670_, _4671_, _4672_, _4673_, _4674_, _4675_, _4676_, _4677_, _4678_, _4679_, _4680_, _4681_, _4682_, _4683_, _4684_, _4685_, _4686_, _4687_, _4688_, _4689_, _4690_, _4691_, _4692_, _4693_, _4694_, _4695_, _4696_, _4697_, _4698_, _4699_, _4700_, _4701_, _4702_, _4703_, _4704_, _4705_, _4706_, _4707_, _4708_, _4709_, _4710_, _4711_, _4712_, _4713_, _4714_, _4715_, _4716_, _4717_, _4718_, _4719_, _4720_, _4721_, _4722_, _4723_, _4724_, _4725_, _4726_, _4727_, _4728_, _4729_, _4730_, _4731_, _4732_, _4733_, _4734_, _4735_, _4736_, _4737_, _4738_, _4739_, _4740_, _4741_, _4742_, _4743_, _4744_, _4745_, _4746_, _4747_, _4748_, _4749_, _4750_, _4751_, _4752_, _4753_, _4754_, _4755_, _4756_, _4757_, _4758_, _4759_, _4760_, _4761_, _4762_, _4763_, _4764_, _4765_, _4766_, _4767_, _4768_, _4769_, _4770_, _4771_, _4772_, _4773_, _4774_, _4775_, _4776_, _4777_, _4778_, _4779_, _4780_, _4781_, _4782_, _4783_, _4784_, _4785_, _4786_, _4787_, _4788_, _4789_, _4790_, _4791_, _4792_, _4793_, _4794_, _4795_, _4796_, _4797_, _4798_, _4799_, _4800_, _4801_, _4802_, _4803_, _4804_, _4805_, _4806_, _4807_, _4808_, _4809_, _4810_, _4811_, _4812_, _4813_, _4814_, _4815_, _4816_, _4817_, _4818_, _4819_, _4820_, _4821_, _4822_, _4823_, _4824_, _4825_, _4826_, _4827_, _4828_, _4829_, _4830_, _4831_, _4832_, _4833_, _4834_, _4835_, _4836_, _4837_, _4838_, _4839_, _4840_, _4841_, _4842_, _4843_, _4844_, _4845_, _4846_, _4847_, _4848_, _4849_, _4850_, _4851_, _4852_, _4853_, _4854_, _4855_, _4856_, _4857_, _4858_, _4859_, _4860_, _4861_, _4862_, _4863_, _4864_, _4865_, _4866_, _4867_, _4868_, _4869_, _4870_, _4871_, _4872_, _4873_, _4874_, _4875_, _4876_, _4877_, _4878_, _4879_, _4880_, _4881_, _4882_, _4883_, _4884_, _4885_, _4886_, _4887_, _4888_, _4889_, _4890_, _4891_, _4892_, _4893_, _4894_, _4895_, _4896_, _4897_, _4898_, _4899_, _4900_, _4901_, _4902_, _4903_, _4904_, _4905_, _4906_, _4907_, _4908_, _4909_, _4910_, _4911_, _4912_, _4913_, _4914_, _4915_, _4916_, _4917_, _4918_, _4919_, _4920_, _4921_, _4922_, _4923_, _4924_, _4925_, _4926_, _4927_, _4928_, _4929_, _4930_, _4931_, _4932_, _4933_, _4934_, _4935_, _4936_, _4937_, _4938_, _4939_, _4940_, _4941_, _4942_, _4943_, _4944_, _4945_, _4946_, _4947_, _4948_, _4949_, _4950_, _4951_, _4952_, _4953_, _4954_, _4955_, _4956_, _4957_, _4958_, _4959_, _4960_, _4961_, _4962_, _4963_, _4964_, _4965_, _4966_, _4967_, _4968_, _4969_, _4970_, _4971_, _4972_, _4973_, _4974_, _4975_, _4976_, _4977_, _4978_, _4979_, _4980_, _4981_, _4982_, _4983_, _4984_, _4985_, _4986_, _4987_, _4988_, _4989_, _4990_, _4991_, _4992_, _4993_, _4994_, _4995_, _4996_, _4997_, _4998_, _4999_, _5000_, _5001_, _5002_, _5003_, _5004_, _5005_, _5006_, _5007_, _5008_, _5009_, _5010_, _5011_, _5012_, _5013_, _5014_, _5015_, _5016_, _5017_, _5018_, _5019_, _5020_, _5021_, _5022_, _5023_, _5024_, _5025_, _5026_, _5027_, _5028_, _5029_, _5030_, _5031_, _5032_, _5033_, _5034_, _5035_, _5036_, _5037_, _5038_, _5039_, _5040_, _5041_, _5042_, _5043_, _5044_, _5045_, _5046_, _5047_, _5048_, _5049_, _5050_, _5051_, _5052_, _5053_, _5054_, _5055_, _5056_, _5057_, _5058_, _5059_, _5060_, _5061_, _5062_, _5063_, _5064_, _5065_, _5066_, _5067_, _5068_, _5069_, _5070_, _5071_, _5072_, _5073_, _5074_, _5075_, _5076_, _5077_, _5078_, _5079_, _5080_, _5081_, _5082_, _5083_, _5084_, _5085_, _5086_, _5087_, _5088_, _5089_, _5090_, _5091_, _5092_, _5093_, _5094_, _5095_, _5096_, _5097_, _5098_, _5099_, _5100_, _5101_, _5102_, _5103_, _5104_, _5105_, _5106_, _5107_, _5108_, _5109_, _5110_, _5111_, _5112_, _5113_, _5114_, _5115_, _5116_, _5117_, _5118_, _5119_, _5120_, _5121_, _5122_, _5123_, _5124_, _5125_, _5126_, _5127_, _5128_, _5129_, _5130_, _5131_, _5132_, _5133_, _5134_, _5135_, _5136_, _5137_, _5138_, _5139_, _5140_, _5141_, _5142_, _5143_, _5144_, _5145_, _5146_, _5147_, _5148_, _5149_, _5150_, _5151_, _5152_, _5153_, _5154_, _5155_, _5156_, _5157_, _5158_, _5159_, _5160_, _5161_, _5162_, _5163_, _5164_, _5165_, _5166_, _5167_, _5168_, _5169_, _5170_, _5171_, _5172_, _5173_, _5174_, _5175_, _5176_, _5177_, _5178_, _5179_, _5180_, _5181_, _5182_, _5183_, _5184_, _5185_, _5186_, _5187_, _5188_, _5189_, _5190_, _5191_, _5192_, _5193_, _5194_, _5195_, _5196_, _5197_, _5198_, _5199_, _5200_, _5201_, _5202_, _5203_, _5204_, _5205_, _5206_, _5207_, _5208_, _5209_, _5210_, _5211_, _5212_, _5213_, _5214_, _5215_, _5216_, _5217_, _5218_, _5219_, _5220_, _5221_, _5222_, _5223_, _5224_, _5225_, _5226_, _5227_, _5228_, _5229_, _5230_, _5231_, _5232_, _5233_, _5234_, _5235_, _5236_, _5237_, _5238_, _5239_, _5240_, _5241_, _5242_, _5243_, _5244_, _5245_, _5246_, _5247_, _5248_, _5249_, _5250_, _5251_, _5252_, _5253_, _5254_, _5255_, _5256_, _5257_, _5258_, _5259_, _5260_, _5261_, _5262_, _5263_, _5264_, _5265_, _5266_, _5267_, _5268_, _5269_, _5270_, _5271_, _5272_, _5273_, _5274_, _5275_, _5276_, _5277_, _5278_, _5279_, _5280_, _5281_, _5282_, _5283_, _5284_, _5285_, _5286_, _5287_, _5288_, _5289_, _5290_, _5291_, _5292_, _5293_, _5294_, _5295_, _5296_, _5297_, _5298_, _5299_, _5300_, _5301_, _5302_, _5303_, _5304_, _5305_, _5306_, _5307_, _5308_, _5309_, _5310_, _5311_, _5312_, _5313_, _5314_, _5315_, _5316_, _5317_, _5318_, _5319_, _5320_, _5321_, _5322_, _5323_, _5324_, _5325_, _5326_, _5327_, _5328_, _5329_, _5330_, _5331_, _5332_, _5333_, _5334_, _5335_, _5336_, _5337_, _5338_, _5339_, _5340_, _5341_, _5342_, _5343_, _5344_, _5345_, _5346_, _5347_, _5348_, _5349_, _5350_, _5351_, _5352_, _5353_, _5354_, _5355_, _5356_, _5357_, _5358_, _5359_, _5360_, _5361_, _5362_, _5363_, _5364_, _5365_, _5366_, _5367_, _5368_, _5369_, _5370_, _5371_, _5372_, _5373_, _5374_, _5375_, _5376_, _5377_, _5378_, _5379_, _5380_, _5381_, _5382_, _5383_, _5384_, _5385_, _5386_, _5387_, _5388_, _5389_, _5390_, _5391_, _5392_, _5393_, _5394_, _5395_, _5396_, _5397_, _5398_, _5399_, _5400_, _5401_, _5402_, _5403_, _5404_, _5405_, _5406_, _5407_, _5408_, _5409_, _5410_, _5411_, _5412_, _5413_, _5414_, _5415_, _5416_, _5417_, _5418_, _5419_, _5420_, _5421_, _5422_, _5423_, _5424_, _5425_, _5426_, _5427_, _5428_, _5429_, _5430_, _5431_, _5432_, _5433_, _5434_, _5435_, _5436_, _5437_, _5438_, _5439_, _5440_, _5441_, _5442_, _5443_, _5444_, _5445_, _5446_, _5447_, _5448_, _5449_, _5450_, _5451_, _5452_, _5453_, _5454_, _5455_, _5456_, _5457_, _5458_, _5459_, _5460_, _5461_, _5462_, _5463_, _5464_, _5465_, _5466_, _5467_, _5468_, _5469_, _5470_, _5471_, _5472_, _5473_, _5474_, _5475_, _5476_, _5477_, _5478_, _5479_, _5480_, _5481_, _5482_, _5483_, _5484_, _5485_, _5486_, _5487_, _5488_, _5489_, _5490_, _5491_, _5492_, _5493_, _5494_, _5495_, _5496_, _5497_, _5498_, _5499_, _5500_, _5501_, _5502_, _5503_, _5504_, _5505_, _5506_, _5507_, _5508_, _5509_, _5510_, _5511_, _5512_, _5513_, _5514_, _5515_, _5516_, _5517_, _5518_, _5519_, _5520_, _5521_, _5522_, _5523_, _5524_, _5525_, _5526_, _5527_, _5528_, _5529_, _5530_, _5531_, _5532_, _5533_, _5534_, _5535_, _5536_, _5537_, _5538_, _5539_, _5540_, _5541_, _5542_, _5543_, _5544_, _5545_, _5546_, _5547_, _5548_, _5549_, _5550_, _5551_, _5552_, _5553_, _5554_, _5555_, _5556_, _5557_, _5558_, _5559_, _5560_, _5561_, _5562_, _5563_, _5564_, _5565_, _5566_, _5567_, _5568_, _5569_, _5570_, _5571_, _5572_, _5573_, _5574_, _5575_, _5576_, _5577_, _5578_, _5579_, _5580_, _5581_, _5582_, _5583_, _5584_, _5585_, _5586_, _5587_, _5588_, _5589_, _5590_, _5591_, _5592_, _5593_, _5594_, _5595_, _5596_, _5597_, _5598_, _5599_, _5600_, _5601_, _5602_, _5603_, _5604_, _5605_, _5606_, _5607_, _5608_, _5609_, _5610_, _5611_, _5612_, _5613_, _5614_, _5615_, _5616_, _5617_, _5618_, _5619_, _5620_, _5621_, _5622_, _5623_, _5624_, _5625_, _5626_, _5627_, _5628_, _5629_, _5630_, _5631_, _5632_, _5633_, _5634_, _5635_, _5636_, _5637_, _5638_, _5639_, _5640_, _5641_, _5642_, _5643_, _5644_, _5645_, _5646_, _5647_, _5648_, _5649_, _5650_, _5651_, _5652_, _5653_, _5654_, _5655_, _5656_, _5657_, _5658_, _5659_, _5660_, _5661_, _5662_, _5663_, _5664_, _5665_, _5666_, _5667_, _5668_, _5669_, _5670_, _5671_, _5672_, _5673_, _5674_, _5675_, _5676_, _5677_, _5678_, _5679_, _5680_, _5681_, _5682_, _5683_, _5684_, _5685_, _5686_, _5687_, _5688_, _5689_, _5690_, _5691_, _5692_, _5693_, _5694_, _5695_, _5696_, _5697_, _5698_, _5699_, _5700_, _5701_, _5702_, _5703_, _5704_, _5705_, _5706_, _5707_, _5708_, _5709_, _5710_, _5711_, _5712_, _5713_, _5714_, _5715_, _5716_, _5717_, _5718_, _5719_, _5720_, _5721_, _5722_, _5723_, _5724_, _5725_, _5726_, _5727_, _5728_, _5729_, _5730_, _5731_, _5732_, _5733_, _5734_, _5735_, _5736_, _5737_, _5738_, _5739_, _5740_, _5741_, _5742_, _5743_, _5744_, _5745_, _5746_, _5747_, _5748_, _5749_, _5750_, _5751_, _5752_, _5753_, _5754_, _5755_, _5756_, _5757_, _5758_, _5759_, _5760_, _5761_, _5762_, _5763_, _5764_, _5765_, _5766_, _5767_, _5768_, _5769_, _5770_, _5771_, _5772_, _5773_, _5774_, _5775_, _5776_, _5777_, _5778_, _5779_, _5780_, _5781_, _5782_, _5783_, _5784_, _5785_, _5786_, _5787_, _5788_, _5789_, _5790_, _5791_, _5792_, _5793_, _5794_, _5795_, _5796_, _5797_, _5798_, _5799_, _5800_, _5801_, _5802_, _5803_, _5804_, _5805_, _5806_, _5807_, _5808_, _5809_, _5810_, _5811_, _5812_, _5813_, _5814_, _5815_, _5816_, _5817_, _5818_;
  input [31:0] G11;
  input [31:0] G12;
  input G11[0], G11[1], G11[2], G11[3], G11[4], G11[5], G11[6], G11[7], G11[8], G11[9], G11[10], G11[11], G11[12], G11[13], G11[14], G11[15], G11[16], G11[17], G11[18], G11[19], G11[20], G11[21], G11[22], G11[23], G11[24], G11[25], G11[26], G11[27], G11[28], G11[29], G11[30], G11[31], G12[0], G12[1], G12[2], G12[3], G12[4], G12[5], G12[6], G12[7], G12[8], G12[9], G12[10], G12[11], G12[12], G12[13], G12[14], G12[15], G12[16], G12[17], G12[18], G12[19], G12[20], G12[21], G12[22], G12[23], G12[24], G12[25], G12[26], G12[27], G12[28], G12[29], G12[30], G12[31];
  output G14[0], G14[1], G14[2], G14[3], G14[4], G14[5], G14[6], G14[7], G14[8], G14[9], G14[10], G14[11], G14[12], G14[13], G14[14], G14[15], G14[16], G14[17], G14[18], G14[19], G14[20], G14[21], G14[22], G14[23], G14[24], G14[25], G14[26], G14[27], G14[28], G14[29], G14[30], G14[31];
  and g_5819_(_5433_, _5517_, _5519_);
  xor g_5820_(_5433_, _5517_, _5520_);
  and g_5821_(_5516_, _5520_, _5521_);
  xor g_5822_(_5516_, _5520_, _5522_);
  or g_5823_(_5447_, _5449_, _5523_);
  and g_5824_(_5522_, _5523_, _5524_);
  xor g_5825_(_5522_, _5523_, _5525_);
  and g_5826_(_5515_, _5525_, _5526_);
  xor g_5827_(_5515_, _5525_, _5527_);
  or g_5828_(_5459_, _5461_, _5528_);
  and g_5829_(G12[5], G11[9], _5529_);
  and g_5830_(G12[2], G11[12], _5530_);
  and g_5831_(G12[4], G11[12], _5531_);
  and g_5832_(_5364_, _5530_, _5532_);
  xor g_5833_(_5364_, _5530_, _5533_);
  and g_5834_(_5529_, _5533_, _5534_);
  xor g_5835_(_5529_, _5533_, _5535_);
  or g_5836_(_5455_, _5457_, _5536_);
  and g_5837_(G12[1], G11[13], _5537_);
  and g_5838_(G12[0], G11[14], _5538_);
  and g_5839_(G12[3], G11[14], _5539_);
  and g_5840_(_5295_, _5538_, _5540_);
  xor g_5841_(_5295_, _5538_, _5541_);
  and g_5842_(_5537_, _5541_, _5542_);
  xor g_5843_(_5537_, _5541_, _5543_);
  and g_5844_(_5536_, _5543_, _5544_);
  xor g_5845_(_5536_, _5543_, _5545_);
  and g_5846_(_5535_, _5545_, _5546_);
  xor g_5847_(_5535_, _5545_, _5547_);
  and g_5848_(_5528_, _5547_, _5548_);
  xor g_5849_(_5528_, _5547_, _5549_);
  and g_5850_(_5527_, _5549_, _5550_);
  xor g_5851_(_5527_, _5549_, _5551_);
  and g_5852_(_5514_, _5551_, _5552_);
  xor g_5853_(_5514_, _5551_, _5553_);
  and g_5854_(_5513_, _5553_, _5554_);
  xor g_5855_(_5513_, _5553_, _5555_);
  and g_5856_(_5488_, _5555_, _5556_);
  xor g_5857_(_5488_, _5555_, _5557_);
  and g_5858_(_5487_, _5557_, _5558_);
  xor g_5859_(_5487_, _5557_, _5559_);
  and g_5860_(_5484_, _5559_, _5560_);
  xor g_5861_(_5484_, _5559_, _5561_);
  and g_5862_(_5475_, _5561_, _5562_);
  xor g_5863_(_5475_, _5561_, _5563_);
  and g_5864_(_5395_, _5478_, _5564_);
  or g_5865_(_5477_, _5564_, _5565_);
  and g_5866_(_5563_, _5564_, _5566_);
  and g_5867_(_5477_, _5563_, _5567_);
  xor g_5868_(_5563_, _5565_, _5568_);
  and g_5869_(_5483_, _5568_, _5569_);
  xor g_5870_(_5483_, _5568_, G14[14]);
  or g_5871_(_5566_, _5569_, _5570_);
  or g_5872_(_5556_, _5558_, _5571_);
  and g_5873_(G11[0], G12[15], _5572_);
  or g_5874_(_5493_, _5495_, _5573_);
  and g_5875_(_5572_, _5573_, _5574_);
  xor g_5876_(_5572_, _5573_, _5575_);
  or g_5877_(_5510_, _5512_, _5576_);
  and g_5878_(_5575_, _5576_, _5577_);
  xor g_5879_(_5575_, _5576_, _5578_);
  or g_5880_(_5552_, _5554_, _5579_);
  or g_5881_(_5505_, _5507_, _5580_);
  and g_5882_(G11[1], G12[14], _5581_);
  and g_5883_(G11[3], G12[12], _5582_);
  and g_5884_(G11[3], G12[13], _5583_);
  and g_5885_(_5492_, _5582_, _5584_);
  xor g_5886_(_5492_, _5582_, _5585_);
  and g_5887_(_5581_, _5585_, _5586_);
  xor g_5888_(_5581_, _5585_, _5587_);
  or g_5889_(_5501_, _5503_, _5588_);
  and g_5890_(G11[4], G12[11], _5589_);
  and g_5891_(G11[6], G12[9], _5590_);
  and g_5892_(G11[6], G12[10], _5591_);
  and g_5893_(_5500_, _5590_, _5592_);
  xor g_5894_(_5500_, _5590_, _5593_);
  and g_5895_(_5589_, _5593_, _5594_);
  xor g_5896_(_5589_, _5593_, _5595_);
  and g_5897_(_5588_, _5595_, _5596_);
  xor g_5898_(_5588_, _5595_, _5597_);
  and g_5899_(_5587_, _5597_, _5598_);
  xor g_5900_(_5587_, _5597_, _5599_);
  or g_5901_(_5524_, _5526_, _5600_);
  and g_5902_(_5599_, _5600_, _5601_);
  xor g_5903_(_5599_, _5600_, _5602_);
  and g_5904_(_5580_, _5602_, _5603_);
  xor g_5905_(_5580_, _5602_, _5604_);
  or g_5906_(_5548_, _5550_, _5605_);
  or g_5907_(_5519_, _5521_, _5606_);
  and g_5908_(G11[7], G12[8], _5607_);
  and g_5909_(G12[6], G11[9], _5608_);
  and g_5910_(G12[7], G11[9], _5609_);
  and g_5911_(_5518_, _5608_, _5610_);
  xor g_5912_(_5518_, _5608_, _5611_);
  and g_5913_(_5607_, _5611_, _5612_);
  xor g_5914_(_5607_, _5611_, _5613_);
  or g_5915_(_5532_, _5534_, _5614_);
  and g_5916_(_5613_, _5614_, _5615_);
  xor g_5917_(_5613_, _5614_, _5616_);
  and g_5918_(_5606_, _5616_, _5617_);
  xor g_5919_(_5606_, _5616_, _5618_);
  or g_5920_(_5544_, _5546_, _5619_);
  and g_5921_(G12[5], G11[10], _5620_);
  and g_5922_(G12[2], G11[13], _5621_);
  and g_5923_(G12[4], G11[13], _5622_);
  and g_5924_(_5446_, _5621_, _5623_);
  xor g_5925_(_5446_, _5621_, _5624_);
  and g_5926_(_5620_, _5624_, _5625_);
  xor g_5927_(_5620_, _5624_, _5626_);
  or g_5928_(_5540_, _5542_, _5627_);
  and g_5929_(G12[1], G11[14], _5628_);
  and g_5930_(G12[0], G11[15], _5629_);
  and g_5931_(G12[3], G11[15], _5630_);
  and g_5932_(_5372_, _5629_, _5631_);
  xor g_5933_(_5372_, _5629_, _5632_);
  and g_5934_(_5628_, _5632_, _5633_);
  xor g_5935_(_5628_, _5632_, _5634_);
  and g_5936_(_5627_, _5634_, _5635_);
  xor g_5937_(_5627_, _5634_, _5636_);
  and g_5938_(_5626_, _5636_, _5637_);
  xor g_5939_(_5626_, _5636_, _5638_);
  and g_5940_(_5619_, _5638_, _5639_);
  xor g_5941_(_5619_, _5638_, _5640_);
  and g_5942_(_5618_, _5640_, _5641_);
  xor g_5943_(_5618_, _5640_, _5642_);
  and g_5944_(_5605_, _5642_, _5643_);
  xor g_5945_(_5605_, _5642_, _5644_);
  and g_5946_(_5604_, _5644_, _5645_);
  xor g_5947_(_5604_, _5644_, _5646_);
  and g_5948_(_5579_, _5646_, _5647_);
  xor g_5949_(_5579_, _5646_, _5648_);
  and g_5950_(_5578_, _5648_, _5649_);
  xor g_5951_(_5578_, _5648_, _5650_);
  and g_5952_(_5571_, _5650_, _5651_);
  xor g_5953_(_5571_, _5650_, _5652_);
  and g_5954_(_5486_, _5652_, _5653_);
  xor g_5955_(_5486_, _5652_, _5654_);
  and g_5956_(_5560_, _5654_, _5655_);
  xor g_5957_(_5560_, _5654_, _5656_);
  or g_5958_(_5562_, _5567_, _5657_);
  xor g_5959_(_5656_, _5657_, _5658_);
  and g_5960_(_5570_, _5658_, _5659_);
  xor g_5961_(_5570_, _5658_, G14[15]);
  and g_5962_(_5567_, _5656_, _5660_);
  or g_5963_(_5659_, _5660_, _5661_);
  and g_5964_(_5562_, _5656_, _5662_);
  or g_5965_(_5651_, _5653_, _5663_);
  or g_5966_(_5647_, _5649_, _5664_);
  and g_5967_(G11[0], G12[16], _5665_);
  and g_5968_(G11[1], G12[15], _5666_);
  and g_5969_(G11[1], G12[16], _5667_);
  and g_5970_(_5572_, _5667_, _5668_);
  xor g_5971_(_5665_, _5666_, _5669_);
  or g_5972_(_5584_, _5586_, _5670_);
  and g_5973_(_5669_, _5670_, _5671_);
  xor g_5974_(_5669_, _5670_, _5672_);
  and g_5975_(_5574_, _5672_, _5673_);
  xor g_5976_(_5574_, _5672_, _5674_);
  or g_5977_(_5601_, _5603_, _5675_);
  and g_5978_(_5674_, _5675_, _5676_);
  xor g_5979_(_5674_, _5675_, _5677_);
  or g_5980_(_5643_, _5645_, _5678_);
  or g_5981_(_5596_, _5598_, _5679_);
  and g_5982_(G11[2], G12[14], _5680_);
  and g_5983_(G11[4], G12[12], _5681_);
  and g_5984_(G11[4], G12[13], _5682_);
  and g_5985_(_5583_, _5681_, _5683_);
  xor g_5986_(_5583_, _5681_, _5684_);
  and g_5987_(_5680_, _5684_, _5685_);
  xor g_5988_(_5680_, _5684_, _5686_);
  or g_5989_(_5592_, _5594_, _5687_);
  and g_5990_(G11[5], G12[11], _5688_);
  and g_5991_(G11[7], G12[9], _5689_);
  and g_5992_(G11[7], G12[10], _5690_);
  and g_5993_(_5591_, _5689_, _5691_);
  xor g_5994_(_5591_, _5689_, _5692_);
  and g_5995_(_5688_, _5692_, _5693_);
  xor g_5996_(_5688_, _5692_, _5694_);
  and g_5997_(_5687_, _5694_, _5695_);
  xor g_5998_(_5687_, _5694_, _5696_);
  and g_5999_(_5686_, _5696_, _5697_);
  xor g_6000_(_5686_, _5696_, _5698_);
  or g_6001_(_5615_, _5617_, _5699_);
  and g_6002_(_5698_, _5699_, _5700_);
  xor g_6003_(_5698_, _5699_, _5701_);
  and g_6004_(_5679_, _5701_, _5702_);
  xor g_6005_(_5679_, _5701_, _5703_);
  or g_6006_(_5639_, _5641_, _5704_);
  or g_6007_(_5610_, _5612_, _5705_);
  and g_6008_(G11[8], G12[8], _5706_);
  and g_6009_(G12[6], G11[10], _5707_);
  and g_6010_(G12[7], G11[10], _5708_);
  and g_6011_(_5609_, _5707_, _5709_);
  xor g_6012_(_5609_, _5707_, _5710_);
  and g_6013_(_5706_, _5710_, _5711_);
  xor g_6014_(_5706_, _5710_, _5712_);
  or g_6015_(_5623_, _5625_, _5713_);
  and g_6016_(_5712_, _5713_, _5714_);
  xor g_6017_(_5712_, _5713_, _5715_);
  and g_6018_(_5705_, _5715_, _5716_);
  xor g_6019_(_5705_, _5715_, _5717_);
  or g_6020_(_5635_, _5637_, _5718_);
  and g_6021_(G12[5], G11[11], _5719_);
  and g_6022_(G12[2], G11[14], _5720_);
  and g_6023_(G12[4], G11[14], _5721_);
  and g_6024_(_5531_, _5720_, _5722_);
  xor g_6025_(_5531_, _5720_, _5723_);
  and g_6026_(_5719_, _5723_, _5724_);
  xor g_6027_(_5719_, _5723_, _5725_);
  or g_6028_(_5631_, _5633_, _5726_);
  and g_6029_(G12[1], G11[15], _5727_);
  and g_6030_(G12[0], G11[16], _5728_);
  and g_6031_(G12[3], G11[16], _5729_);
  and g_6032_(_5454_, _5728_, _5730_);
  xor g_6033_(_5454_, _5728_, _5731_);
  and g_6034_(_5727_, _5731_, _5732_);
  xor g_6035_(_5727_, _5731_, _5733_);
  and g_6036_(_5726_, _5733_, _5734_);
  xor g_6037_(_5726_, _5733_, _5735_);
  and g_6038_(_5725_, _5735_, _5736_);
  xor g_6039_(_5725_, _5735_, _5737_);
  and g_6040_(_5718_, _5737_, _5738_);
  xor g_6041_(_5718_, _5737_, _5739_);
  and g_6042_(_5717_, _5739_, _5740_);
  xor g_6043_(_5717_, _5739_, _5741_);
  and g_6044_(_5704_, _5741_, _5742_);
  xor g_6045_(_5704_, _5741_, _5743_);
  and g_6046_(_5703_, _5743_, _5744_);
  xor g_6047_(_5703_, _5743_, _5745_);
  and g_6048_(_5678_, _5745_, _5746_);
  xor g_6049_(_5678_, _5745_, _5747_);
  and g_6050_(_5677_, _5747_, _5748_);
  xor g_6051_(_5677_, _5747_, _5749_);
  and g_6052_(_5664_, _5749_, _5750_);
  xor g_6053_(_5664_, _5749_, _5751_);
  and g_6054_(_5577_, _5751_, _5752_);
  xor g_6055_(_5577_, _5751_, _5753_);
  and g_6056_(_5663_, _5753_, _5754_);
  xor g_6057_(_5663_, _5753_, _5755_);
  and g_6058_(_5655_, _5755_, _5756_);
  xor g_6059_(_5655_, _5755_, _5757_);
  and g_6060_(_5662_, _5757_, _5758_);
  xor g_6061_(_5662_, _5757_, _5759_);
  and g_6062_(_5661_, _5759_, _5760_);
  xor g_6063_(_5661_, _5759_, G14[16]);
  or g_6064_(_5758_, _5760_, _5761_);
  or g_6065_(_5750_, _5752_, _5762_);
  or g_6066_(_5746_, _5748_, _5763_);
  or g_6067_(_5700_, _5702_, _5764_);
  and g_6068_(G11[0], G12[17], _5765_);
  and g_6069_(G11[2], G12[15], _5766_);
  and g_6070_(G11[2], G12[16], _5767_);
  and g_6071_(_5667_, _5766_, _5768_);
  xor g_6072_(_5667_, _5766_, _5769_);
  and g_6073_(_5765_, _5769_, _5770_);
  xor g_6074_(_5765_, _5769_, _5771_);
  or g_6075_(_5683_, _5685_, _5772_);
  and g_6076_(_5771_, _5772_, _5773_);
  or g_6077_(_5771_, _5772_, _5774_);
  xor g_6078_(_5771_, _5772_, _5775_);
  or g_6079_(_5668_, _5671_, _5776_);
  xor g_6080_(_5775_, _5776_, _5777_);
  and g_6081_(_5764_, _5777_, _5778_);
  xor g_6082_(_5764_, _5777_, _5779_);
  and g_6083_(_5673_, _5779_, _5780_);
  xor g_6084_(_5673_, _5779_, _5781_);
  or g_6085_(_5742_, _5744_, _5782_);
  or g_6086_(_5695_, _5697_, _5783_);
  and g_6087_(G11[3], G12[14], _5784_);
  and g_6088_(G11[5], G12[12], _5785_);
  and g_6089_(G11[5], G12[13], _5786_);
  and g_6090_(_5682_, _5785_, _5787_);
  xor g_6091_(_5682_, _5785_, _5788_);
  and g_6092_(_5784_, _5788_, _5789_);
  xor g_6093_(_5784_, _5788_, _5790_);
  or g_6094_(_5691_, _5693_, _5791_);
  and g_6095_(G11[6], G12[11], _5792_);
  and g_6096_(G11[8], G12[9], _5793_);
  and g_6097_(G11[8], G12[10], _5794_);
  and g_6098_(_5690_, _5793_, _5795_);
  xor g_6099_(_5690_, _5793_, _5797_);
  and g_6100_(_5792_, _5797_, _5798_);
  xor g_6101_(_5792_, _5797_, _5799_);
  and g_6102_(_5791_, _5799_, _5800_);
  xor g_6103_(_5791_, _5799_, _5801_);
  and g_6104_(_5790_, _5801_, _5802_);
  xor g_6105_(_5790_, _5801_, _5803_);
  or g_6106_(_5714_, _5716_, _5804_);
  and g_6107_(_5803_, _5804_, _5805_);
  xor g_6108_(_5803_, _5804_, _5806_);
  and g_6109_(_5783_, _5806_, _5808_);
  xor g_6110_(_5783_, _5806_, _5809_);
  or g_6111_(_5738_, _5740_, _5810_);
  or g_6112_(_5709_, _5711_, _5811_);
  and g_6113_(G12[8], G11[9], _5812_);
  and g_6114_(G12[6], G11[11], _5813_);
  and g_6115_(G12[7], G11[11], _5814_);
  and g_6116_(_5708_, _5813_, _5815_);
  xor g_6117_(_5708_, _5813_, _5816_);
  and g_6118_(_5812_, _5816_, _5817_);
  xor g_6119_(_5812_, _5816_, _2876_);
  or g_6120_(_5722_, _5724_, _2877_);
  and g_6121_(_2876_, _2877_, _2878_);
  xor g_6122_(_2876_, _2877_, _2879_);
  and g_6123_(_5811_, _2879_, _2880_);
  xor g_6124_(_5811_, _2879_, _2881_);
  or g_6125_(_5734_, _5736_, _2882_);
  and g_6126_(G12[5], G11[12], _2883_);
  and g_6127_(G12[2], G11[15], _2884_);
  and g_6128_(G12[4], G11[15], _2885_);
  and g_6129_(_5622_, _2884_, _2887_);
  xor g_6130_(_5622_, _2884_, _2888_);
  and g_6131_(_2883_, _2888_, _2889_);
  xor g_6132_(_2883_, _2888_, _2890_);
  or g_6133_(_5730_, _5732_, _2891_);
  and g_6134_(G12[1], G11[16], _2892_);
  and g_6135_(G12[0], G11[17], _2893_);
  and g_6136_(G12[3], G11[17], _2894_);
  and g_6137_(_5539_, _2893_, _2895_);
  xor g_6138_(_5539_, _2893_, _2896_);
  and g_6139_(_2892_, _2896_, _2898_);
  xor g_6140_(_2892_, _2896_, _2899_);
  and g_6141_(_2891_, _2899_, _2900_);
  xor g_6142_(_2891_, _2899_, _2901_);
  and g_6143_(_2890_, _2901_, _2902_);
  xor g_6144_(_2890_, _2901_, _2903_);
  and g_6145_(_2882_, _2903_, _2904_);
  xor g_6146_(_2882_, _2903_, _2905_);
  and g_6147_(_2881_, _2905_, _2906_);
  xor g_6148_(_2881_, _2905_, _2907_);
  and g_6149_(_5810_, _2907_, _2908_);
  xor g_6150_(_5810_, _2907_, _2909_);
  and g_6151_(_5809_, _2909_, _2910_);
  xor g_6152_(_5809_, _2909_, _2911_);
  and g_6153_(_5782_, _2911_, _2912_);
  xor g_6154_(_5782_, _2911_, _2913_);
  and g_6155_(_5781_, _2913_, _2914_);
  xor g_6156_(_5781_, _2913_, _2915_);
  and g_6157_(_5763_, _2915_, _2916_);
  xor g_6158_(_5763_, _2915_, _2917_);
  and g_6159_(_5676_, _2917_, _2919_);
  xor g_6160_(_5676_, _2917_, _2920_);
  and g_6161_(_5762_, _2920_, _2921_);
  xor g_6162_(_5762_, _2920_, _2922_);
  and g_6163_(_5754_, _2922_, _2923_);
  xor g_6164_(_5754_, _2922_, _2924_);
  and g_6165_(_5756_, _2924_, _2925_);
  or g_6166_(_5756_, _2924_, _2926_);
  xor g_6167_(_5756_, _2924_, _2927_);
  xor g_6168_(_5761_, _2927_, G14[17]);
  and g_6169_(_5760_, _2927_, _2929_);
  and g_6170_(_5758_, _2926_, _2930_);
  or g_6171_(_2925_, _2930_, _2931_);
  or g_6172_(_2929_, _2931_, _2932_);
  or g_6173_(_2916_, _2919_, _2933_);
  or g_6174_(_5778_, _5780_, _2934_);
  or g_6175_(_2912_, _2914_, _2935_);
  and g_6176_(_5671_, _5775_, _2936_);
  and g_6177_(G11[0], G12[18], _2937_);
  or g_6178_(_5768_, _5770_, _2938_);
  and g_6179_(G11[1], G12[17], _2939_);
  and g_6180_(G11[3], G12[15], _2940_);
  and g_6181_(G11[3], G12[16], _2941_);
  and g_6182_(_5767_, _2940_, _2942_);
  xor g_6183_(_5767_, _2940_, _2943_);
  and g_6184_(_2939_, _2943_, _2944_);
  xor g_6185_(_2939_, _2943_, _2945_);
  or g_6186_(_5787_, _5789_, _2946_);
  and g_6187_(_2945_, _2946_, _2947_);
  xor g_6188_(_2945_, _2946_, _2948_);
  and g_6189_(_2938_, _2948_, _2950_);
  xor g_6190_(_2938_, _2948_, _2951_);
  or g_6191_(_5668_, _5773_, _2952_);
  and g_6192_(_5774_, _2952_, _2953_);
  and g_6193_(_2951_, _2953_, _2954_);
  xor g_6194_(_2951_, _2953_, _2955_);
  and g_6195_(_2937_, _2955_, _2956_);
  xor g_6196_(_2937_, _2955_, _2957_);
  or g_6197_(_5805_, _5808_, _2958_);
  and g_6198_(_2957_, _2958_, _2959_);
  xor g_6199_(_2957_, _2958_, _2961_);
  and g_6200_(_2936_, _2961_, _2962_);
  xor g_6201_(_2936_, _2961_, _2963_);
  or g_6202_(_2908_, _2910_, _2964_);
  or g_6203_(_5800_, _5802_, _2965_);
  and g_6204_(G11[4], G12[14], _2966_);
  and g_6205_(G11[6], G12[12], _2967_);
  and g_6206_(G11[6], G12[13], _2968_);
  and g_6207_(_5786_, _2967_, _2969_);
  xor g_6208_(_5786_, _2967_, _2970_);
  and g_6209_(_2966_, _2970_, _2972_);
  xor g_6210_(_2966_, _2970_, _2973_);
  or g_6211_(_5795_, _5798_, _2974_);
  and g_6212_(G11[7], G12[11], _2975_);
  and g_6213_(G11[9], G12[9], _2976_);
  and g_6214_(G11[9], G12[10], _2977_);
  and g_6215_(_5794_, _2976_, _2978_);
  xor g_6216_(_5794_, _2976_, _2979_);
  and g_6217_(_2975_, _2979_, _2980_);
  xor g_6218_(_2975_, _2979_, _2981_);
  and g_6219_(_2974_, _2981_, _2983_);
  xor g_6220_(_2974_, _2981_, _2984_);
  and g_6221_(_2973_, _2984_, _2985_);
  xor g_6222_(_2973_, _2984_, _2986_);
  or g_6223_(_2878_, _2880_, _2987_);
  and g_6224_(_2986_, _2987_, _2988_);
  xor g_6225_(_2986_, _2987_, _2989_);
  and g_6226_(_2965_, _2989_, _2990_);
  xor g_6227_(_2965_, _2989_, _2991_);
  or g_6228_(_2904_, _2906_, _2992_);
  or g_6229_(_5815_, _5817_, _2994_);
  and g_6230_(G12[8], G11[10], _2995_);
  and g_6231_(G12[6], G11[12], _2996_);
  and g_6232_(G12[7], G11[12], _2997_);
  and g_6233_(_5814_, _2996_, _2998_);
  xor g_6234_(_5814_, _2996_, _2999_);
  and g_6235_(_2995_, _2999_, _3000_);
  xor g_6236_(_2995_, _2999_, _3001_);
  or g_6237_(_2887_, _2889_, _3002_);
  and g_6238_(_3001_, _3002_, _3003_);
  xor g_6239_(_3001_, _3002_, _3005_);
  and g_6240_(_2994_, _3005_, _3006_);
  xor g_6241_(_2994_, _3005_, _3007_);
  or g_6242_(_2900_, _2902_, _3008_);
  and g_6243_(G12[5], G11[13], _3009_);
  and g_6244_(G12[2], G11[16], _3010_);
  and g_6245_(G12[4], G11[16], _3011_);
  and g_6246_(_5721_, _3010_, _3012_);
  xor g_6247_(_5721_, _3010_, _3013_);
  and g_6248_(_3009_, _3013_, _3014_);
  xor g_6249_(_3009_, _3013_, _3016_);
  or g_6250_(_2895_, _2898_, _3017_);
  and g_6251_(G12[1], G11[17], _3018_);
  and g_6252_(G12[0], G11[18], _3019_);
  and g_6253_(G12[3], G11[18], _3020_);
  and g_6254_(_5630_, _3019_, _3021_);
  xor g_6255_(_5630_, _3019_, _3022_);
  and g_6256_(_3018_, _3022_, _3023_);
  xor g_6257_(_3018_, _3022_, _3024_);
  and g_6258_(_3017_, _3024_, _3025_);
  xor g_6259_(_3017_, _3024_, _3027_);
  and g_6260_(_3016_, _3027_, _3028_);
  xor g_6261_(_3016_, _3027_, _3029_);
  and g_6262_(_3008_, _3029_, _3030_);
  xor g_6263_(_3008_, _3029_, _3031_);
  and g_6264_(_3007_, _3031_, _3032_);
  xor g_6265_(_3007_, _3031_, _3033_);
  and g_6266_(_2992_, _3033_, _3034_);
  xor g_6267_(_2992_, _3033_, _3035_);
  and g_6268_(_2991_, _3035_, _3036_);
  xor g_6269_(_2991_, _3035_, _3037_);
  and g_6270_(_2964_, _3037_, _3038_);
  xor g_6271_(_2964_, _3037_, _3039_);
  and g_6272_(_2963_, _3039_, _3040_);
  xor g_6273_(_2963_, _3039_, _3041_);
  and g_6274_(_2935_, _3041_, _3042_);
  xor g_6275_(_2935_, _3041_, _3043_);
  and g_6276_(_2934_, _3043_, _3044_);
  xor g_6277_(_2934_, _3043_, _3045_);
  and g_6278_(_2933_, _3045_, _3046_);
  xor g_6279_(_2933_, _3045_, _3048_);
  and g_6280_(_2921_, _3048_, _3049_);
  xor g_6281_(_2921_, _3048_, _3050_);
  and g_6282_(_2923_, _3050_, _3051_);
  xor g_6283_(_2923_, _3050_, _3052_);
  and g_6284_(_2932_, _3052_, _3053_);
  xor g_6285_(_2932_, _3052_, G14[18]);
  or g_6286_(_3051_, _3053_, _3054_);
  or g_6287_(_3042_, _3044_, _3055_);
  or g_6288_(_2959_, _2962_, _3056_);
  or g_6289_(_3038_, _3040_, _3058_);
  or g_6290_(_2954_, _2956_, _3059_);
  and g_6291_(G11[0], G12[19], _3060_);
  and g_6292_(G11[1], G12[18], _3061_);
  and g_6293_(G11[1], G12[19], _3062_);
  and g_6294_(_2937_, _3062_, _3063_);
  xor g_6295_(_3060_, _3061_, _3064_);
  or g_6296_(_2947_, _2950_, _3065_);
  or g_6297_(_2942_, _2944_, _3066_);
  and g_6298_(G11[2], G12[17], _3067_);
  and g_6299_(G11[4], G12[15], _3069_);
  and g_6300_(G11[4], G12[16], _3070_);
  and g_6301_(_2941_, _3069_, _3071_);
  xor g_6302_(_2941_, _3069_, _3072_);
  and g_6303_(_3067_, _3072_, _3073_);
  xor g_6304_(_3067_, _3072_, _3074_);
  or g_6305_(_2969_, _2972_, _3075_);
  and g_6306_(_3074_, _3075_, _3076_);
  xor g_6307_(_3074_, _3075_, _3077_);
  and g_6308_(_3066_, _3077_, _3078_);
  xor g_6309_(_3066_, _3077_, _3080_);
  and g_6310_(_3065_, _3080_, _3081_);
  xor g_6311_(_3065_, _3080_, _3082_);
  and g_6312_(_3064_, _3082_, _3083_);
  xor g_6313_(_3064_, _3082_, _3084_);
  or g_6314_(_2988_, _2990_, _3085_);
  and g_6315_(_3084_, _3085_, _3086_);
  xor g_6316_(_3084_, _3085_, _3087_);
  and g_6317_(_3059_, _3087_, _3088_);
  xor g_6318_(_3059_, _3087_, _3089_);
  or g_6319_(_3034_, _3036_, _3091_);
  or g_6320_(_2983_, _2985_, _3092_);
  and g_6321_(G11[5], G12[14], _3093_);
  and g_6322_(G11[7], G12[12], _3094_);
  and g_6323_(G11[7], G12[13], _3095_);
  and g_6324_(_2968_, _3094_, _3096_);
  xor g_6325_(_2968_, _3094_, _3097_);
  and g_6326_(_3093_, _3097_, _3098_);
  xor g_6327_(_3093_, _3097_, _3099_);
  or g_6328_(_2978_, _2980_, _3100_);
  and g_6329_(G11[8], G12[11], _3102_);
  and g_6330_(G11[10], G12[9], _3103_);
  and g_6331_(G11[10], G12[10], _3104_);
  and g_6332_(_2977_, _3103_, _3105_);
  xor g_6333_(_2977_, _3103_, _3106_);
  and g_6334_(_3102_, _3106_, _3107_);
  xor g_6335_(_3102_, _3106_, _3108_);
  and g_6336_(_3100_, _3108_, _3109_);
  xor g_6337_(_3100_, _3108_, _3110_);
  and g_6338_(_3099_, _3110_, _3111_);
  xor g_6339_(_3099_, _3110_, _3113_);
  or g_6340_(_3003_, _3006_, _3114_);
  and g_6341_(_3113_, _3114_, _3115_);
  xor g_6342_(_3113_, _3114_, _3116_);
  and g_6343_(_3092_, _3116_, _3117_);
  xor g_6344_(_3092_, _3116_, _3118_);
  or g_6345_(_3030_, _3032_, _3119_);
  or g_6346_(_2998_, _3000_, _3120_);
  and g_6347_(G12[8], G11[11], _3121_);
  and g_6348_(G12[6], G11[13], _3122_);
  and g_6349_(G12[7], G11[13], _3124_);
  and g_6350_(_2997_, _3122_, _3125_);
  xor g_6351_(_2997_, _3122_, _3126_);
  and g_6352_(_3121_, _3126_, _3127_);
  xor g_6353_(_3121_, _3126_, _3128_);
  or g_6354_(_3012_, _3014_, _3129_);
  and g_6355_(_3128_, _3129_, _3130_);
  xor g_6356_(_3128_, _3129_, _3131_);
  and g_6357_(_3120_, _3131_, _3132_);
  xor g_6358_(_3120_, _3131_, _3133_);
  or g_6359_(_3025_, _3028_, _3135_);
  and g_6360_(G12[5], G11[14], _3136_);
  and g_6361_(G12[2], G11[17], _3137_);
  and g_6362_(G12[4], G11[17], _3138_);
  and g_6363_(_2885_, _3137_, _3139_);
  xor g_6364_(_2885_, _3137_, _3140_);
  and g_6365_(_3136_, _3140_, _3141_);
  xor g_6366_(_3136_, _3140_, _3142_);
  or g_6367_(_3021_, _3023_, _3143_);
  and g_6368_(G12[1], G11[18], _3144_);
  and g_6369_(G12[0], G11[19], _3146_);
  and g_6370_(G12[3], G11[19], _3147_);
  and g_6371_(_5729_, _3146_, _3148_);
  xor g_6372_(_5729_, _3146_, _3149_);
  and g_6373_(_3144_, _3149_, _3150_);
  xor g_6374_(_3144_, _3149_, _3151_);
  and g_6375_(_3143_, _3151_, _3152_);
  xor g_6376_(_3143_, _3151_, _3153_);
  and g_6377_(_3142_, _3153_, _3154_);
  xor g_6378_(_3142_, _3153_, _3155_);
  and g_6379_(_3135_, _3155_, _3157_);
  xor g_6380_(_3135_, _3155_, _3158_);
  and g_6381_(_3133_, _3158_, _3159_);
  xor g_6382_(_3133_, _3158_, _3160_);
  and g_6383_(_3119_, _3160_, _3161_);
  xor g_6384_(_3119_, _3160_, _3162_);
  and g_6385_(_3118_, _3162_, _3163_);
  xor g_6386_(_3118_, _3162_, _3164_);
  and g_6387_(_3091_, _3164_, _3165_);
  xor g_6388_(_3091_, _3164_, _3166_);
  and g_6389_(_3089_, _3166_, _3168_);
  xor g_6390_(_3089_, _3166_, _3169_);
  and g_6391_(_3058_, _3169_, _3170_);
  xor g_6392_(_3058_, _3169_, _3171_);
  and g_6393_(_3056_, _3171_, _3172_);
  xor g_6394_(_3056_, _3171_, _3173_);
  and g_6395_(_3055_, _3173_, _3174_);
  xor g_6396_(_3055_, _3173_, _3175_);
  and g_6397_(_3046_, _3175_, _3176_);
  xor g_6398_(_3046_, _3175_, _3177_);
  and g_6399_(_3049_, _3177_, _3179_);
  xor g_6400_(_3049_, _3177_, _3180_);
  xor g_6401_(_3054_, _3180_, G14[19]);
  and g_6402_(_3053_, _3180_, _3181_);
  and g_6403_(_3051_, _3177_, _3182_);
  or g_6404_(_3179_, _3182_, _3183_);
  or g_6405_(_3181_, _3183_, _3184_);
  or g_6406_(_3170_, _3172_, _3185_);
  or g_6407_(_3086_, _3088_, _3186_);
  or g_6408_(_3165_, _3168_, _3187_);
  or g_6409_(_3081_, _3083_, _3189_);
  and g_6410_(G11[0], G12[20], _3190_);
  and g_6411_(G11[2], G12[18], _3191_);
  and g_6412_(G11[2], G12[19], _3192_);
  and g_6413_(_3062_, _3191_, _3193_);
  xor g_6414_(_3062_, _3191_, _3194_);
  and g_6415_(_3190_, _3194_, _3195_);
  xor g_6416_(_3190_, _3194_, _3196_);
  and g_6417_(_3063_, _3196_, _3197_);
  xor g_6418_(_3063_, _3196_, _3198_);
  or g_6419_(_3076_, _3078_, _3199_);
  or g_6420_(_3071_, _3073_, _3200_);
  and g_6421_(G11[3], G12[17], _3201_);
  and g_6422_(G11[5], G12[15], _3202_);
  and g_6423_(G11[5], G12[16], _3203_);
  and g_6424_(_3070_, _3202_, _3204_);
  xor g_6425_(_3070_, _3202_, _3205_);
  and g_6426_(_3201_, _3205_, _3206_);
  xor g_6427_(_3201_, _3205_, _3207_);
  or g_6428_(_3096_, _3098_, _3208_);
  and g_6429_(_3207_, _3208_, _3210_);
  xor g_6430_(_3207_, _3208_, _3211_);
  and g_6431_(_3200_, _3211_, _3212_);
  xor g_6432_(_3200_, _3211_, _3213_);
  and g_6433_(_3199_, _3213_, _3214_);
  xor g_6434_(_3199_, _3213_, _3215_);
  and g_6435_(_3198_, _3215_, _3216_);
  xor g_6436_(_3198_, _3215_, _3217_);
  or g_6437_(_3115_, _3117_, _3218_);
  and g_6438_(_3217_, _3218_, _3219_);
  xor g_6439_(_3217_, _3218_, _3221_);
  and g_6440_(_3189_, _3221_, _3222_);
  xor g_6441_(_3189_, _3221_, _3223_);
  or g_6442_(_3161_, _3163_, _3224_);
  or g_6443_(_3109_, _3111_, _3225_);
  and g_6444_(G11[6], G12[14], _3226_);
  and g_6445_(G11[8], G12[12], _3227_);
  and g_6446_(G11[8], G12[13], _3228_);
  and g_6447_(_3095_, _3227_, _3229_);
  xor g_6448_(_3095_, _3227_, _3230_);
  and g_6449_(_3226_, _3230_, _3232_);
  xor g_6450_(_3226_, _3230_, _3233_);
  or g_6451_(_3105_, _3107_, _3234_);
  and g_6452_(G11[9], G12[11], _3235_);
  and g_6453_(G12[9], G11[11], _3236_);
  and g_6454_(G12[10], G11[11], _3237_);
  and g_6455_(_3104_, _3236_, _3238_);
  xor g_6456_(_3104_, _3236_, _3239_);
  and g_6457_(_3235_, _3239_, _3240_);
  xor g_6458_(_3235_, _3239_, _3241_);
  and g_6459_(_3234_, _3241_, _3243_);
  xor g_6460_(_3234_, _3241_, _3244_);
  and g_6461_(_3233_, _3244_, _3245_);
  xor g_6462_(_3233_, _3244_, _3246_);
  or g_6463_(_3130_, _3132_, _3247_);
  and g_6464_(_3246_, _3247_, _3248_);
  xor g_6465_(_3246_, _3247_, _3249_);
  and g_6466_(_3225_, _3249_, _3250_);
  xor g_6467_(_3225_, _3249_, _3251_);
  or g_6468_(_3157_, _3159_, _3252_);
  or g_6469_(_3125_, _3127_, _3254_);
  and g_6470_(G12[8], G11[12], _3255_);
  and g_6471_(G12[6], G11[14], _3256_);
  and g_6472_(G12[7], G11[14], _3257_);
  and g_6473_(_3124_, _3256_, _3258_);
  xor g_6474_(_3124_, _3256_, _3259_);
  and g_6475_(_3255_, _3259_, _3260_);
  xor g_6476_(_3255_, _3259_, _3261_);
  or g_6477_(_3139_, _3141_, _3262_);
  and g_6478_(_3261_, _3262_, _3263_);
  xor g_6479_(_3261_, _3262_, _3265_);
  and g_6480_(_3254_, _3265_, _3266_);
  xor g_6481_(_3254_, _3265_, _3267_);
  or g_6482_(_3152_, _3154_, _3268_);
  and g_6483_(G12[5], G11[15], _3269_);
  and g_6484_(G12[2], G11[18], _3270_);
  and g_6485_(G12[4], G11[18], _3271_);
  and g_6486_(_3011_, _3270_, _3272_);
  xor g_6487_(_3011_, _3270_, _3273_);
  and g_6488_(_3269_, _3273_, _3274_);
  xor g_6489_(_3269_, _3273_, _3276_);
  or g_6490_(_3148_, _3150_, _3277_);
  and g_6491_(G12[1], G11[19], _3278_);
  and g_6492_(G12[0], G11[20], _3279_);
  and g_6493_(G12[3], G11[20], _3280_);
  and g_6494_(_2894_, _3279_, _3281_);
  xor g_6495_(_2894_, _3279_, _3282_);
  and g_6496_(_3278_, _3282_, _3283_);
  xor g_6497_(_3278_, _3282_, _3284_);
  and g_6498_(_3277_, _3284_, _3285_);
  xor g_6499_(_3277_, _3284_, _3287_);
  and g_6500_(_3276_, _3287_, _3288_);
  xor g_6501_(_3276_, _3287_, _3289_);
  and g_6502_(_3268_, _3289_, _3290_);
  xor g_6503_(_3268_, _3289_, _3291_);
  and g_6504_(_3267_, _3291_, _3292_);
  xor g_6505_(_3267_, _3291_, _3293_);
  and g_6506_(_3252_, _3293_, _3294_);
  xor g_6507_(_3252_, _3293_, _3295_);
  and g_6508_(_3251_, _3295_, _3296_);
  xor g_6509_(_3251_, _3295_, _3298_);
  and g_6510_(_3224_, _3298_, _3299_);
  xor g_6511_(_3224_, _3298_, _3300_);
  and g_6512_(_3223_, _3300_, _3301_);
  xor g_6513_(_3223_, _3300_, _3302_);
  and g_6514_(_3187_, _3302_, _3303_);
  xor g_6515_(_3187_, _3302_, _3304_);
  and g_6516_(_3186_, _3304_, _3305_);
  xor g_6517_(_3186_, _3304_, _3306_);
  and g_6518_(_3185_, _3306_, _3307_);
  xor g_6519_(_3185_, _3306_, _3309_);
  and g_6520_(_3174_, _3309_, _3310_);
  xor g_6521_(_3174_, _3309_, _3311_);
  and g_6522_(_3176_, _3311_, _3312_);
  xor g_6523_(_3176_, _3311_, _3313_);
  and g_6524_(_3184_, _3313_, _3314_);
  xor g_6525_(_3184_, _3313_, G14[20]);
  or g_6526_(_3312_, _3314_, _3315_);
  or g_6527_(_3303_, _3305_, _3316_);
  or g_6528_(_3219_, _3222_, _3317_);
  and g_6529_(_3197_, _3317_, _3319_);
  xor g_6530_(_3197_, _3317_, _3320_);
  or g_6531_(_3299_, _3301_, _3321_);
  or g_6532_(_3214_, _3216_, _3322_);
  and g_6533_(G11[0], G12[21], _3323_);
  or g_6534_(_3193_, _3195_, _3324_);
  and g_6535_(G11[1], G12[20], _3325_);
  and g_6536_(G11[3], G12[18], _3326_);
  and g_6537_(G11[3], G12[19], _3327_);
  and g_6538_(_3192_, _3326_, _3328_);
  xor g_6539_(_3192_, _3326_, _3330_);
  and g_6540_(_3325_, _3330_, _3331_);
  xor g_6541_(_3325_, _3330_, _3332_);
  and g_6542_(_3324_, _3332_, _3333_);
  xor g_6543_(_3324_, _3332_, _3334_);
  and g_6544_(_3323_, _3334_, _3335_);
  xor g_6545_(_3323_, _3334_, _3336_);
  or g_6546_(_3210_, _3212_, _3337_);
  or g_6547_(_3204_, _3206_, _3338_);
  and g_6548_(G11[4], G12[17], _3339_);
  and g_6549_(G11[6], G12[15], _3341_);
  and g_6550_(G11[6], G12[16], _3342_);
  and g_6551_(_3203_, _3341_, _3343_);
  xor g_6552_(_3203_, _3341_, _3344_);
  and g_6553_(_3339_, _3344_, _3345_);
  xor g_6554_(_3339_, _3344_, _3346_);
  or g_6555_(_3229_, _3232_, _3347_);
  and g_6556_(_3346_, _3347_, _3348_);
  xor g_6557_(_3346_, _3347_, _3349_);
  and g_6558_(_3338_, _3349_, _3350_);
  xor g_6559_(_3338_, _3349_, _3352_);
  and g_6560_(_3337_, _3352_, _3353_);
  xor g_6561_(_3337_, _3352_, _3354_);
  and g_6562_(_3336_, _3354_, _3355_);
  xor g_6563_(_3336_, _3354_, _3356_);
  or g_6564_(_3248_, _3250_, _3357_);
  and g_6565_(_3356_, _3357_, _3358_);
  xor g_6566_(_3356_, _3357_, _3359_);
  and g_6567_(_3322_, _3359_, _3360_);
  xor g_6568_(_3322_, _3359_, _3361_);
  or g_6569_(_3294_, _3296_, _3363_);
  or g_6570_(_3243_, _3245_, _3364_);
  and g_6571_(G11[7], G12[14], _3365_);
  and g_6572_(G11[9], G12[12], _3366_);
  and g_6573_(G11[9], G12[13], _3367_);
  and g_6574_(_3228_, _3366_, _3368_);
  xor g_6575_(_3228_, _3366_, _3369_);
  and g_6576_(_3365_, _3369_, _3370_);
  xor g_6577_(_3365_, _3369_, _3371_);
  or g_6578_(_3238_, _3240_, _3372_);
  and g_6579_(G11[10], G12[11], _3374_);
  and g_6580_(G12[9], G11[12], _3375_);
  and g_6581_(G12[10], G11[12], _3376_);
  and g_6582_(_3237_, _3375_, _3377_);
  xor g_6583_(_3237_, _3375_, _3378_);
  and g_6584_(_3374_, _3378_, _3379_);
  xor g_6585_(_3374_, _3378_, _3380_);
  and g_6586_(_3372_, _3380_, _3381_);
  xor g_6587_(_3372_, _3380_, _3382_);
  and g_6588_(_3371_, _3382_, _3383_);
  xor g_6589_(_3371_, _3382_, _3385_);
  or g_6590_(_3263_, _3266_, _3386_);
  and g_6591_(_3385_, _3386_, _3387_);
  xor g_6592_(_3385_, _3386_, _3388_);
  and g_6593_(_3364_, _3388_, _3389_);
  xor g_6594_(_3364_, _3388_, _3390_);
  or g_6595_(_3290_, _3292_, _3391_);
  or g_6596_(_3258_, _3260_, _3392_);
  and g_6597_(G12[8], G11[13], _3393_);
  and g_6598_(G12[6], G11[15], _3394_);
  and g_6599_(G12[7], G11[15], _3396_);
  and g_6600_(_3257_, _3394_, _3397_);
  xor g_6601_(_3257_, _3394_, _3398_);
  and g_6602_(_3393_, _3398_, _3399_);
  xor g_6603_(_3393_, _3398_, _3400_);
  or g_6604_(_3272_, _3274_, _3401_);
  and g_6605_(_3400_, _3401_, _3402_);
  xor g_6606_(_3400_, _3401_, _3403_);
  and g_6607_(_3392_, _3403_, _3404_);
  xor g_6608_(_3392_, _3403_, _3405_);
  or g_6609_(_3285_, _3288_, _3407_);
  and g_6610_(G12[5], G11[16], _3408_);
  and g_6611_(G12[2], G11[19], _3409_);
  and g_6612_(G12[4], G11[19], _3410_);
  and g_6613_(_3138_, _3409_, _3411_);
  xor g_6614_(_3138_, _3409_, _3412_);
  and g_6615_(_3408_, _3412_, _3413_);
  xor g_6616_(_3408_, _3412_, _3414_);
  or g_6617_(_3281_, _3283_, _3415_);
  and g_6618_(G12[1], G11[20], _3416_);
  and g_6619_(G12[0], G11[21], _3418_);
  and g_6620_(G12[3], G11[21], _3419_);
  and g_6621_(_3020_, _3418_, _3420_);
  xor g_6622_(_3020_, _3418_, _3421_);
  and g_6623_(_3416_, _3421_, _3422_);
  xor g_6624_(_3416_, _3421_, _3423_);
  and g_6625_(_3415_, _3423_, _3424_);
  xor g_6626_(_3415_, _3423_, _3425_);
  and g_6627_(_3414_, _3425_, _3426_);
  xor g_6628_(_3414_, _3425_, _3427_);
  and g_6629_(_3407_, _3427_, _3429_);
  xor g_6630_(_3407_, _3427_, _3430_);
  and g_6631_(_3405_, _3430_, _3431_);
  xor g_6632_(_3405_, _3430_, _3432_);
  and g_6633_(_3391_, _3432_, _3433_);
  xor g_6634_(_3391_, _3432_, _3434_);
  and g_6635_(_3390_, _3434_, _3435_);
  xor g_6636_(_3390_, _3434_, _3436_);
  and g_6637_(_3363_, _3436_, _3437_);
  xor g_6638_(_3363_, _3436_, _3438_);
  and g_6639_(_3361_, _3438_, _3440_);
  xor g_6640_(_3361_, _3438_, _3441_);
  and g_6641_(_3321_, _3441_, _3442_);
  xor g_6642_(_3321_, _3441_, _3443_);
  and g_6643_(_3320_, _3443_, _3444_);
  xor g_6644_(_3320_, _3443_, _3445_);
  and g_6645_(_3316_, _3445_, _3446_);
  xor g_6646_(_3316_, _3445_, _3447_);
  and g_6647_(_3307_, _3447_, _3448_);
  xor g_6648_(_3307_, _3447_, _3449_);
  and g_6649_(_3310_, _3449_, _3451_);
  xor g_6650_(_3310_, _3449_, _3452_);
  xor g_6651_(_3315_, _3452_, G14[21]);
  and g_6652_(_3314_, _3452_, _3453_);
  and g_6653_(_3312_, _3449_, _3454_);
  or g_6654_(_3451_, _3454_, _3455_);
  or g_6655_(_3453_, _3455_, _3456_);
  or g_6656_(_3442_, _3444_, _3457_);
  or g_6657_(_3333_, _3335_, _3458_);
  or g_6658_(_3358_, _3360_, _3459_);
  and g_6659_(_3458_, _3459_, _3461_);
  xor g_6660_(_3458_, _3459_, _3462_);
  or g_6661_(_3437_, _3440_, _3463_);
  or g_6662_(_3353_, _3355_, _3464_);
  and g_6663_(G11[0], G12[22], _3465_);
  and g_6664_(G11[1], G12[21], _3466_);
  and g_6665_(G11[1], G12[22], _3467_);
  and g_6666_(_3323_, _3467_, _3468_);
  xor g_6667_(_3465_, _3466_, _3469_);
  or g_6668_(_3328_, _3331_, _3470_);
  and g_6669_(G11[2], G12[20], _3471_);
  and g_6670_(G11[4], G12[18], _3472_);
  and g_6671_(G11[4], G12[19], _3473_);
  and g_6672_(_3327_, _3472_, _3474_);
  xor g_6673_(_3327_, _3472_, _3475_);
  and g_6674_(_3471_, _3475_, _3476_);
  xor g_6675_(_3471_, _3475_, _3477_);
  and g_6676_(_3470_, _3477_, _3478_);
  xor g_6677_(_3470_, _3477_, _3479_);
  and g_6678_(_3469_, _3479_, _3480_);
  xor g_6679_(_3469_, _3479_, _3482_);
  or g_6680_(_3348_, _3350_, _3483_);
  or g_6681_(_3343_, _3345_, _3484_);
  and g_6682_(G11[5], G12[17], _3485_);
  and g_6683_(G11[7], G12[15], _3486_);
  and g_6684_(G11[7], G12[16], _3487_);
  and g_6685_(_3342_, _3486_, _3488_);
  xor g_6686_(_3342_, _3486_, _3489_);
  and g_6687_(_3485_, _3489_, _3490_);
  xor g_6688_(_3485_, _3489_, _3491_);
  or g_6689_(_3368_, _3370_, _3493_);
  and g_6690_(_3491_, _3493_, _3494_);
  xor g_6691_(_3491_, _3493_, _3495_);
  and g_6692_(_3484_, _3495_, _3496_);
  xor g_6693_(_3484_, _3495_, _3497_);
  and g_6694_(_3483_, _3497_, _3498_);
  xor g_6695_(_3483_, _3497_, _3499_);
  and g_6696_(_3482_, _3499_, _3500_);
  xor g_6697_(_3482_, _3499_, _3501_);
  or g_6698_(_3387_, _3389_, _3502_);
  and g_6699_(_3501_, _3502_, _3504_);
  xor g_6700_(_3501_, _3502_, _3505_);
  and g_6701_(_3464_, _3505_, _3506_);
  xor g_6702_(_3464_, _3505_, _3507_);
  or g_6703_(_3433_, _3435_, _3508_);
  or g_6704_(_3381_, _3383_, _3509_);
  and g_6705_(G11[8], G12[14], _3510_);
  and g_6706_(G11[10], G12[12], _3511_);
  and g_6707_(G11[10], G12[13], _3512_);
  and g_6708_(_3367_, _3511_, _3513_);
  xor g_6709_(_3367_, _3511_, _3515_);
  and g_6710_(_3510_, _3515_, _3516_);
  xor g_6711_(_3510_, _3515_, _3517_);
  or g_6712_(_3377_, _3379_, _3518_);
  and g_6713_(G11[11], G12[11], _3519_);
  and g_6714_(G12[9], G11[13], _3520_);
  and g_6715_(G12[10], G11[13], _3521_);
  and g_6716_(_3376_, _3520_, _3522_);
  xor g_6717_(_3376_, _3520_, _3523_);
  and g_6718_(_3519_, _3523_, _3524_);
  xor g_6719_(_3519_, _3523_, _3526_);
  and g_6720_(_3518_, _3526_, _3527_);
  xor g_6721_(_3518_, _3526_, _3528_);
  and g_6722_(_3517_, _3528_, _3529_);
  xor g_6723_(_3517_, _3528_, _3530_);
  or g_6724_(_3402_, _3404_, _3531_);
  and g_6725_(_3530_, _3531_, _3532_);
  xor g_6726_(_3530_, _3531_, _3533_);
  and g_6727_(_3509_, _3533_, _3534_);
  xor g_6728_(_3509_, _3533_, _3535_);
  or g_6729_(_3429_, _3431_, _3537_);
  or g_6730_(_3397_, _3399_, _3538_);
  and g_6731_(G12[8], G11[14], _3539_);
  and g_6732_(G12[6], G11[16], _3540_);
  and g_6733_(G12[7], G11[16], _3541_);
  and g_6734_(_3396_, _3540_, _3542_);
  xor g_6735_(_3396_, _3540_, _3543_);
  and g_6736_(_3539_, _3543_, _3544_);
  xor g_6737_(_3539_, _3543_, _3545_);
  or g_6738_(_3411_, _3413_, _3546_);
  and g_6739_(_3545_, _3546_, _3548_);
  xor g_6740_(_3545_, _3546_, _3549_);
  and g_6741_(_3538_, _3549_, _3550_);
  xor g_6742_(_3538_, _3549_, _3551_);
  or g_6743_(_3424_, _3426_, _3552_);
  and g_6744_(G12[5], G11[17], _3553_);
  and g_6745_(G12[2], G11[20], _3554_);
  and g_6746_(G12[4], G11[20], _3555_);
  and g_6747_(_3271_, _3554_, _3556_);
  xor g_6748_(_3271_, _3554_, _3557_);
  and g_6749_(_3553_, _3557_, _3559_);
  xor g_6750_(_3553_, _3557_, _3560_);
  or g_6751_(_3420_, _3422_, _3561_);
  and g_6752_(G12[1], G11[21], _3562_);
  and g_6753_(G12[0], G11[22], _3563_);
  and g_6754_(G12[3], G11[22], _3564_);
  and g_6755_(_3147_, _3563_, _3565_);
  xor g_6756_(_3147_, _3563_, _3566_);
  and g_6757_(_3562_, _3566_, _3567_);
  xor g_6758_(_3562_, _3566_, _3568_);
  and g_6759_(_3561_, _3568_, _3570_);
  xor g_6760_(_3561_, _3568_, _3571_);
  and g_6761_(_3560_, _3571_, _3572_);
  xor g_6762_(_3560_, _3571_, _3573_);
  and g_6763_(_3552_, _3573_, _3574_);
  xor g_6764_(_3552_, _3573_, _3575_);
  and g_6765_(_3551_, _3575_, _3576_);
  xor g_6766_(_3551_, _3575_, _3577_);
  and g_6767_(_3537_, _3577_, _3578_);
  xor g_6768_(_3537_, _3577_, _3579_);
  and g_6769_(_3535_, _3579_, _3581_);
  xor g_6770_(_3535_, _3579_, _3582_);
  and g_6771_(_3508_, _3582_, _3583_);
  xor g_6772_(_3508_, _3582_, _3584_);
  and g_6773_(_3507_, _3584_, _3585_);
  xor g_6774_(_3507_, _3584_, _3586_);
  and g_6775_(_3463_, _3586_, _3587_);
  xor g_6776_(_3463_, _3586_, _3588_);
  and g_6777_(_3462_, _3588_, _3589_);
  xor g_6778_(_3462_, _3588_, _3590_);
  and g_6779_(_3457_, _3590_, _3592_);
  xor g_6780_(_3457_, _3590_, _3593_);
  and g_6781_(_3319_, _3593_, _3594_);
  xor g_6782_(_3319_, _3593_, _3595_);
  and g_6783_(_3446_, _3595_, _3596_);
  xor g_6784_(_3446_, _3595_, _3597_);
  and g_6785_(_3448_, _3597_, _3598_);
  xor g_6786_(_3448_, _3597_, _3599_);
  and g_6787_(_3456_, _3599_, _3600_);
  xor g_6788_(_3456_, _3599_, G14[22]);
  or g_6789_(_3598_, _3600_, _3602_);
  or g_6790_(_3592_, _3594_, _3603_);
  or g_6791_(_3587_, _3589_, _3604_);
  or g_6792_(_3504_, _3506_, _3605_);
  and g_6793_(_3468_, _3478_, _3606_);
  xor g_6794_(_3468_, _3478_, _3607_);
  or g_6795_(_3480_, _3607_, _3608_);
  and g_6796_(_3605_, _3608_, _3609_);
  xor g_6797_(_3605_, _3608_, _3610_);
  or g_6798_(_3583_, _3585_, _3611_);
  or g_6799_(_3498_, _3500_, _3613_);
  and g_6800_(G11[0], G12[23], _3614_);
  and g_6801_(G11[2], G12[21], _3615_);
  and g_6802_(G11[2], G12[22], _3616_);
  and g_6803_(_3467_, _3615_, _3617_);
  xor g_6804_(_3467_, _3615_, _3618_);
  and g_6805_(_3614_, _3618_, _3619_);
  xor g_6806_(_3614_, _3618_, _3620_);
  or g_6807_(_3474_, _3476_, _3621_);
  and g_6808_(G11[3], G12[20], _3622_);
  and g_6809_(G11[5], G12[18], _3624_);
  and g_6810_(G11[5], G12[19], _3625_);
  and g_6811_(_3473_, _3624_, _3626_);
  xor g_6812_(_3473_, _3624_, _3627_);
  and g_6813_(_3622_, _3627_, _3628_);
  xor g_6814_(_3622_, _3627_, _3629_);
  and g_6815_(_3621_, _3629_, _3630_);
  xor g_6816_(_3621_, _3629_, _3631_);
  and g_6817_(_3620_, _3631_, _3632_);
  xor g_6818_(_3620_, _3631_, _3633_);
  or g_6819_(_3494_, _3496_, _3635_);
  or g_6820_(_3488_, _3490_, _3636_);
  and g_6821_(G11[6], G12[17], _3637_);
  and g_6822_(G11[8], G12[15], _3638_);
  and g_6823_(G11[8], G12[16], _3639_);
  and g_6824_(_3487_, _3638_, _3640_);
  xor g_6825_(_3487_, _3638_, _3641_);
  and g_6826_(_3637_, _3641_, _3642_);
  xor g_6827_(_3637_, _3641_, _3643_);
  or g_6828_(_3513_, _3516_, _3644_);
  and g_6829_(_3643_, _3644_, _3646_);
  xor g_6830_(_3643_, _3644_, _3647_);
  and g_6831_(_3636_, _3647_, _3648_);
  xor g_6832_(_3636_, _3647_, _3649_);
  and g_6833_(_3635_, _3649_, _3650_);
  xor g_6834_(_3635_, _3649_, _3651_);
  and g_6835_(_3633_, _3651_, _3652_);
  xor g_6836_(_3633_, _3651_, _3653_);
  or g_6837_(_3532_, _3534_, _3654_);
  and g_6838_(_3653_, _3654_, _3655_);
  xor g_6839_(_3653_, _3654_, _3657_);
  and g_6840_(_3613_, _3657_, _3658_);
  xor g_6841_(_3613_, _3657_, _3659_);
  or g_6842_(_3578_, _3581_, _3660_);
  or g_6843_(_3527_, _3529_, _3661_);
  and g_6844_(G11[9], G12[14], _3662_);
  and g_6845_(G11[11], G12[12], _3663_);
  and g_6846_(G11[11], G12[13], _3664_);
  and g_6847_(_3512_, _3663_, _3665_);
  xor g_6848_(_3512_, _3663_, _3666_);
  and g_6849_(_3662_, _3666_, _3668_);
  xor g_6850_(_3662_, _3666_, _3669_);
  or g_6851_(_3522_, _3524_, _3670_);
  and g_6852_(G12[11], G11[12], _3671_);
  and g_6853_(G12[9], G11[14], _3672_);
  and g_6854_(G12[10], G11[14], _3673_);
  and g_6855_(_3521_, _3672_, _3674_);
  xor g_6856_(_3521_, _3672_, _3675_);
  and g_6857_(_3671_, _3675_, _3676_);
  xor g_6858_(_3671_, _3675_, _3677_);
  and g_6859_(_3670_, _3677_, _3679_);
  xor g_6860_(_3670_, _3677_, _3680_);
  and g_6861_(_3669_, _3680_, _3681_);
  xor g_6862_(_3669_, _3680_, _3682_);
  or g_6863_(_3548_, _3550_, _3683_);
  and g_6864_(_3682_, _3683_, _3684_);
  xor g_6865_(_3682_, _3683_, _3685_);
  and g_6866_(_3661_, _3685_, _3686_);
  xor g_6867_(_3661_, _3685_, _3687_);
  or g_6868_(_3574_, _3576_, _3688_);
  or g_6869_(_3542_, _3544_, _3690_);
  and g_6870_(G12[8], G11[15], _3691_);
  and g_6871_(G12[6], G11[17], _3692_);
  and g_6872_(G12[7], G11[17], _3693_);
  and g_6873_(_3541_, _3692_, _3694_);
  xor g_6874_(_3541_, _3692_, _3695_);
  and g_6875_(_3691_, _3695_, _3696_);
  xor g_6876_(_3691_, _3695_, _3697_);
  or g_6877_(_3556_, _3559_, _3698_);
  and g_6878_(_3697_, _3698_, _3699_);
  xor g_6879_(_3697_, _3698_, _3701_);
  and g_6880_(_3690_, _3701_, _3702_);
  xor g_6881_(_3690_, _3701_, _3703_);
  or g_6882_(_3570_, _3572_, _3704_);
  and g_6883_(G12[5], G11[18], _3705_);
  and g_6884_(G12[2], G11[21], _3706_);
  and g_6885_(G12[4], G11[21], _3707_);
  and g_6886_(_3410_, _3706_, _3708_);
  xor g_6887_(_3410_, _3706_, _3709_);
  and g_6888_(_3705_, _3709_, _3710_);
  xor g_6889_(_3705_, _3709_, _3712_);
  or g_6890_(_3565_, _3567_, _3713_);
  and g_6891_(G12[1], G11[22], _3714_);
  and g_6892_(G12[0], G11[23], _3715_);
  and g_6893_(G12[3], G11[23], _3716_);
  and g_6894_(_3280_, _3715_, _3717_);
  xor g_6895_(_3280_, _3715_, _3718_);
  and g_6896_(_3714_, _3718_, _3719_);
  xor g_6897_(_3714_, _3718_, _3720_);
  and g_6898_(_3713_, _3720_, _3721_);
  xor g_6899_(_3713_, _3720_, _3723_);
  and g_6900_(_3712_, _3723_, _3724_);
  xor g_6901_(_3712_, _3723_, _3725_);
  and g_6902_(_3704_, _3725_, _3726_);
  xor g_6903_(_3704_, _3725_, _3727_);
  and g_6904_(_3703_, _3727_, _3728_);
  xor g_6905_(_3703_, _3727_, _3729_);
  and g_6906_(_3688_, _3729_, _3730_);
  xor g_6907_(_3688_, _3729_, _3731_);
  and g_6908_(_3687_, _3731_, _3732_);
  xor g_6909_(_3687_, _3731_, _3734_);
  and g_6910_(_3660_, _3734_, _3735_);
  xor g_6911_(_3660_, _3734_, _3736_);
  and g_6912_(_3659_, _3736_, _3737_);
  xor g_6913_(_3659_, _3736_, _3738_);
  and g_6914_(_3611_, _3738_, _3739_);
  xor g_6915_(_3611_, _3738_, _3740_);
  and g_6916_(_3610_, _3740_, _3741_);
  xor g_6917_(_3610_, _3740_, _3742_);
  and g_6918_(_3604_, _3742_, _3743_);
  xor g_6919_(_3604_, _3742_, _3745_);
  and g_6920_(_3461_, _3745_, _3746_);
  xor g_6921_(_3461_, _3745_, _3747_);
  and g_6922_(_3603_, _3747_, _3748_);
  xor g_6923_(_3603_, _3747_, _3749_);
  and g_6924_(_3596_, _3749_, _3750_);
  xor g_6925_(_3596_, _3749_, _3751_);
  and g_6926_(_3602_, _3751_, _3752_);
  xor g_6927_(_3602_, _3751_, G14[23]);
  or g_6928_(_3743_, _3746_, _3753_);
  or g_6929_(_3739_, _3741_, _3755_);
  and g_6930_(G11[0], G12[24], _3756_);
  or g_6931_(_3617_, _3619_, _3757_);
  and g_6932_(_3756_, _3757_, _3758_);
  xor g_6933_(_3756_, _3757_, _3759_);
  or g_6934_(_3630_, _3632_, _3760_);
  and g_6935_(_3759_, _3760_, _3761_);
  xor g_6936_(_3759_, _3760_, _3762_);
  and g_6937_(_3606_, _3762_, _3763_);
  xor g_6938_(_3606_, _3762_, _3764_);
  or g_6939_(_3655_, _3658_, _3766_);
  and g_6940_(_3764_, _3766_, _3767_);
  xor g_6941_(_3764_, _3766_, _3768_);
  or g_6942_(_3735_, _3737_, _3769_);
  or g_6943_(_3650_, _3652_, _3770_);
  and g_6944_(G11[1], G12[23], _3771_);
  and g_6945_(G11[3], G12[21], _3772_);
  and g_6946_(G11[3], G12[22], _3773_);
  and g_6947_(_3616_, _3772_, _3774_);
  xor g_6948_(_3616_, _3772_, _3775_);
  and g_6949_(_3771_, _3775_, _3776_);
  xor g_6950_(_3771_, _3775_, _3777_);
  or g_6951_(_3626_, _3628_, _3778_);
  and g_6952_(G11[4], G12[20], _3779_);
  and g_6953_(G11[6], G12[18], _3780_);
  and g_6954_(G11[6], G12[19], _3781_);
  and g_6955_(_3625_, _3780_, _3782_);
  xor g_6956_(_3625_, _3780_, _3783_);
  and g_6957_(_3779_, _3783_, _3784_);
  xor g_6958_(_3779_, _3783_, _3785_);
  and g_6959_(_3778_, _3785_, _3787_);
  xor g_6960_(_3778_, _3785_, _3788_);
  and g_6961_(_3777_, _3788_, _3789_);
  xor g_6962_(_3777_, _3788_, _3790_);
  or g_6963_(_3646_, _3648_, _3791_);
  or g_6964_(_3640_, _3642_, _3792_);
  and g_6965_(G11[7], G12[17], _3793_);
  and g_6966_(G11[9], G12[15], _3794_);
  and g_6967_(G11[9], G12[16], _3795_);
  and g_6968_(_3639_, _3794_, _3796_);
  xor g_6969_(_3639_, _3794_, _3798_);
  and g_6970_(_3793_, _3798_, _3799_);
  xor g_6971_(_3793_, _3798_, _3800_);
  or g_6972_(_3665_, _3668_, _3801_);
  and g_6973_(_3800_, _3801_, _3802_);
  xor g_6974_(_3800_, _3801_, _3803_);
  and g_6975_(_3792_, _3803_, _3804_);
  xor g_6976_(_3792_, _3803_, _3805_);
  and g_6977_(_3791_, _3805_, _3806_);
  xor g_6978_(_3791_, _3805_, _3807_);
  and g_6979_(_3790_, _3807_, _3809_);
  xor g_6980_(_3790_, _3807_, _3810_);
  or g_6981_(_3684_, _3686_, _3811_);
  and g_6982_(_3810_, _3811_, _3812_);
  xor g_6983_(_3810_, _3811_, _3813_);
  and g_6984_(_3770_, _3813_, _3814_);
  xor g_6985_(_3770_, _3813_, _3815_);
  or g_6986_(_3730_, _3732_, _3816_);
  or g_6987_(_3679_, _3681_, _3817_);
  and g_6988_(G11[10], G12[14], _3818_);
  and g_6989_(G11[12], G12[12], _3820_);
  and g_6990_(G11[12], G12[13], _3821_);
  and g_6991_(_3664_, _3820_, _3822_);
  xor g_6992_(_3664_, _3820_, _3823_);
  and g_6993_(_3818_, _3823_, _3824_);
  xor g_6994_(_3818_, _3823_, _3825_);
  or g_6995_(_3674_, _3676_, _3826_);
  and g_6996_(G12[11], G11[13], _3827_);
  and g_6997_(G12[9], G11[15], _3828_);
  and g_6998_(G12[10], G11[15], _3829_);
  and g_6999_(_3673_, _3828_, _3831_);
  xor g_7000_(_3673_, _3828_, _3832_);
  and g_7001_(_3827_, _3832_, _3833_);
  xor g_7002_(_3827_, _3832_, _3834_);
  and g_7003_(_3826_, _3834_, _3835_);
  xor g_7004_(_3826_, _3834_, _3836_);
  and g_7005_(_3825_, _3836_, _3837_);
  xor g_7006_(_3825_, _3836_, _3838_);
  or g_7007_(_3699_, _3702_, _3839_);
  and g_7008_(_3838_, _3839_, _3840_);
  xor g_7009_(_3838_, _3839_, _3842_);
  and g_7010_(_3817_, _3842_, _3843_);
  xor g_7011_(_3817_, _3842_, _3844_);
  or g_7012_(_3726_, _3728_, _3845_);
  or g_7013_(_3694_, _3696_, _3846_);
  and g_7014_(G12[8], G11[16], _3847_);
  and g_7015_(G12[6], G11[18], _3848_);
  and g_7016_(G12[7], G11[18], _3849_);
  and g_7017_(_3693_, _3848_, _3850_);
  xor g_7018_(_3693_, _3848_, _3851_);
  and g_7019_(_3847_, _3851_, _3853_);
  xor g_7020_(_3847_, _3851_, _3854_);
  or g_7021_(_3708_, _3710_, _3855_);
  and g_7022_(_3854_, _3855_, _3856_);
  xor g_7023_(_3854_, _3855_, _3857_);
  and g_7024_(_3846_, _3857_, _3858_);
  xor g_7025_(_3846_, _3857_, _3859_);
  or g_7026_(_3721_, _3724_, _3860_);
  and g_7027_(G12[5], G11[19], _3861_);
  and g_7028_(G12[2], G11[22], _3862_);
  and g_7029_(G12[4], G11[22], _3864_);
  and g_7030_(_3555_, _3862_, _3865_);
  xor g_7031_(_3555_, _3862_, _3866_);
  and g_7032_(_3861_, _3866_, _3867_);
  xor g_7033_(_3861_, _3866_, _3868_);
  or g_7034_(_3717_, _3719_, _3869_);
  and g_7035_(G12[1], G11[23], _3870_);
  and g_7036_(G12[0], G11[24], _3871_);
  and g_7037_(G12[3], G11[24], _3872_);
  and g_7038_(_3419_, _3871_, _3873_);
  xor g_7039_(_3419_, _3871_, _3875_);
  and g_7040_(_3870_, _3875_, _3876_);
  xor g_7041_(_3870_, _3875_, _3877_);
  and g_7042_(_3869_, _3877_, _3878_);
  xor g_7043_(_3869_, _3877_, _3879_);
  and g_7044_(_3868_, _3879_, _3880_);
  xor g_7045_(_3868_, _3879_, _3881_);
  and g_7046_(_3860_, _3881_, _3882_);
  xor g_7047_(_3860_, _3881_, _3883_);
  and g_7048_(_3859_, _3883_, _3884_);
  xor g_7049_(_3859_, _3883_, _3886_);
  and g_7050_(_3845_, _3886_, _3887_);
  xor g_7051_(_3845_, _3886_, _3888_);
  and g_7052_(_3844_, _3888_, _3889_);
  xor g_7053_(_3844_, _3888_, _3890_);
  and g_7054_(_3816_, _3890_, _3891_);
  xor g_7055_(_3816_, _3890_, _3892_);
  and g_7056_(_3815_, _3892_, _3893_);
  xor g_7057_(_3815_, _3892_, _3894_);
  and g_7058_(_3769_, _3894_, _3895_);
  xor g_7059_(_3769_, _3894_, _3897_);
  and g_7060_(_3768_, _3897_, _3898_);
  xor g_7061_(_3768_, _3897_, _3899_);
  and g_7062_(_3755_, _3899_, _3900_);
  xor g_7063_(_3755_, _3899_, _3901_);
  and g_7064_(_3609_, _3901_, _3902_);
  xor g_7065_(_3609_, _3901_, _3903_);
  and g_7066_(_3753_, _3903_, _3904_);
  xor g_7067_(_3753_, _3903_, _3905_);
  and g_7068_(_3748_, _3905_, _3906_);
  xor g_7069_(_3748_, _3905_, _3908_);
  or g_7070_(_3750_, _3752_, _3909_);
  and g_7071_(_3908_, _3909_, _3910_);
  xor g_7072_(_3908_, _3909_, G14[24]);
  or g_7073_(_3906_, _3910_, _3911_);
  or g_7074_(_3900_, _3902_, _3912_);
  or g_7075_(_3895_, _3898_, _3913_);
  or g_7076_(_3812_, _3814_, _3914_);
  and g_7077_(G11[0], G12[25], _3915_);
  and g_7078_(G11[1], G12[24], _3916_);
  and g_7079_(G11[1], G12[25], _3918_);
  and g_7080_(_3756_, _3918_, _3919_);
  xor g_7081_(_3915_, _3916_, _3920_);
  or g_7082_(_3774_, _3776_, _3921_);
  and g_7083_(_3920_, _3921_, _3922_);
  xor g_7084_(_3920_, _3921_, _3923_);
  or g_7085_(_3787_, _3789_, _3924_);
  and g_7086_(_3923_, _3924_, _3925_);
  or g_7087_(_3923_, _3924_, _3926_);
  xor g_7088_(_3923_, _3924_, _3927_);
  or g_7089_(_3758_, _3761_, _3929_);
  xor g_7090_(_3927_, _3929_, _3930_);
  and g_7091_(_3914_, _3930_, _3931_);
  xor g_7092_(_3914_, _3930_, _3932_);
  and g_7093_(_3763_, _3932_, _3933_);
  xor g_7094_(_3763_, _3932_, _3934_);
  or g_7095_(_3891_, _3893_, _3935_);
  or g_7096_(_3806_, _3809_, _3936_);
  and g_7097_(G11[2], G12[23], _3937_);
  and g_7098_(G11[4], G12[21], _3938_);
  and g_7099_(G11[4], G12[22], _3940_);
  and g_7100_(_3773_, _3938_, _3941_);
  xor g_7101_(_3773_, _3938_, _3942_);
  and g_7102_(_3937_, _3942_, _3943_);
  xor g_7103_(_3937_, _3942_, _3944_);
  or g_7104_(_3782_, _3784_, _3945_);
  and g_7105_(G11[5], G12[20], _3946_);
  and g_7106_(G11[7], G12[18], _3947_);
  and g_7107_(G11[7], G12[19], _3948_);
  and g_7108_(_3781_, _3947_, _3949_);
  xor g_7109_(_3781_, _3947_, _3951_);
  and g_7110_(_3946_, _3951_, _3952_);
  xor g_7111_(_3946_, _3951_, _3953_);
  and g_7112_(_3945_, _3953_, _3954_);
  xor g_7113_(_3945_, _3953_, _3955_);
  and g_7114_(_3944_, _3955_, _3956_);
  xor g_7115_(_3944_, _3955_, _3957_);
  or g_7116_(_3802_, _3804_, _3958_);
  or g_7117_(_3796_, _3799_, _3959_);
  and g_7118_(G11[8], G12[17], _3960_);
  and g_7119_(G11[10], G12[15], _3962_);
  and g_7120_(G11[10], G12[16], _3963_);
  and g_7121_(_3795_, _3962_, _3964_);
  xor g_7122_(_3795_, _3962_, _3965_);
  and g_7123_(_3960_, _3965_, _3966_);
  xor g_7124_(_3960_, _3965_, _3967_);
  or g_7125_(_3822_, _3824_, _3968_);
  and g_7126_(_3967_, _3968_, _3969_);
  xor g_7127_(_3967_, _3968_, _3970_);
  and g_7128_(_3959_, _3970_, _3971_);
  xor g_7129_(_3959_, _3970_, _3973_);
  and g_7130_(_3958_, _3973_, _3974_);
  xor g_7131_(_3958_, _3973_, _3975_);
  and g_7132_(_3957_, _3975_, _3976_);
  xor g_7133_(_3957_, _3975_, _3977_);
  or g_7134_(_3840_, _3843_, _3978_);
  and g_7135_(_3977_, _3978_, _3979_);
  xor g_7136_(_3977_, _3978_, _3980_);
  and g_7137_(_3936_, _3980_, _3981_);
  xor g_7138_(_3936_, _3980_, _3982_);
  or g_7139_(_3887_, _3889_, _3984_);
  or g_7140_(_3835_, _3837_, _3985_);
  and g_7141_(G11[11], G12[14], _3986_);
  and g_7142_(G12[12], G11[13], _3987_);
  and g_7143_(G11[13], G12[13], _3988_);
  and g_7144_(_3821_, _3987_, _3989_);
  xor g_7145_(_3821_, _3987_, _3990_);
  and g_7146_(_3986_, _3990_, _3991_);
  xor g_7147_(_3986_, _3990_, _3992_);
  or g_7148_(_3831_, _3833_, _3993_);
  and g_7149_(G12[11], G11[14], _3995_);
  and g_7150_(G12[9], G11[16], _3996_);
  and g_7151_(G12[10], G11[16], _3997_);
  and g_7152_(_3829_, _3996_, _3998_);
  xor g_7153_(_3829_, _3996_, _3999_);
  and g_7154_(_3995_, _3999_, _4000_);
  xor g_7155_(_3995_, _3999_, _4001_);
  and g_7156_(_3993_, _4001_, _4002_);
  xor g_7157_(_3993_, _4001_, _4003_);
  and g_7158_(_3992_, _4003_, _4004_);
  xor g_7159_(_3992_, _4003_, _4006_);
  or g_7160_(_3856_, _3858_, _4007_);
  and g_7161_(_4006_, _4007_, _4008_);
  xor g_7162_(_4006_, _4007_, _4009_);
  and g_7163_(_3985_, _4009_, _4010_);
  xor g_7164_(_3985_, _4009_, _4011_);
  or g_7165_(_3882_, _3884_, _4012_);
  or g_7166_(_3850_, _3853_, _4013_);
  and g_7167_(G12[8], G11[17], _4014_);
  and g_7168_(G12[6], G11[19], _4015_);
  and g_7169_(G12[7], G11[19], _4017_);
  and g_7170_(_3849_, _4015_, _4018_);
  xor g_7171_(_3849_, _4015_, _4019_);
  and g_7172_(_4014_, _4019_, _4020_);
  xor g_7173_(_4014_, _4019_, _4021_);
  or g_7174_(_3865_, _3867_, _4022_);
  and g_7175_(_4021_, _4022_, _4023_);
  xor g_7176_(_4021_, _4022_, _4024_);
  and g_7177_(_4013_, _4024_, _4025_);
  xor g_7178_(_4013_, _4024_, _4026_);
  or g_7179_(_3878_, _3880_, _4028_);
  and g_7180_(G12[5], G11[20], _4029_);
  and g_7181_(G12[2], G11[23], _4030_);
  and g_7182_(G12[4], G11[23], _4031_);
  and g_7183_(_3707_, _4030_, _4032_);
  xor g_7184_(_3707_, _4030_, _4033_);
  and g_7185_(_4029_, _4033_, _4034_);
  xor g_7186_(_4029_, _4033_, _4035_);
  or g_7187_(_3873_, _3876_, _4036_);
  and g_7188_(G12[1], G11[24], _4037_);
  and g_7189_(G12[0], G11[25], _4039_);
  and g_7190_(G12[3], G11[25], _4040_);
  and g_7191_(_3564_, _4039_, _4041_);
  xor g_7192_(_3564_, _4039_, _4042_);
  and g_7193_(_4037_, _4042_, _4043_);
  xor g_7194_(_4037_, _4042_, _4044_);
  and g_7195_(_4036_, _4044_, _4045_);
  xor g_7196_(_4036_, _4044_, _4046_);
  and g_7197_(_4035_, _4046_, _4047_);
  xor g_7198_(_4035_, _4046_, _4048_);
  and g_7199_(_4028_, _4048_, _4050_);
  xor g_7200_(_4028_, _4048_, _4051_);
  and g_7201_(_4026_, _4051_, _4052_);
  xor g_7202_(_4026_, _4051_, _4053_);
  and g_7203_(_4012_, _4053_, _4054_);
  xor g_7204_(_4012_, _4053_, _4055_);
  and g_7205_(_4011_, _4055_, _4056_);
  xor g_7206_(_4011_, _4055_, _4057_);
  and g_7207_(_3984_, _4057_, _4058_);
  xor g_7208_(_3984_, _4057_, _4059_);
  and g_7209_(_3982_, _4059_, _4061_);
  xor g_7210_(_3982_, _4059_, _4062_);
  and g_7211_(_3935_, _4062_, _4063_);
  xor g_7212_(_3935_, _4062_, _4064_);
  and g_7213_(_3934_, _4064_, _4065_);
  xor g_7214_(_3934_, _4064_, _4066_);
  and g_7215_(_3913_, _4066_, _4067_);
  xor g_7216_(_3913_, _4066_, _4068_);
  and g_7217_(_3767_, _4068_, _4069_);
  xor g_7218_(_3767_, _4068_, _4070_);
  and g_7219_(_3912_, _4070_, _4072_);
  xor g_7220_(_3912_, _4070_, _4073_);
  and g_7221_(_3904_, _4073_, _4074_);
  xor g_7222_(_3904_, _4073_, _4075_);
  and g_7223_(_3911_, _4075_, _4076_);
  xor g_7224_(_3911_, _4075_, G14[25]);
  or g_7225_(_4067_, _4069_, _4077_);
  or g_7226_(_3931_, _3933_, _4078_);
  or g_7227_(_4063_, _4065_, _4079_);
  and g_7228_(_3761_, _3927_, _4080_);
  and g_7229_(G11[0], G12[26], _4082_);
  and g_7230_(G11[2], G12[24], _4083_);
  and g_7231_(G11[2], G12[25], _4084_);
  and g_7232_(_3918_, _4083_, _4085_);
  xor g_7233_(_3918_, _4083_, _4086_);
  and g_7234_(_4082_, _4086_, _4087_);
  xor g_7235_(_4082_, _4086_, _4088_);
  or g_7236_(_3941_, _3943_, _4089_);
  and g_7237_(_4088_, _4089_, _4090_);
  xor g_7238_(_4088_, _4089_, _4091_);
  and g_7239_(_3919_, _4091_, _4093_);
  xor g_7240_(_3919_, _4091_, _4094_);
  or g_7241_(_3954_, _3956_, _4095_);
  and g_7242_(_4094_, _4095_, _4096_);
  xor g_7243_(_4094_, _4095_, _4097_);
  and g_7244_(_3922_, _4097_, _4098_);
  xor g_7245_(_3922_, _4097_, _4099_);
  not g_7246_(_4099_, _4100_);
  or g_7247_(_3758_, _3925_, _4101_);
  and g_7248_(_3926_, _4101_, _4102_);
  and g_7249_(_4099_, _4102_, _4104_);
  xor g_7250_(_4099_, _4102_, _4105_);
  xor g_7251_(_4100_, _4102_, _4106_);
  or g_7252_(_3979_, _3981_, _4107_);
  and g_7253_(_4105_, _4107_, _4108_);
  xor g_7254_(_4106_, _4107_, _4109_);
  not g_7255_(_4109_, _4110_);
  and g_7256_(_4080_, _4110_, _4111_);
  xor g_7257_(_4080_, _4110_, _4112_);
  or g_7258_(_4058_, _4061_, _4113_);
  or g_7259_(_3974_, _3976_, _4115_);
  and g_7260_(G11[3], G12[23], _4116_);
  and g_7261_(G11[5], G12[21], _4117_);
  and g_7262_(G11[5], G12[22], _4118_);
  and g_7263_(_3940_, _4117_, _4119_);
  xor g_7264_(_3940_, _4117_, _4120_);
  and g_7265_(_4116_, _4120_, _4121_);
  xor g_7266_(_4116_, _4120_, _4122_);
  or g_7267_(_3949_, _3952_, _4123_);
  and g_7268_(G11[6], G12[20], _4124_);
  and g_7269_(G11[8], G12[18], _4126_);
  and g_7270_(G11[8], G12[19], _4127_);
  and g_7271_(_3948_, _4126_, _4128_);
  xor g_7272_(_3948_, _4126_, _4129_);
  and g_7273_(_4124_, _4129_, _4130_);
  xor g_7274_(_4124_, _4129_, _4131_);
  and g_7275_(_4123_, _4131_, _4132_);
  xor g_7276_(_4123_, _4131_, _4133_);
  and g_7277_(_4122_, _4133_, _4134_);
  xor g_7278_(_4122_, _4133_, _4135_);
  or g_7279_(_3969_, _3971_, _4137_);
  or g_7280_(_3964_, _3966_, _4138_);
  and g_7281_(G11[9], G12[17], _4139_);
  and g_7282_(G11[11], G12[15], _4140_);
  and g_7283_(G11[11], G12[16], _4141_);
  and g_7284_(_3963_, _4140_, _4142_);
  xor g_7285_(_3963_, _4140_, _4143_);
  and g_7286_(_4139_, _4143_, _4144_);
  xor g_7287_(_4139_, _4143_, _4145_);
  or g_7288_(_3989_, _3991_, _4146_);
  and g_7289_(_4145_, _4146_, _4148_);
  xor g_7290_(_4145_, _4146_, _4149_);
  and g_7291_(_4138_, _4149_, _4150_);
  xor g_7292_(_4138_, _4149_, _4151_);
  and g_7293_(_4137_, _4151_, _4152_);
  xor g_7294_(_4137_, _4151_, _4153_);
  and g_7295_(_4135_, _4153_, _4154_);
  xor g_7296_(_4135_, _4153_, _4155_);
  or g_7297_(_4008_, _4010_, _4156_);
  and g_7298_(_4155_, _4156_, _4157_);
  xor g_7299_(_4155_, _4156_, _4159_);
  and g_7300_(_4115_, _4159_, _4160_);
  xor g_7301_(_4115_, _4159_, _4161_);
  or g_7302_(_4054_, _4056_, _4162_);
  or g_7303_(_4002_, _4004_, _4163_);
  and g_7304_(G11[12], G12[14], _4164_);
  and g_7305_(G12[12], G11[14], _4165_);
  and g_7306_(G12[13], G11[14], _4166_);
  and g_7307_(_3988_, _4165_, _4167_);
  xor g_7308_(_3988_, _4165_, _4168_);
  and g_7309_(_4164_, _4168_, _4170_);
  xor g_7310_(_4164_, _4168_, _4171_);
  or g_7311_(_3998_, _4000_, _4172_);
  and g_7312_(G12[11], G11[15], _4173_);
  and g_7313_(G12[9], G11[17], _4174_);
  and g_7314_(G12[10], G11[17], _4175_);
  and g_7315_(_3997_, _4174_, _4176_);
  xor g_7316_(_3997_, _4174_, _4177_);
  and g_7317_(_4173_, _4177_, _4178_);
  xor g_7318_(_4173_, _4177_, _4179_);
  and g_7319_(_4172_, _4179_, _4180_);
  xor g_7320_(_4172_, _4179_, _4181_);
  and g_7321_(_4171_, _4181_, _4182_);
  xor g_7322_(_4171_, _4181_, _4183_);
  or g_7323_(_4023_, _4025_, _4184_);
  and g_7324_(_4183_, _4184_, _4185_);
  xor g_7325_(_4183_, _4184_, _4186_);
  and g_7326_(_4163_, _4186_, _4187_);
  xor g_7327_(_4163_, _4186_, _4188_);
  or g_7328_(_4050_, _4052_, _4189_);
  or g_7329_(_4018_, _4020_, _4191_);
  and g_7330_(G12[8], G11[18], _4192_);
  and g_7331_(G12[6], G11[20], _4193_);
  and g_7332_(G12[7], G11[20], _4194_);
  and g_7333_(_4017_, _4193_, _4195_);
  xor g_7334_(_4017_, _4193_, _4196_);
  and g_7335_(_4192_, _4196_, _4197_);
  xor g_7336_(_4192_, _4196_, _4198_);
  or g_7337_(_4032_, _4034_, _4199_);
  and g_7338_(_4198_, _4199_, _4200_);
  xor g_7339_(_4198_, _4199_, _4202_);
  and g_7340_(_4191_, _4202_, _4203_);
  xor g_7341_(_4191_, _4202_, _4204_);
  or g_7342_(_4045_, _4047_, _4205_);
  and g_7343_(G12[5], G11[21], _4206_);
  and g_7344_(G12[2], G11[24], _4207_);
  and g_7345_(G12[4], G11[24], _4208_);
  and g_7346_(_3864_, _4207_, _4209_);
  xor g_7347_(_3864_, _4207_, _4210_);
  and g_7348_(_4206_, _4210_, _4211_);
  xor g_7349_(_4206_, _4210_, _4213_);
  or g_7350_(_4041_, _4043_, _4214_);
  and g_7351_(G12[1], G11[25], _4215_);
  and g_7352_(G12[0], G11[26], _4216_);
  and g_7353_(G12[3], G11[26], _4217_);
  and g_7354_(_3715_, _4217_, _4218_);
  xor g_7355_(_3716_, _4216_, _4219_);
  and g_7356_(_4215_, _4219_, _4220_);
  xor g_7357_(_4215_, _4219_, _4221_);
  and g_7358_(_4214_, _4221_, _4222_);
  xor g_7359_(_4214_, _4221_, _4224_);
  and g_7360_(_4213_, _4224_, _4225_);
  xor g_7361_(_4213_, _4224_, _4226_);
  and g_7362_(_4205_, _4226_, _4227_);
  xor g_7363_(_4205_, _4226_, _4228_);
  and g_7364_(_4204_, _4228_, _4229_);
  xor g_7365_(_4204_, _4228_, _4230_);
  and g_7366_(_4189_, _4230_, _4231_);
  xor g_7367_(_4189_, _4230_, _4232_);
  and g_7368_(_4188_, _4232_, _4233_);
  xor g_7369_(_4188_, _4232_, _4235_);
  and g_7370_(_4162_, _4235_, _4236_);
  xor g_7371_(_4162_, _4235_, _4237_);
  and g_7372_(_4161_, _4237_, _4238_);
  xor g_7373_(_4161_, _4237_, _4239_);
  and g_7374_(_4113_, _4239_, _4240_);
  xor g_7375_(_4113_, _4239_, _4241_);
  and g_7376_(_4112_, _4241_, _4242_);
  xor g_7377_(_4112_, _4241_, _4243_);
  and g_7378_(_4079_, _4243_, _4244_);
  xor g_7379_(_4079_, _4243_, _4246_);
  and g_7380_(_4078_, _4246_, _4247_);
  xor g_7381_(_4078_, _4246_, _4248_);
  and g_7382_(_4077_, _4248_, _4249_);
  xor g_7383_(_4077_, _4248_, _4250_);
  and g_7384_(_4072_, _4250_, _4251_);
  xor g_7385_(_4072_, _4250_, _4252_);
  or g_7386_(_4074_, _4076_, _4253_);
  and g_7387_(_4252_, _4253_, _4254_);
  xor g_7388_(_4252_, _4253_, G14[26]);
  or g_7389_(_4251_, _4254_, _4256_);
  or g_7390_(_4244_, _4247_, _4257_);
  or g_7391_(_4108_, _4111_, _4258_);
  or g_7392_(_4240_, _4242_, _4259_);
  and g_7393_(G11[0], G12[27], _4260_);
  or g_7394_(_4096_, _4098_, _4261_);
  or g_7395_(_4090_, _4093_, _4262_);
  or g_7396_(_4085_, _4087_, _4263_);
  and g_7397_(G11[1], G12[26], _4264_);
  and g_7398_(G11[3], G12[24], _4265_);
  and g_7399_(G11[3], G12[25], _4267_);
  and g_7400_(_4084_, _4265_, _4268_);
  xor g_7401_(_4084_, _4265_, _4269_);
  and g_7402_(_4264_, _4269_, _4270_);
  xor g_7403_(_4264_, _4269_, _4271_);
  or g_7404_(_4119_, _4121_, _4272_);
  and g_7405_(_4271_, _4272_, _4273_);
  xor g_7406_(_4271_, _4272_, _4274_);
  and g_7407_(_4263_, _4274_, _4275_);
  xor g_7408_(_4263_, _4274_, _4276_);
  or g_7409_(_4132_, _4134_, _4278_);
  and g_7410_(_4276_, _4278_, _4279_);
  xor g_7411_(_4276_, _4278_, _4280_);
  and g_7412_(_4262_, _4280_, _4281_);
  xor g_7413_(_4262_, _4280_, _4282_);
  and g_7414_(_4261_, _4282_, _4283_);
  xor g_7415_(_4261_, _4282_, _4284_);
  and g_7416_(_4260_, _4284_, _4285_);
  xor g_7417_(_4260_, _4284_, _4286_);
  or g_7418_(_4157_, _4160_, _4287_);
  and g_7419_(_4286_, _4287_, _4289_);
  xor g_7420_(_4286_, _4287_, _4290_);
  and g_7421_(_4104_, _4290_, _4291_);
  xor g_7422_(_4104_, _4290_, _4292_);
  or g_7423_(_4236_, _4238_, _4293_);
  or g_7424_(_4152_, _4154_, _4294_);
  and g_7425_(G11[4], G12[23], _4295_);
  and g_7426_(G11[6], G12[21], _4296_);
  and g_7427_(G11[6], G12[22], _4297_);
  and g_7428_(_4118_, _4296_, _4298_);
  xor g_7429_(_4118_, _4296_, _4300_);
  and g_7430_(_4295_, _4300_, _4301_);
  xor g_7431_(_4295_, _4300_, _4302_);
  or g_7432_(_4128_, _4130_, _4303_);
  and g_7433_(G11[7], G12[20], _4304_);
  and g_7434_(G11[9], G12[18], _4305_);
  and g_7435_(G11[9], G12[19], _4306_);
  and g_7436_(_4127_, _4305_, _4307_);
  xor g_7437_(_4127_, _4305_, _4308_);
  and g_7438_(_4304_, _4308_, _4309_);
  xor g_7439_(_4304_, _4308_, _4311_);
  and g_7440_(_4303_, _4311_, _4312_);
  xor g_7441_(_4303_, _4311_, _4313_);
  and g_7442_(_4302_, _4313_, _4314_);
  xor g_7443_(_4302_, _4313_, _4315_);
  or g_7444_(_4148_, _4150_, _4316_);
  or g_7445_(_4142_, _4144_, _4317_);
  and g_7446_(G11[10], G12[17], _4318_);
  and g_7447_(G11[12], G12[15], _4319_);
  and g_7448_(G11[12], G12[16], _4320_);
  and g_7449_(_4141_, _4319_, _4322_);
  xor g_7450_(_4141_, _4319_, _4323_);
  and g_7451_(_4318_, _4323_, _4324_);
  xor g_7452_(_4318_, _4323_, _4325_);
  or g_7453_(_4167_, _4170_, _4326_);
  and g_7454_(_4325_, _4326_, _4327_);
  xor g_7455_(_4325_, _4326_, _4328_);
  and g_7456_(_4317_, _4328_, _4329_);
  xor g_7457_(_4317_, _4328_, _4330_);
  and g_7458_(_4316_, _4330_, _4331_);
  xor g_7459_(_4316_, _4330_, _4333_);
  and g_7460_(_4315_, _4333_, _4334_);
  xor g_7461_(_4315_, _4333_, _4335_);
  or g_7462_(_4185_, _4187_, _4336_);
  and g_7463_(_4335_, _4336_, _4337_);
  xor g_7464_(_4335_, _4336_, _4338_);
  and g_7465_(_4294_, _4338_, _4339_);
  xor g_7466_(_4294_, _4338_, _4340_);
  or g_7467_(_4231_, _4233_, _4341_);
  or g_7468_(_4180_, _4182_, _4342_);
  and g_7469_(G11[13], G12[14], _4344_);
  and g_7470_(G12[12], G11[15], _4345_);
  and g_7471_(G12[13], G11[15], _4346_);
  and g_7472_(_4166_, _4345_, _4347_);
  xor g_7473_(_4166_, _4345_, _4348_);
  and g_7474_(_4344_, _4348_, _4349_);
  xor g_7475_(_4344_, _4348_, _4350_);
  or g_7476_(_4176_, _4178_, _4351_);
  and g_7477_(G12[11], G11[16], _4352_);
  and g_7478_(G12[9], G11[18], _4353_);
  and g_7479_(G12[10], G11[18], _4355_);
  and g_7480_(_4175_, _4353_, _4356_);
  xor g_7481_(_4175_, _4353_, _4357_);
  and g_7482_(_4352_, _4357_, _4358_);
  xor g_7483_(_4352_, _4357_, _4359_);
  and g_7484_(_4351_, _4359_, _4360_);
  xor g_7485_(_4351_, _4359_, _4361_);
  and g_7486_(_4350_, _4361_, _4362_);
  xor g_7487_(_4350_, _4361_, _4363_);
  or g_7488_(_4200_, _4203_, _4364_);
  and g_7489_(_4363_, _4364_, _4366_);
  xor g_7490_(_4363_, _4364_, _4367_);
  and g_7491_(_4342_, _4367_, _4368_);
  xor g_7492_(_4342_, _4367_, _4369_);
  or g_7493_(_4227_, _4229_, _4370_);
  or g_7494_(_4195_, _4197_, _4371_);
  and g_7495_(G12[8], G11[19], _4372_);
  and g_7496_(G12[6], G11[21], _4373_);
  and g_7497_(G12[7], G11[21], _4374_);
  and g_7498_(_4194_, _4373_, _4375_);
  xor g_7499_(_4194_, _4373_, _4377_);
  and g_7500_(_4372_, _4377_, _4378_);
  xor g_7501_(_4372_, _4377_, _4379_);
  or g_7502_(_4209_, _4211_, _4380_);
  and g_7503_(_4379_, _4380_, _4381_);
  xor g_7504_(_4379_, _4380_, _4382_);
  and g_7505_(_4371_, _4382_, _4383_);
  xor g_7506_(_4371_, _4382_, _4384_);
  or g_7507_(_4222_, _4225_, _4385_);
  and g_7508_(G12[5], G11[22], _4386_);
  and g_7509_(G12[2], G11[25], _4388_);
  and g_7510_(G12[4], G11[25], _4389_);
  and g_7511_(_4031_, _4388_, _4390_);
  xor g_7512_(_4031_, _4388_, _4391_);
  and g_7513_(_4386_, _4391_, _4392_);
  xor g_7514_(_4386_, _4391_, _4393_);
  or g_7515_(_4218_, _4220_, _4394_);
  and g_7516_(G12[1], G11[26], _4395_);
  and g_7517_(G12[0], G11[27], _4396_);
  and g_7518_(G12[3], G11[27], _4397_);
  and g_7519_(_3871_, _4397_, _4399_);
  xor g_7520_(_3872_, _4396_, _4400_);
  and g_7521_(_4395_, _4400_, _4401_);
  xor g_7522_(_4395_, _4400_, _4402_);
  and g_7523_(_4394_, _4402_, _4403_);
  xor g_7524_(_4394_, _4402_, _4404_);
  and g_7525_(_4393_, _4404_, _4405_);
  xor g_7526_(_4393_, _4404_, _4406_);
  and g_7527_(_4385_, _4406_, _4407_);
  xor g_7528_(_4385_, _4406_, _4408_);
  and g_7529_(_4384_, _4408_, _4410_);
  xor g_7530_(_4384_, _4408_, _4411_);
  and g_7531_(_4370_, _4411_, _4412_);
  xor g_7532_(_4370_, _4411_, _4413_);
  and g_7533_(_4369_, _4413_, _4414_);
  xor g_7534_(_4369_, _4413_, _4415_);
  and g_7535_(_4341_, _4415_, _4416_);
  xor g_7536_(_4341_, _4415_, _4417_);
  and g_7537_(_4340_, _4417_, _4418_);
  xor g_7538_(_4340_, _4417_, _4419_);
  and g_7539_(_4293_, _4419_, _4421_);
  xor g_7540_(_4293_, _4419_, _4422_);
  and g_7541_(_4292_, _4422_, _4423_);
  xor g_7542_(_4292_, _4422_, _4424_);
  and g_7543_(_4259_, _4424_, _4425_);
  xor g_7544_(_4259_, _4424_, _4426_);
  and g_7545_(_4258_, _4426_, _4427_);
  xor g_7546_(_4258_, _4426_, _4428_);
  and g_7547_(_4257_, _4428_, _4429_);
  xor g_7548_(_4257_, _4428_, _4430_);
  and g_7549_(_4249_, _4430_, _4432_);
  xor g_7550_(_4249_, _4430_, _4433_);
  and g_7551_(_4256_, _4433_, _4434_);
  xor g_7552_(_4256_, _4433_, G14[27]);
  or g_7553_(_4425_, _4427_, _4435_);
  or g_7554_(_4289_, _4291_, _4436_);
  or g_7555_(_4421_, _4423_, _4437_);
  or g_7556_(_4283_, _4285_, _4438_);
  and g_7557_(G11[0], G12[28], _4439_);
  and g_7558_(G11[1], G12[27], _4440_);
  and g_7559_(G11[1], G12[28], _4442_);
  and g_7560_(_4260_, _4442_, _4443_);
  xor g_7561_(_4439_, _4440_, _4444_);
  or g_7562_(_4279_, _4281_, _4445_);
  or g_7563_(_4273_, _4275_, _4446_);
  or g_7564_(_4268_, _4270_, _4447_);
  and g_7565_(G11[2], G12[26], _4448_);
  and g_7566_(G11[4], G12[24], _4449_);
  and g_7567_(G11[4], G12[25], _4450_);
  and g_7568_(_4267_, _4449_, _4451_);
  xor g_7569_(_4267_, _4449_, _4453_);
  and g_7570_(_4448_, _4453_, _4454_);
  xor g_7571_(_4448_, _4453_, _4455_);
  or g_7572_(_4298_, _4301_, _4456_);
  and g_7573_(_4455_, _4456_, _4457_);
  xor g_7574_(_4455_, _4456_, _4458_);
  and g_7575_(_4447_, _4458_, _4459_);
  xor g_7576_(_4447_, _4458_, _4460_);
  or g_7577_(_4312_, _4314_, _4461_);
  and g_7578_(_4460_, _4461_, _4462_);
  xor g_7579_(_4460_, _4461_, _4464_);
  and g_7580_(_4446_, _4464_, _4465_);
  xor g_7581_(_4446_, _4464_, _4466_);
  and g_7582_(_4445_, _4466_, _4467_);
  xor g_7583_(_4445_, _4466_, _4468_);
  and g_7584_(_4444_, _4468_, _4469_);
  xor g_7585_(_4444_, _4468_, _4470_);
  or g_7586_(_4337_, _4339_, _4471_);
  and g_7587_(_4470_, _4471_, _4472_);
  xor g_7588_(_4470_, _4471_, _4473_);
  and g_7589_(_4438_, _4473_, _4475_);
  xor g_7590_(_4438_, _4473_, _4476_);
  or g_7591_(_4416_, _4418_, _4477_);
  or g_7592_(_4331_, _4334_, _4478_);
  and g_7593_(G11[5], G12[23], _4479_);
  and g_7594_(G11[7], G12[21], _4480_);
  and g_7595_(G11[7], G12[22], _4481_);
  and g_7596_(_4297_, _4480_, _4482_);
  xor g_7597_(_4297_, _4480_, _4483_);
  and g_7598_(_4479_, _4483_, _4484_);
  xor g_7599_(_4479_, _4483_, _4486_);
  or g_7600_(_4307_, _4309_, _4487_);
  and g_7601_(G11[8], G12[20], _4488_);
  and g_7602_(G11[10], G12[18], _4489_);
  and g_7603_(G11[10], G12[19], _4490_);
  and g_7604_(_4306_, _4489_, _4491_);
  xor g_7605_(_4306_, _4489_, _4492_);
  and g_7606_(_4488_, _4492_, _4493_);
  xor g_7607_(_4488_, _4492_, _4494_);
  and g_7608_(_4487_, _4494_, _4495_);
  xor g_7609_(_4487_, _4494_, _4497_);
  and g_7610_(_4486_, _4497_, _4498_);
  xor g_7611_(_4486_, _4497_, _4499_);
  or g_7612_(_4327_, _4329_, _4500_);
  or g_7613_(_4322_, _4324_, _4501_);
  and g_7614_(G11[11], G12[17], _4502_);
  and g_7615_(G11[13], G12[15], _4503_);
  and g_7616_(G11[13], G12[16], _4504_);
  and g_7617_(_4320_, _4503_, _4505_);
  xor g_7618_(_4320_, _4503_, _4506_);
  and g_7619_(_4502_, _4506_, _4508_);
  xor g_7620_(_4502_, _4506_, _4509_);
  or g_7621_(_4347_, _4349_, _4510_);
  and g_7622_(_4509_, _4510_, _4511_);
  xor g_7623_(_4509_, _4510_, _4512_);
  and g_7624_(_4501_, _4512_, _4513_);
  xor g_7625_(_4501_, _4512_, _4514_);
  and g_7626_(_4500_, _4514_, _4515_);
  xor g_7627_(_4500_, _4514_, _4516_);
  and g_7628_(_4499_, _4516_, _4517_);
  xor g_7629_(_4499_, _4516_, _4519_);
  or g_7630_(_4366_, _4368_, _4520_);
  and g_7631_(_4519_, _4520_, _4521_);
  xor g_7632_(_4519_, _4520_, _4522_);
  and g_7633_(_4478_, _4522_, _4523_);
  xor g_7634_(_4478_, _4522_, _4524_);
  or g_7635_(_4412_, _4414_, _4525_);
  or g_7636_(_4360_, _4362_, _4526_);
  and g_7637_(G11[14], G12[14], _4527_);
  and g_7638_(G12[12], G11[16], _4528_);
  and g_7639_(G12[13], G11[16], _4530_);
  and g_7640_(_4346_, _4528_, _4531_);
  xor g_7641_(_4346_, _4528_, _4532_);
  and g_7642_(_4527_, _4532_, _4533_);
  xor g_7643_(_4527_, _4532_, _4534_);
  or g_7644_(_4356_, _4358_, _4535_);
  and g_7645_(G12[11], G11[17], _4536_);
  and g_7646_(G12[9], G11[19], _4537_);
  and g_7647_(G12[10], G11[19], _4538_);
  and g_7648_(_4355_, _4537_, _4539_);
  xor g_7649_(_4355_, _4537_, _4541_);
  and g_7650_(_4536_, _4541_, _4542_);
  xor g_7651_(_4536_, _4541_, _4543_);
  and g_7652_(_4535_, _4543_, _4544_);
  xor g_7653_(_4535_, _4543_, _4545_);
  and g_7654_(_4534_, _4545_, _4546_);
  xor g_7655_(_4534_, _4545_, _4547_);
  or g_7656_(_4381_, _4383_, _4548_);
  and g_7657_(_4547_, _4548_, _4549_);
  xor g_7658_(_4547_, _4548_, _4550_);
  and g_7659_(_4526_, _4550_, _4552_);
  xor g_7660_(_4526_, _4550_, _4553_);
  or g_7661_(_4407_, _4410_, _4554_);
  or g_7662_(_4375_, _4378_, _4555_);
  and g_7663_(G12[8], G11[20], _4556_);
  and g_7664_(G12[6], G11[22], _4557_);
  and g_7665_(G12[7], G11[22], _4558_);
  and g_7666_(_4374_, _4557_, _4559_);
  xor g_7667_(_4374_, _4557_, _4560_);
  and g_7668_(_4556_, _4560_, _4561_);
  xor g_7669_(_4556_, _4560_, _4563_);
  or g_7670_(_4390_, _4392_, _4564_);
  and g_7671_(_4563_, _4564_, _4565_);
  xor g_7672_(_4563_, _4564_, _4566_);
  and g_7673_(_4555_, _4566_, _4567_);
  xor g_7674_(_4555_, _4566_, _4568_);
  or g_7675_(_4403_, _4405_, _4569_);
  and g_7676_(G12[5], G11[23], _4570_);
  and g_7677_(G12[2], G11[26], _4571_);
  and g_7678_(G12[4], G11[26], _4572_);
  and g_7679_(_4207_, _4572_, _4574_);
  xor g_7680_(_4208_, _4571_, _4575_);
  and g_7681_(_4570_, _4575_, _4576_);
  xor g_7682_(_4570_, _4575_, _4577_);
  or g_7683_(_4399_, _4401_, _4578_);
  and g_7684_(G12[1], G11[27], _4579_);
  and g_7685_(G12[0], G11[28], _4580_);
  and g_7686_(G12[3], G11[28], _4581_);
  and g_7687_(_4039_, _4581_, _4582_);
  xor g_7688_(_4040_, _4580_, _4583_);
  and g_7689_(_4579_, _4583_, _4585_);
  xor g_7690_(_4579_, _4583_, _4586_);
  and g_7691_(_4578_, _4586_, _4587_);
  xor g_7692_(_4578_, _4586_, _4588_);
  and g_7693_(_4577_, _4588_, _4589_);
  xor g_7694_(_4577_, _4588_, _4590_);
  and g_7695_(_4569_, _4590_, _4591_);
  xor g_7696_(_4569_, _4590_, _4592_);
  and g_7697_(_4568_, _4592_, _4593_);
  xor g_7698_(_4568_, _4592_, _4594_);
  and g_7699_(_4554_, _4594_, _4596_);
  xor g_7700_(_4554_, _4594_, _4597_);
  and g_7701_(_4553_, _4597_, _4598_);
  xor g_7702_(_4553_, _4597_, _4599_);
  and g_7703_(_4525_, _4599_, _4600_);
  xor g_7704_(_4525_, _4599_, _4601_);
  and g_7705_(_4524_, _4601_, _4602_);
  xor g_7706_(_4524_, _4601_, _4603_);
  and g_7707_(_4477_, _4603_, _4604_);
  xor g_7708_(_4477_, _4603_, _4605_);
  and g_7709_(_4476_, _4605_, _4607_);
  xor g_7710_(_4476_, _4605_, _4608_);
  and g_7711_(_4437_, _4608_, _4609_);
  xor g_7712_(_4437_, _4608_, _4610_);
  and g_7713_(_4436_, _4610_, _4611_);
  xor g_7714_(_4436_, _4610_, _4612_);
  and g_7715_(_4435_, _4612_, _4613_);
  xor g_7716_(_4435_, _4612_, _4614_);
  and g_7717_(_4429_, _4614_, _4615_);
  xor g_7718_(_4429_, _4614_, _4616_);
  or g_7719_(_4432_, _4434_, _4618_);
  and g_7720_(_4616_, _4618_, _4619_);
  xor g_7721_(_4616_, _4618_, G14[28]);
  or g_7722_(_4615_, _4619_, _4620_);
  or g_7723_(_4609_, _4611_, _4621_);
  or g_7724_(_4472_, _4475_, _4622_);
  or g_7725_(_4604_, _4607_, _4623_);
  or g_7726_(_4467_, _4469_, _4624_);
  and g_7727_(G11[0], G12[29], _4625_);
  and g_7728_(G11[2], G12[27], _4626_);
  and g_7729_(G11[2], G12[28], _4628_);
  and g_7730_(_4442_, _4626_, _4629_);
  xor g_7731_(_4442_, _4626_, _4630_);
  and g_7732_(_4625_, _4630_, _4631_);
  xor g_7733_(_4625_, _4630_, _4632_);
  and g_7734_(_4443_, _4632_, _4633_);
  not g_7735_(_4633_, _4634_);
  xor g_7736_(_4443_, _4632_, _4635_);
  or g_7737_(_4462_, _4465_, _4636_);
  or g_7738_(_4457_, _4459_, _4637_);
  or g_7739_(_4451_, _4454_, _4639_);
  and g_7740_(G11[3], G12[26], _4640_);
  and g_7741_(G11[5], G12[24], _4641_);
  and g_7742_(G11[5], G12[25], _4642_);
  and g_7743_(_4450_, _4641_, _4643_);
  xor g_7744_(_4450_, _4641_, _4644_);
  and g_7745_(_4640_, _4644_, _4645_);
  xor g_7746_(_4640_, _4644_, _4646_);
  or g_7747_(_4482_, _4484_, _4647_);
  and g_7748_(_4646_, _4647_, _4648_);
  xor g_7749_(_4646_, _4647_, _4649_);
  and g_7750_(_4639_, _4649_, _4650_);
  xor g_7751_(_4639_, _4649_, _4651_);
  or g_7752_(_4495_, _4498_, _4652_);
  and g_7753_(_4651_, _4652_, _4653_);
  xor g_7754_(_4651_, _4652_, _4654_);
  and g_7755_(_4637_, _4654_, _4655_);
  xor g_7756_(_4637_, _4654_, _4656_);
  and g_7757_(_4636_, _4656_, _4657_);
  xor g_7758_(_4636_, _4656_, _4658_);
  and g_7759_(_4635_, _4658_, _4660_);
  xor g_7760_(_4635_, _4658_, _4661_);
  or g_7761_(_4521_, _4523_, _4662_);
  and g_7762_(_4661_, _4662_, _4663_);
  xor g_7763_(_4661_, _4662_, _4664_);
  and g_7764_(_4624_, _4664_, _4665_);
  xor g_7765_(_4624_, _4664_, _4666_);
  or g_7766_(_4600_, _4602_, _4667_);
  or g_7767_(_4515_, _4517_, _4668_);
  and g_7768_(G11[6], G12[23], _4669_);
  and g_7769_(G11[8], G12[21], _4671_);
  and g_7770_(G11[8], G12[22], _4672_);
  and g_7771_(_4481_, _4671_, _4673_);
  xor g_7772_(_4481_, _4671_, _4674_);
  and g_7773_(_4669_, _4674_, _4675_);
  xor g_7774_(_4669_, _4674_, _4676_);
  or g_7775_(_4491_, _4493_, _4677_);
  and g_7776_(G11[9], G12[20], _4678_);
  and g_7777_(G11[11], G12[18], _4679_);
  and g_7778_(G11[11], G12[19], _4680_);
  and g_7779_(_4490_, _4679_, _4682_);
  xor g_7780_(_4490_, _4679_, _4683_);
  and g_7781_(_4678_, _4683_, _4684_);
  xor g_7782_(_4678_, _4683_, _4685_);
  and g_7783_(_4677_, _4685_, _4686_);
  xor g_7784_(_4677_, _4685_, _4687_);
  and g_7785_(_4676_, _4687_, _4688_);
  xor g_7786_(_4676_, _4687_, _4689_);
  or g_7787_(_4511_, _4513_, _4690_);
  or g_7788_(_4505_, _4508_, _4691_);
  and g_7789_(G11[12], G12[17], _4693_);
  and g_7790_(G11[14], G12[15], _4694_);
  and g_7791_(G11[14], G12[16], _4695_);
  and g_7792_(_4504_, _4694_, _4696_);
  xor g_7793_(_4504_, _4694_, _4697_);
  and g_7794_(_4693_, _4697_, _4698_);
  xor g_7795_(_4693_, _4697_, _4699_);
  or g_7796_(_4531_, _4533_, _4700_);
  and g_7797_(_4699_, _4700_, _4701_);
  xor g_7798_(_4699_, _4700_, _4702_);
  and g_7799_(_4691_, _4702_, _4704_);
  xor g_7800_(_4691_, _4702_, _4705_);
  and g_7801_(_4690_, _4705_, _4706_);
  xor g_7802_(_4690_, _4705_, _4707_);
  and g_7803_(_4689_, _4707_, _4708_);
  xor g_7804_(_4689_, _4707_, _4709_);
  or g_7805_(_4549_, _4552_, _4710_);
  and g_7806_(_4709_, _4710_, _4711_);
  xor g_7807_(_4709_, _4710_, _4712_);
  and g_7808_(_4668_, _4712_, _4713_);
  xor g_7809_(_4668_, _4712_, _4715_);
  or g_7810_(_4596_, _4598_, _4716_);
  or g_7811_(_4544_, _4546_, _4717_);
  and g_7812_(G12[14], G11[15], _4718_);
  and g_7813_(G12[12], G11[17], _4719_);
  and g_7814_(G12[13], G11[17], _4720_);
  and g_7815_(_4530_, _4719_, _4721_);
  xor g_7816_(_4530_, _4719_, _4722_);
  and g_7817_(_4718_, _4722_, _4723_);
  xor g_7818_(_4718_, _4722_, _4724_);
  or g_7819_(_4539_, _4542_, _4726_);
  and g_7820_(G12[11], G11[18], _4727_);
  and g_7821_(G12[9], G11[20], _4728_);
  and g_7822_(G12[10], G11[20], _4729_);
  and g_7823_(_4538_, _4728_, _4730_);
  xor g_7824_(_4538_, _4728_, _4731_);
  and g_7825_(_4727_, _4731_, _4732_);
  xor g_7826_(_4727_, _4731_, _4733_);
  and g_7827_(_4726_, _4733_, _4734_);
  xor g_7828_(_4726_, _4733_, _4735_);
  and g_7829_(_4724_, _4735_, _4737_);
  xor g_7830_(_4724_, _4735_, _4738_);
  or g_7831_(_4565_, _4567_, _4739_);
  and g_7832_(_4738_, _4739_, _4740_);
  xor g_7833_(_4738_, _4739_, _4741_);
  and g_7834_(_4717_, _4741_, _4742_);
  xor g_7835_(_4717_, _4741_, _4743_);
  or g_7836_(_4591_, _4593_, _4744_);
  or g_7837_(_4559_, _4561_, _4745_);
  and g_7838_(G12[8], G11[21], _4746_);
  and g_7839_(G12[6], G11[23], _4748_);
  and g_7840_(G12[7], G11[23], _4749_);
  and g_7841_(_4558_, _4748_, _4750_);
  xor g_7842_(_4558_, _4748_, _4751_);
  and g_7843_(_4746_, _4751_, _4752_);
  xor g_7844_(_4746_, _4751_, _4753_);
  or g_7845_(_4574_, _4576_, _4754_);
  and g_7846_(_4753_, _4754_, _4755_);
  xor g_7847_(_4753_, _4754_, _4756_);
  and g_7848_(_4745_, _4756_, _4757_);
  xor g_7849_(_4745_, _4756_, _4759_);
  or g_7850_(_4587_, _4589_, _4760_);
  and g_7851_(G12[5], G11[24], _4761_);
  and g_7852_(G12[2], G11[27], _4762_);
  and g_7853_(G12[4], G11[27], _4763_);
  and g_7854_(_4388_, _4763_, _4764_);
  xor g_7855_(_4389_, _4762_, _4765_);
  and g_7856_(_4761_, _4765_, _4766_);
  xor g_7857_(_4761_, _4765_, _4767_);
  or g_7858_(_4582_, _4585_, _4768_);
  and g_7859_(G12[1], G11[28], _4770_);
  and g_7860_(G12[0], G11[29], _4771_);
  and g_7861_(_4217_, _4771_, _4772_);
  xor g_7862_(_4217_, _4771_, _4773_);
  and g_7863_(_4770_, _4773_, _4774_);
  xor g_7864_(_4770_, _4773_, _4775_);
  and g_7865_(_4768_, _4775_, _4776_);
  xor g_7866_(_4768_, _4775_, _4777_);
  and g_7867_(_4767_, _4777_, _4778_);
  xor g_7868_(_4767_, _4777_, _4779_);
  and g_7869_(_4760_, _4779_, _4781_);
  xor g_7870_(_4760_, _4779_, _4782_);
  and g_7871_(_4759_, _4782_, _4783_);
  xor g_7872_(_4759_, _4782_, _4784_);
  and g_7873_(_4744_, _4784_, _4785_);
  xor g_7874_(_4744_, _4784_, _4786_);
  and g_7875_(_4743_, _4786_, _4787_);
  xor g_7876_(_4743_, _4786_, _4788_);
  and g_7877_(_4716_, _4788_, _4789_);
  xor g_7878_(_4716_, _4788_, _4790_);
  and g_7879_(_4715_, _4790_, _4792_);
  xor g_7880_(_4715_, _4790_, _4793_);
  and g_7881_(_4667_, _4793_, _4794_);
  xor g_7882_(_4667_, _4793_, _4795_);
  and g_7883_(_4666_, _4795_, _4796_);
  xor g_7884_(_4666_, _4795_, _4797_);
  and g_7885_(_4623_, _4797_, _4798_);
  xor g_7886_(_4623_, _4797_, _4799_);
  and g_7887_(_4622_, _4799_, _4800_);
  xor g_7888_(_4622_, _4799_, _4801_);
  and g_7889_(_4621_, _4801_, _4803_);
  xor g_7890_(_4621_, _4801_, _4804_);
  and g_7891_(_4613_, _4804_, _4805_);
  xor g_7892_(_4613_, _4804_, _4806_);
  and g_7893_(_4620_, _4806_, _4807_);
  xor g_7894_(_4620_, _4806_, G14[29]);
  or g_7895_(_4798_, _4800_, _4808_);
  or g_7896_(_4663_, _4665_, _4809_);
  or g_7897_(_4794_, _4796_, _4810_);
  or g_7898_(_4657_, _4660_, _4811_);
  not g_7899_(_4811_, _4813_);
  and g_7900_(G11[0], G12[30], _4814_);
  or g_7901_(_4629_, _4631_, _4815_);
  and g_7902_(G11[1], G12[29], _4816_);
  and g_7903_(G11[3], G12[27], _4817_);
  and g_7904_(G11[3], G12[28], _4818_);
  and g_7905_(_4626_, _4818_, _4819_);
  xor g_7906_(_4628_, _4817_, _4820_);
  and g_7907_(_4816_, _4820_, _4821_);
  xor g_7908_(_4816_, _4820_, _4822_);
  and g_7909_(_4815_, _4822_, _4824_);
  xor g_7910_(_4815_, _4822_, _4825_);
  and g_7911_(_4814_, _4825_, _4826_);
  xor g_7912_(_4814_, _4825_, _4827_);
  and g_7913_(_4633_, _4827_, _4828_);
  xor g_7914_(_4634_, _4827_, _4829_);
  not g_7915_(_4829_, _4830_);
  or g_7916_(_4653_, _4655_, _4831_);
  or g_7917_(_4648_, _4650_, _4832_);
  or g_7918_(_4643_, _4645_, _4833_);
  and g_7919_(G11[4], G12[26], _4835_);
  and g_7920_(G11[6], G12[24], _4836_);
  and g_7921_(G11[6], G12[25], _4837_);
  and g_7922_(_4641_, _4837_, _4838_);
  xor g_7923_(_4642_, _4836_, _4839_);
  and g_7924_(_4835_, _4839_, _4840_);
  xor g_7925_(_4835_, _4839_, _4841_);
  or g_7926_(_4673_, _4675_, _4842_);
  and g_7927_(_4841_, _4842_, _4843_);
  xor g_7928_(_4841_, _4842_, _4844_);
  and g_7929_(_4833_, _4844_, _4846_);
  xor g_7930_(_4833_, _4844_, _4847_);
  or g_7931_(_4686_, _4688_, _4848_);
  and g_7932_(_4847_, _4848_, _4849_);
  xor g_7933_(_4847_, _4848_, _4850_);
  and g_7934_(_4832_, _4850_, _4851_);
  xor g_7935_(_4832_, _4850_, _4852_);
  and g_7936_(_4831_, _4852_, _4853_);
  xor g_7937_(_4831_, _4852_, _4854_);
  and g_7938_(_4830_, _4854_, _4855_);
  xor g_7939_(_4829_, _4854_, _4857_);
  or g_7940_(_4711_, _4713_, _4858_);
  not g_7941_(_4858_, _4859_);
  or g_7942_(_4857_, _4859_, _4860_);
  xor g_7943_(_4857_, _4858_, _4861_);
  or g_7944_(_4813_, _4861_, _4862_);
  xor g_7945_(_4813_, _4861_, _4863_);
  or g_7946_(_4789_, _4792_, _4864_);
  or g_7947_(_4706_, _4708_, _4865_);
  and g_7948_(G11[7], G12[23], _4866_);
  and g_7949_(G11[9], G12[21], _4868_);
  and g_7950_(G11[9], G12[22], _4869_);
  and g_7951_(_4671_, _4869_, _4870_);
  xor g_7952_(_4672_, _4868_, _4871_);
  and g_7953_(_4866_, _4871_, _4872_);
  xor g_7954_(_4866_, _4871_, _4873_);
  or g_7955_(_4682_, _4684_, _4874_);
  and g_7956_(G11[10], G12[20], _4875_);
  and g_7957_(G11[12], G12[18], _4876_);
  and g_7958_(G11[12], G12[19], _4877_);
  and g_7959_(_4679_, _4877_, _4879_);
  xor g_7960_(_4680_, _4876_, _4880_);
  and g_7961_(_4875_, _4880_, _4881_);
  xor g_7962_(_4875_, _4880_, _4882_);
  and g_7963_(_4874_, _4882_, _4883_);
  xor g_7964_(_4874_, _4882_, _4884_);
  and g_7965_(_4873_, _4884_, _4885_);
  xor g_7966_(_4873_, _4884_, _4886_);
  or g_7967_(_4701_, _4704_, _4887_);
  or g_7968_(_4696_, _4698_, _4888_);
  not g_7969_(_4888_, _4890_);
  and g_7970_(G11[13], G12[17], _4891_);
  and g_7971_(G11[15], G12[15], _4892_);
  and g_7972_(G11[15], G12[16], _4893_);
  and g_7973_(_4694_, _4893_, _4894_);
  xor g_7974_(_4695_, _4892_, _4895_);
  and g_7975_(_4891_, _4895_, _4896_);
  xor g_7976_(_4891_, _4895_, _4897_);
  or g_7977_(_4721_, _4723_, _4898_);
  and g_7978_(_4897_, _4898_, _4899_);
  xor g_7979_(_4897_, _4898_, _4901_);
  and g_7980_(_4888_, _4901_, _4902_);
  xor g_7981_(_4890_, _4901_, _4903_);
  not g_7982_(_4903_, _4904_);
  and g_7983_(_4887_, _4904_, _4905_);
  xor g_7984_(_4887_, _4904_, _4906_);
  and g_7985_(_4886_, _4906_, _4907_);
  xor g_7986_(_4886_, _4906_, _4908_);
  or g_7987_(_4740_, _4742_, _4909_);
  and g_7988_(_4908_, _4909_, _4910_);
  xor g_7989_(_4908_, _4909_, _4912_);
  and g_7990_(_4865_, _4912_, _4913_);
  xor g_7991_(_4865_, _4912_, _4914_);
  or g_7992_(_4785_, _4787_, _4915_);
  or g_7993_(_4734_, _4737_, _4916_);
  and g_7994_(G12[14], G11[16], _4917_);
  and g_7995_(G12[12], G11[18], _4918_);
  and g_7996_(G12[13], G11[18], _4919_);
  and g_7997_(_4719_, _4919_, _4920_);
  xor g_7998_(_4720_, _4918_, _4921_);
  and g_7999_(_4917_, _4921_, _4923_);
  xor g_8000_(_4917_, _4921_, _4924_);
  or g_8001_(_4730_, _4732_, _4925_);
  and g_8002_(G12[11], G11[19], _4926_);
  and g_8003_(G12[9], G11[21], _4927_);
  and g_8004_(G12[10], G11[21], _4928_);
  and g_8005_(_4728_, _4928_, _4929_);
  xor g_8006_(_4729_, _4927_, _4930_);
  and g_8007_(_4926_, _4930_, _4931_);
  xor g_8008_(_4926_, _4930_, _4932_);
  and g_8009_(_4925_, _4932_, _4934_);
  xor g_8010_(_4925_, _4932_, _4935_);
  and g_8011_(_4924_, _4935_, _4936_);
  xor g_8012_(_4924_, _4935_, _4937_);
  or g_8013_(_4755_, _4757_, _4938_);
  and g_8014_(_4937_, _4938_, _4939_);
  xor g_8015_(_4937_, _4938_, _4940_);
  and g_8016_(_4916_, _4940_, _4941_);
  xor g_8017_(_4916_, _4940_, _4942_);
  or g_8018_(_4781_, _4783_, _4943_);
  or g_8019_(_4750_, _4752_, _4945_);
  and g_8020_(G12[8], G11[22], _4946_);
  and g_8021_(G12[6], G11[24], _4947_);
  and g_8022_(G12[7], G11[24], _4948_);
  and g_8023_(_4748_, _4948_, _4949_);
  xor g_8024_(_4749_, _4947_, _4950_);
  and g_8025_(_4946_, _4950_, _4951_);
  xor g_8026_(_4946_, _4950_, _4952_);
  or g_8027_(_4764_, _4766_, _4953_);
  and g_8028_(_4952_, _4953_, _4954_);
  xor g_8029_(_4952_, _4953_, _4956_);
  and g_8030_(_4945_, _4956_, _4957_);
  xor g_8031_(_4945_, _4956_, _4958_);
  or g_8032_(_4776_, _4778_, _4959_);
  and g_8033_(G12[5], G11[25], _4960_);
  and g_8034_(G12[2], G11[28], _4961_);
  and g_8035_(_4572_, _4961_, _4962_);
  xor g_8036_(_4572_, _4961_, _4963_);
  and g_8037_(_4960_, _4963_, _4964_);
  xor g_8038_(_4960_, _4963_, _4965_);
  or g_8039_(_4772_, _4774_, _4967_);
  and g_8040_(G12[1], G11[29], _4968_);
  and g_8041_(G12[0], G11[30], _4969_);
  and g_8042_(_4397_, _4969_, _4970_);
  xor g_8043_(_4397_, _4969_, _4971_);
  and g_8044_(_4968_, _4971_, _4972_);
  xor g_8045_(_4968_, _4971_, _4973_);
  and g_8046_(_4967_, _4973_, _4974_);
  xor g_8047_(_4967_, _4973_, _4975_);
  and g_8048_(_4965_, _4975_, _4976_);
  xor g_8049_(_4965_, _4975_, _4978_);
  and g_8050_(_4959_, _4978_, _4979_);
  xor g_8051_(_4959_, _4978_, _4980_);
  and g_8052_(_4958_, _4980_, _4981_);
  xor g_8053_(_4958_, _4980_, _4982_);
  and g_8054_(_4943_, _4982_, _4983_);
  xor g_8055_(_4943_, _4982_, _4984_);
  and g_8056_(_4942_, _4984_, _4985_);
  xor g_8057_(_4942_, _4984_, _4986_);
  and g_8058_(_4915_, _4986_, _4987_);
  xor g_8059_(_4915_, _4986_, _4989_);
  and g_8060_(_4914_, _4989_, _4990_);
  xor g_8061_(_4914_, _4989_, _4991_);
  and g_8062_(_4864_, _4991_, _4992_);
  xor g_8063_(_4864_, _4991_, _4993_);
  and g_8064_(_4863_, _4993_, _4994_);
  xor g_8065_(_4863_, _4993_, _4995_);
  and g_8066_(_4810_, _4995_, _4996_);
  xor g_8067_(_4810_, _4995_, _4997_);
  and g_8068_(_4809_, _4997_, _4998_);
  xor g_8069_(_4809_, _4997_, _5000_);
  and g_8070_(_4808_, _5000_, _5001_);
  xor g_8071_(_4808_, _5000_, _5002_);
  and g_8072_(_4803_, _5002_, _5003_);
  xor g_8073_(_4803_, _5002_, _5004_);
  or g_8074_(_4805_, _4807_, _5005_);
  and g_8075_(_5004_, _5005_, _5006_);
  xor g_8076_(_5004_, _5005_, G14[30]);
  or g_8077_(_5003_, _5006_, _5007_);
  or g_8078_(_4996_, _4998_, _5008_);
  and g_8079_(_4860_, _4862_, _5010_);
  or g_8080_(_4992_, _4994_, _5011_);
  or g_8081_(_4853_, _4855_, _5012_);
  or g_8082_(_4987_, _4990_, _5013_);
  xor g_8083_(_5012_, _5013_, _5014_);
  or g_8084_(_4979_, _4981_, _5015_);
  and g_8085_(G11[8], G12[23], _5016_);
  or g_8086_(_4879_, _4881_, _5017_);
  xor g_8087_(_5016_, _5017_, _5018_);
  and g_8088_(G11[11], G12[20], _5019_);
  or g_8089_(_4920_, _4923_, _5021_);
  and g_8090_(G11[14], G12[17], _5022_);
  and g_8091_(G12[15], G11[16], _5023_);
  xor g_8092_(_4893_, _5023_, _5024_);
  xor g_8093_(_5022_, _5024_, _5025_);
  xor g_8094_(_5021_, _5025_, _5026_);
  and g_8095_(G11[13], G12[18], _5027_);
  xor g_8096_(_4877_, _5027_, _5028_);
  and g_8097_(G11[10], G12[21], _5029_);
  xor g_8098_(_4869_, _5029_, _5030_);
  xor g_8099_(_5028_, _5030_, _5032_);
  xor g_8100_(_5019_, _5032_, _5033_);
  xor g_8101_(_5018_, _5026_, _5034_);
  xor g_8102_(_5033_, _5034_, _5035_);
  or g_8103_(_4894_, _4896_, _5036_);
  or g_8104_(_4899_, _4902_, _5037_);
  xor g_8105_(_5036_, _5037_, _5038_);
  and g_8106_(G12[6], G11[25], _5039_);
  xor g_8107_(_4948_, _5039_, _5040_);
  or g_8108_(_4962_, _4964_, _5041_);
  and g_8109_(G12[8], G11[23], _5043_);
  xor g_8110_(_5040_, _5043_, _5044_);
  xor g_8111_(_5041_, _5044_, _5045_);
  or g_8112_(_4970_, _4972_, _5046_);
  and g_8113_(G12[1], G11[30], _5047_);
  xor g_8114_(_5046_, _5047_, _5048_);
  or g_8115_(_5796_, _5807_, _5049_);
  and g_8116_(G12[0], G11[31], _5050_);
  xor g_8117_(_4581_, _5050_, _5051_);
  and g_8118_(G12[2], G11[29], _5052_);
  xor g_8119_(_4763_, _5052_, _5054_);
  xor g_8120_(_5051_, _5054_, _5055_);
  xor g_8121_(_5049_, _5055_, _5056_);
  xor g_8122_(_5048_, _5056_, _5057_);
  xor g_8123_(_5045_, _5057_, _5058_);
  xor g_8124_(_5035_, _5038_, _5059_);
  xor g_8125_(_5058_, _5059_, _5060_);
  xor g_8126_(_5015_, _5060_, _5061_);
  or g_8127_(_4939_, _4941_, _5062_);
  or g_8128_(_4934_, _4936_, _5063_);
  or g_8129_(_4954_, _4957_, _5065_);
  or g_8130_(_4929_, _4931_, _5066_);
  and g_8131_(G12[11], G11[20], _5067_);
  and g_8132_(G12[9], G11[22], _5068_);
  xor g_8133_(_4928_, _5068_, _5069_);
  xor g_8134_(_5067_, _5069_, _5070_);
  xor g_8135_(_5066_, _5070_, _5071_);
  and g_8136_(G12[14], G11[17], _5072_);
  and g_8137_(G12[12], G11[19], _5073_);
  xor g_8138_(_4919_, _5073_, _5074_);
  xor g_8139_(_5072_, _5074_, _5076_);
  xor g_8140_(_5071_, _5076_, _5077_);
  xor g_8141_(_5065_, _5077_, _5078_);
  xor g_8142_(_5063_, _5078_, _5079_);
  or g_8143_(_4949_, _4951_, _5080_);
  or g_8144_(_4974_, _4976_, _5081_);
  xor g_8145_(_5080_, _5081_, _5082_);
  xor g_8146_(_5079_, _5082_, _5083_);
  xor g_8147_(_5062_, _5083_, _5084_);
  xor g_8148_(_5061_, _5084_, _5085_);
  or g_8149_(_4910_, _4913_, _5087_);
  or g_8150_(_4849_, _4851_, _5088_);
  or g_8151_(_4843_, _4846_, _5089_);
  or g_8152_(_4824_, _4826_, _5090_);
  or g_8153_(_4819_, _4821_, _5091_);
  and g_8154_(G11[1], G12[30], _5092_);
  and g_8155_(G11[2], G12[29], _5093_);
  xor g_8156_(_5092_, _5093_, _5094_);
  and g_8157_(G11[4], G12[27], _5095_);
  xor g_8158_(_4818_, _5095_, _5096_);
  xor g_8159_(_5094_, _5096_, _5098_);
  xor g_8160_(_5091_, _5098_, _5099_);
  and g_8161_(G11[0], G12[31], _5100_);
  xor g_8162_(_5099_, _5100_, _5101_);
  xor g_8163_(_5090_, _5101_, _5102_);
  or g_8164_(_4883_, _4885_, _5103_);
  or g_8165_(_4838_, _4840_, _5104_);
  or g_8166_(_4870_, _4872_, _5105_);
  and g_8167_(G11[5], G12[26], _5106_);
  and g_8168_(G11[7], G12[24], _5107_);
  xor g_8169_(_4837_, _5107_, _5109_);
  xor g_8170_(_5106_, _5109_, _5110_);
  xor g_8171_(_5105_, _5110_, _5111_);
  xor g_8172_(_5104_, _5111_, _5112_);
  xor g_8173_(_5103_, _5112_, _5113_);
  xor g_8174_(_5089_, _5113_, _5114_);
  xor g_8175_(_5102_, _5114_, _5115_);
  xor g_8176_(_5088_, _5115_, _5116_);
  xor g_8177_(_5087_, _5116_, _5117_);
  or g_8178_(_4905_, _4907_, _5118_);
  or g_8179_(_4983_, _4985_, _5120_);
  xor g_8180_(_5118_, _5120_, _5121_);
  xor g_8181_(_5085_, _5121_, _5122_);
  xor g_8182_(_5117_, _5122_, _5123_);
  xor g_8183_(_5014_, _5123_, _5124_);
  xor g_8184_(_5011_, _5124_, _5125_);
  xor g_8185_(_5010_, _5125_, _5126_);
  xor g_8186_(_5008_, _5126_, _5127_);
  xor g_8187_(_4828_, _5001_, _5128_);
  xor g_8188_(_5127_, _5128_, _5129_);
  xor g_8189_(_5007_, _5129_, G14[31]);
  xor g_8190_(_5137_, _5192_, G14[9]);
  not g_8191_(G12[5], _5796_);
  not g_8192_(G11[26], _5807_);
  and g_8193_(G12[1], G11[0], _5818_);
  and g_8194_(G12[0], G11[1], _2886_);
  not g_8195_(_2886_, _2897_);
  and g_8196_(G12[0], G11[0], G14[0]);
  and g_8197_(G11[1], G12[1], _2918_);
  and g_8198_(G14[0], _2918_, _2928_);
  xor g_8199_(_5818_, _2886_, G14[1]);
  and g_8200_(G11[0], G12[2], _2949_);
  and g_8201_(G12[0], G11[2], _2960_);
  and g_8202_(G12[1], G11[2], _2971_);
  and g_8203_(_2886_, _2971_, _2982_);
  xor g_8204_(_2918_, _2960_, _2993_);
  and g_8205_(_2928_, _2993_, _3004_);
  xor g_8206_(_2928_, _2993_, _3015_);
  and g_8207_(_2949_, _3015_, _3026_);
  xor g_8208_(_2949_, _3015_, G14[2]);
  or g_8209_(_3004_, _3026_, _3047_);
  and g_8210_(G11[1], G12[2], _3057_);
  and g_8211_(G12[0], G11[3], _3068_);
  and g_8212_(G11[0], G12[3], _3079_);
  and g_8213_(G12[3], G11[3], _3090_);
  and g_8214_(G14[0], _3090_, _3101_);
  or g_8215_(_3068_, _3079_, _3112_);
  xor g_8216_(_3068_, _3079_, _3123_);
  not g_8217_(_3123_, _3134_);
  and g_8218_(_2897_, _2971_, _3145_);
  xor g_8219_(_3123_, _3145_, _3156_);
  and g_8220_(_3057_, _3156_, _3167_);
  xor g_8221_(_3057_, _3156_, _3178_);
  and g_8222_(_3047_, _3178_, _3188_);
  xor g_8223_(_3047_, _3178_, G14[3]);
  and g_8224_(_2982_, _3134_, _3209_);
  or g_8225_(_3167_, _3209_, _3220_);
  and g_8226_(G11[0], G12[4], _3231_);
  and g_8227_(G11[2], G12[2], _3242_);
  and g_8228_(G11[2], G12[4], _3253_);
  and g_8229_(_2949_, _3253_, _3264_);
  xor g_8230_(_3231_, _3242_, _3275_);
  and g_8231_(G12[1], G11[3], _3286_);
  and g_8232_(G12[0], G11[4], _3297_);
  and g_8233_(G11[1], G12[3], _3308_);
  and g_8234_(G12[3], G11[4], _3318_);
  and g_8235_(_2886_, _3318_, _3329_);
  xor g_8236_(_3297_, _3308_, _3340_);
  and g_8237_(_3286_, _3340_, _3351_);
  xor g_8238_(_3286_, _3340_, _3362_);
  and g_8239_(_2971_, _3112_, _3373_);
  or g_8240_(_3101_, _3373_, _3384_);
  and g_8241_(_3362_, _3384_, _3395_);
  xor g_8242_(_3362_, _3384_, _3406_);
  and g_8243_(_3275_, _3406_, _3417_);
  xor g_8244_(_3275_, _3406_, _3428_);
  and g_8245_(_3220_, _3428_, _3439_);
  xor g_8246_(_3220_, _3428_, _3450_);
  and g_8247_(_3188_, _3450_, _3460_);
  xor g_8248_(_3188_, _3450_, G14[4]);
  or g_8249_(_3395_, _3417_, _3481_);
  and g_8250_(G11[0], G12[5], _3492_);
  and g_8251_(G11[1], G12[4], _3503_);
  and g_8252_(G12[2], G11[3], _3514_);
  and g_8253_(G11[3], G12[4], _3525_);
  and g_8254_(_3057_, _3525_, _3536_);
  xor g_8255_(_3503_, _3514_, _3547_);
  and g_8256_(_3492_, _3547_, _3558_);
  xor g_8257_(_3492_, _3547_, _3569_);
  or g_8258_(_3329_, _3351_, _3580_);
  and g_8259_(G12[1], G11[4], _3591_);
  and g_8260_(G12[0], G11[5], _3601_);
  and g_8261_(G11[2], G12[3], _3612_);
  and g_8262_(G12[3], G11[5], _3623_);
  and g_8263_(_2960_, _3623_, _3634_);
  xor g_8264_(_3601_, _3612_, _3645_);
  and g_8265_(_3591_, _3645_, _3656_);
  xor g_8266_(_3591_, _3645_, _3667_);
  and g_8267_(_3580_, _3667_, _3678_);
  xor g_8268_(_3580_, _3667_, _3689_);
  and g_8269_(_3569_, _3689_, _3700_);
  xor g_8270_(_3569_, _3689_, _3711_);
  and g_8271_(_3481_, _3711_, _3722_);
  xor g_8272_(_3481_, _3711_, _3733_);
  and g_8273_(_3264_, _3733_, _3744_);
  xor g_8274_(_3264_, _3733_, _3754_);
  or g_8275_(_3439_, _3460_, _3765_);
  xor g_8276_(_3754_, _3765_, G14[5]);
  and g_8277_(_3460_, _3754_, _3786_);
  and g_8278_(_3439_, _3754_, _3797_);
  or g_8279_(_3722_, _3744_, _3808_);
  and g_8280_(G11[0], G12[6], _3819_);
  or g_8281_(_3536_, _3558_, _3830_);
  and g_8282_(_3819_, _3830_, _3841_);
  xor g_8283_(_3819_, _3830_, _3852_);
  or g_8284_(_3678_, _3700_, _3863_);
  and g_8285_(G11[1], G12[5], _3874_);
  and g_8286_(G12[2], G11[4], _3885_);
  and g_8287_(G11[4], G12[4], _3896_);
  and g_8288_(_3253_, _3885_, _3907_);
  xor g_8289_(_3253_, _3885_, _3917_);
  and g_8290_(_3874_, _3917_, _3928_);
  xor g_8291_(_3874_, _3917_, _3939_);
  or g_8292_(_3634_, _3656_, _3950_);
  and g_8293_(G12[1], G11[5], _3961_);
  and g_8294_(G12[0], G11[6], _3972_);
  and g_8295_(G12[3], G11[6], _3983_);
  and g_8296_(_3090_, _3972_, _3994_);
  xor g_8297_(_3090_, _3972_, _4005_);
  and g_8298_(_3961_, _4005_, _4016_);
  xor g_8299_(_3961_, _4005_, _4027_);
  and g_8300_(_3950_, _4027_, _4038_);
  xor g_8301_(_3950_, _4027_, _4049_);
  and g_8302_(_3939_, _4049_, _4060_);
  xor g_8303_(_3939_, _4049_, _4071_);
  and g_8304_(_3863_, _4071_, _4081_);
  xor g_8305_(_3863_, _4071_, _4092_);
  and g_8306_(_3852_, _4092_, _4103_);
  xor g_8307_(_3852_, _4092_, _4114_);
  and g_8308_(_3808_, _4114_, _4125_);
  xor g_8309_(_3808_, _4114_, _4136_);
  and g_8310_(_3797_, _4136_, _4147_);
  xor g_8311_(_3797_, _4136_, _4158_);
  and g_8312_(_3786_, _4158_, _4169_);
  xor g_8313_(_3786_, _4158_, G14[6]);
  or g_8314_(_4081_, _4103_, _4190_);
  and g_8315_(G11[0], G12[7], _4201_);
  and g_8316_(G11[1], G12[6], _4212_);
  and g_8317_(G11[1], G12[7], _4223_);
  and g_8318_(_3819_, _4223_, _4234_);
  xor g_8319_(_4201_, _4212_, _4245_);
  or g_8320_(_3907_, _3928_, _4255_);
  and g_8321_(_4245_, _4255_, _4266_);
  xor g_8322_(_4245_, _4255_, _4277_);
  or g_8323_(_4038_, _4060_, _4288_);
  and g_8324_(G11[2], G12[5], _4299_);
  and g_8325_(G12[2], G11[5], _4310_);
  and g_8326_(G12[4], G11[5], _4321_);
  and g_8327_(_3525_, _4310_, _4332_);
  xor g_8328_(_3525_, _4310_, _4343_);
  and g_8329_(_4299_, _4343_, _4354_);
  xor g_8330_(_4299_, _4343_, _4365_);
  or g_8331_(_3994_, _4016_, _4376_);
  and g_8332_(G12[1], G11[6], _4387_);
  and g_8333_(G12[0], G11[7], _4398_);
  and g_8334_(G12[3], G11[7], _4409_);
  and g_8335_(_3318_, _4398_, _4420_);
  xor g_8336_(_3318_, _4398_, _4431_);
  and g_8337_(_4387_, _4431_, _4441_);
  xor g_8338_(_4387_, _4431_, _4452_);
  and g_8339_(_4376_, _4452_, _4463_);
  xor g_8340_(_4376_, _4452_, _4474_);
  and g_8341_(_4365_, _4474_, _4485_);
  xor g_8342_(_4365_, _4474_, _4496_);
  and g_8343_(_4288_, _4496_, _4507_);
  xor g_8344_(_4288_, _4496_, _4518_);
  and g_8345_(_4277_, _4518_, _4529_);
  xor g_8346_(_4277_, _4518_, _4540_);
  and g_8347_(_4190_, _4540_, _4551_);
  xor g_8348_(_4190_, _4540_, _4562_);
  and g_8349_(_3841_, _4562_, _4573_);
  xor g_8350_(_3841_, _4562_, _4584_);
  and g_8351_(_4125_, _4584_, _4595_);
  xor g_8352_(_4125_, _4584_, _4606_);
  and g_8353_(_4147_, _4606_, _4617_);
  xor g_8354_(_4147_, _4606_, _4627_);
  and g_8355_(_4169_, _4627_, _4638_);
  xor g_8356_(_4169_, _4627_, G14[7]);
  or g_8357_(_4551_, _4573_, _4659_);
  or g_8358_(_4507_, _4529_, _4670_);
  and g_8359_(G11[0], G12[8], _4681_);
  and g_8360_(G11[2], G12[6], _4692_);
  and g_8361_(G11[2], G12[7], _4703_);
  and g_8362_(_4223_, _4692_, _4714_);
  xor g_8363_(_4223_, _4692_, _4725_);
  and g_8364_(_4681_, _4725_, _4736_);
  xor g_8365_(_4681_, _4725_, _4747_);
  or g_8366_(_4332_, _4354_, _4758_);
  and g_8367_(_4747_, _4758_, _4769_);
  xor g_8368_(_4747_, _4758_, _4780_);
  and g_8369_(_4234_, _4780_, _4791_);
  xor g_8370_(_4234_, _4780_, _4802_);
  or g_8371_(_4463_, _4485_, _4812_);
  and g_8372_(G11[3], G12[5], _4823_);
  and g_8373_(G12[2], G11[6], _4834_);
  and g_8374_(G12[4], G11[6], _4845_);
  and g_8375_(_3896_, _4834_, _4856_);
  xor g_8376_(_3896_, _4834_, _4867_);
  and g_8377_(_4823_, _4867_, _4878_);
  xor g_8378_(_4823_, _4867_, _4889_);
  or g_8379_(_4420_, _4441_, _4900_);
  and g_8380_(G12[1], G11[7], _4911_);
  and g_8381_(G12[0], G11[8], _4922_);
  and g_8382_(G12[3], G11[8], _4933_);
  and g_8383_(_3623_, _4922_, _4944_);
  xor g_8384_(_3623_, _4922_, _4955_);
  and g_8385_(_4911_, _4955_, _4966_);
  xor g_8386_(_4911_, _4955_, _4977_);
  and g_8387_(_4900_, _4977_, _4988_);
  xor g_8388_(_4900_, _4977_, _4999_);
  and g_8389_(_4889_, _4999_, _5009_);
  xor g_8390_(_4889_, _4999_, _5020_);
  and g_8391_(_4812_, _5020_, _5031_);
  xor g_8392_(_4812_, _5020_, _5042_);
  and g_8393_(_4802_, _5042_, _5053_);
  xor g_8394_(_4802_, _5042_, _5064_);
  and g_8395_(_4670_, _5064_, _5075_);
  xor g_8396_(_4670_, _5064_, _5086_);
  and g_8397_(_4266_, _5086_, _5097_);
  xor g_8398_(_4266_, _5086_, _5108_);
  and g_8399_(_4659_, _5108_, _5119_);
  xor g_8400_(_4659_, _5108_, _5130_);
  and g_8401_(_4595_, _5130_, _5131_);
  not g_8402_(_5131_, _5132_);
  and g_8403_(_4617_, _5130_, _5133_);
  xor g_8404_(_4617_, _5130_, _5134_);
  or g_8405_(_4595_, _5134_, _5135_);
  and g_8406_(_5132_, _5135_, _5136_);
  and g_8407_(_4638_, _5136_, _5137_);
  xor g_8408_(_4638_, _5136_, G14[8]);
  or g_8409_(_5075_, _5097_, _5138_);
  or g_8410_(_5031_, _5053_, _5139_);
  or g_8411_(_4988_, _5009_, _5140_);
  or g_8412_(_4944_, _4966_, _5141_);
  and g_8413_(G12[0], G11[9], _5142_);
  and g_8414_(G12[3], G11[9], _5143_);
  and g_8415_(_3983_, _5142_, _5144_);
  xor g_8416_(_3983_, _5142_, _5145_);
  and g_8417_(G12[1], G11[8], _5146_);
  and g_8418_(_5145_, _5146_, _5147_);
  xor g_8419_(_5145_, _5146_, _5148_);
  and g_8420_(_5141_, _5148_, _5149_);
  xor g_8421_(_5141_, _5148_, _5150_);
  and g_8422_(G11[4], G12[5], _5151_);
  and g_8423_(G12[2], G11[7], _5152_);
  and g_8424_(G12[4], G11[7], _5153_);
  and g_8425_(_4321_, _5152_, _5154_);
  xor g_8426_(_4321_, _5152_, _5155_);
  and g_8427_(_5151_, _5155_, _5156_);
  xor g_8428_(_5151_, _5155_, _5157_);
  and g_8429_(_5150_, _5157_, _5158_);
  xor g_8430_(_5150_, _5157_, _5159_);
  and g_8431_(_5140_, _5159_, _5160_);
  xor g_8432_(_5140_, _5159_, _5161_);
  or g_8433_(_4714_, _4736_, _5162_);
  and g_8434_(G11[3], G12[6], _5163_);
  and g_8435_(G11[3], G12[7], _5164_);
  and g_8436_(_4703_, _5163_, _5165_);
  xor g_8437_(_4703_, _5163_, _5166_);
  and g_8438_(G11[1], G12[8], _5167_);
  and g_8439_(_5166_, _5167_, _5168_);
  xor g_8440_(_5166_, _5167_, _5169_);
  or g_8441_(_4856_, _4878_, _5170_);
  and g_8442_(_5169_, _5170_, _5171_);
  xor g_8443_(_5169_, _5170_, _5172_);
  and g_8444_(_5162_, _5172_, _5173_);
  xor g_8445_(_5162_, _5172_, _5174_);
  and g_8446_(_5161_, _5174_, _5175_);
  xor g_8447_(_5161_, _5174_, _5176_);
  and g_8448_(_5139_, _5176_, _5177_);
  xor g_8449_(_5139_, _5176_, _5178_);
  and g_8450_(G11[0], G12[9], _5179_);
  or g_8451_(_4769_, _4791_, _5180_);
  and g_8452_(_5179_, _5180_, _5181_);
  xor g_8453_(_5179_, _5180_, _5182_);
  and g_8454_(_5178_, _5182_, _5183_);
  xor g_8455_(_5178_, _5182_, _5184_);
  and g_8456_(_5138_, _5184_, _5185_);
  xor g_8457_(_5138_, _5184_, _5186_);
  and g_8458_(_5119_, _5186_, _5187_);
  xor g_8459_(_5119_, _5186_, _5188_);
  and g_8460_(_5131_, _5188_, _5189_);
  xor g_8461_(_5131_, _5188_, _5190_);
  and g_8462_(_5133_, _5190_, _5191_);
  xor g_8463_(_5133_, _5190_, _5192_);
  and g_8464_(_5137_, _5192_, _5193_);
  or g_8465_(_5191_, _5193_, _5194_);
  or g_8466_(_5177_, _5183_, _5195_);
  and g_8467_(G11[0], G12[10], _5196_);
  and g_8468_(G11[1], G12[9], _5197_);
  and g_8469_(G11[1], G12[10], _5198_);
  and g_8470_(_5179_, _5198_, _5199_);
  xor g_8471_(_5196_, _5197_, _5200_);
  or g_8472_(_5171_, _5173_, _5201_);
  and g_8473_(_5200_, _5201_, _5202_);
  xor g_8474_(_5200_, _5201_, _5203_);
  or g_8475_(_5160_, _5175_, _5204_);
  or g_8476_(_5165_, _5168_, _5205_);
  and g_8477_(G11[2], G12[8], _5206_);
  and g_8478_(G11[4], G12[6], _5207_);
  and g_8479_(G11[4], G12[7], _5208_);
  and g_8480_(_5164_, _5207_, _5209_);
  xor g_8481_(_5164_, _5207_, _5210_);
  and g_8482_(_5206_, _5210_, _5211_);
  xor g_8483_(_5206_, _5210_, _5212_);
  or g_8484_(_5154_, _5156_, _5213_);
  and g_8485_(_5212_, _5213_, _5214_);
  xor g_8486_(_5212_, _5213_, _5215_);
  and g_8487_(_5205_, _5215_, _5216_);
  xor g_8488_(_5205_, _5215_, _5217_);
  or g_8489_(_5149_, _5158_, _5218_);
  and g_8490_(G11[5], G12[5], _5219_);
  and g_8491_(G12[2], G11[8], _5220_);
  and g_8492_(G12[4], G11[8], _5221_);
  and g_8493_(_4845_, _5220_, _5222_);
  xor g_8494_(_4845_, _5220_, _5223_);
  and g_8495_(_5219_, _5223_, _5224_);
  xor g_8496_(_5219_, _5223_, _5225_);
  or g_8497_(_5144_, _5147_, _5226_);
  and g_8498_(G12[1], G11[9], _5227_);
  and g_8499_(G12[0], G11[10], _5228_);
  and g_8500_(G12[3], G11[10], _5229_);
  and g_8501_(_4409_, _5228_, _5230_);
  xor g_8502_(_4409_, _5228_, _5231_);
  and g_8503_(_5227_, _5231_, _5232_);
  xor g_8504_(_5227_, _5231_, _5233_);
  and g_8505_(_5226_, _5233_, _5234_);
  xor g_8506_(_5226_, _5233_, _5235_);
  and g_8507_(_5225_, _5235_, _5236_);
  xor g_8508_(_5225_, _5235_, _5237_);
  and g_8509_(_5218_, _5237_, _5238_);
  xor g_8510_(_5218_, _5237_, _5239_);
  and g_8511_(_5217_, _5239_, _5240_);
  xor g_8512_(_5217_, _5239_, _5241_);
  and g_8513_(_5204_, _5241_, _5242_);
  xor g_8514_(_5204_, _5241_, _5243_);
  and g_8515_(_5203_, _5243_, _5244_);
  xor g_8516_(_5203_, _5243_, _5245_);
  and g_8517_(_5195_, _5245_, _5246_);
  xor g_8518_(_5195_, _5245_, _5247_);
  and g_8519_(_5181_, _5247_, _5248_);
  xor g_8520_(_5181_, _5247_, _5249_);
  and g_8521_(_5185_, _5249_, _5250_);
  xor g_8522_(_5185_, _5249_, _5251_);
  or g_8523_(_5187_, _5189_, _5252_);
  xor g_8524_(_5251_, _5252_, _5253_);
  and g_8525_(_5194_, _5253_, _5254_);
  xor g_8526_(_5194_, _5253_, G14[10]);
  and g_8527_(_5189_, _5251_, _5255_);
  or g_8528_(_5246_, _5248_, _5256_);
  or g_8529_(_5242_, _5244_, _5257_);
  and g_8530_(G11[0], G12[11], _5258_);
  and g_8531_(G11[2], G12[9], _5259_);
  and g_8532_(G11[2], G12[10], _5260_);
  and g_8533_(_5198_, _5259_, _5261_);
  xor g_8534_(_5198_, _5259_, _5262_);
  and g_8535_(_5258_, _5262_, _5263_);
  xor g_8536_(_5258_, _5262_, _5264_);
  and g_8537_(_5199_, _5264_, _5265_);
  xor g_8538_(_5199_, _5264_, _5266_);
  or g_8539_(_5214_, _5216_, _5267_);
  and g_8540_(_5266_, _5267_, _5268_);
  xor g_8541_(_5266_, _5267_, _5269_);
  or g_8542_(_5238_, _5240_, _5270_);
  or g_8543_(_5209_, _5211_, _5271_);
  and g_8544_(G11[3], G12[8], _5272_);
  and g_8545_(G11[5], G12[6], _5273_);
  and g_8546_(G11[5], G12[7], _5274_);
  and g_8547_(_5208_, _5273_, _5275_);
  xor g_8548_(_5208_, _5273_, _5276_);
  and g_8549_(_5272_, _5276_, _5277_);
  xor g_8550_(_5272_, _5276_, _5278_);
  or g_8551_(_5222_, _5224_, _5279_);
  and g_8552_(_5278_, _5279_, _5280_);
  xor g_8553_(_5278_, _5279_, _5281_);
  and g_8554_(_5271_, _5281_, _5282_);
  xor g_8555_(_5271_, _5281_, _5283_);
  or g_8556_(_5234_, _5236_, _5284_);
  and g_8557_(G12[5], G11[6], _5285_);
  and g_8558_(G12[2], G11[9], _5286_);
  and g_8559_(G12[4], G11[9], _5287_);
  and g_8560_(_5153_, _5286_, _5288_);
  xor g_8561_(_5153_, _5286_, _5289_);
  and g_8562_(_5285_, _5289_, _5290_);
  xor g_8563_(_5285_, _5289_, _5291_);
  or g_8564_(_5230_, _5232_, _5292_);
  and g_8565_(G12[1], G11[10], _5293_);
  and g_8566_(G12[0], G11[11], _5294_);
  and g_8567_(G12[3], G11[11], _5295_);
  and g_8568_(_4933_, _5294_, _5296_);
  xor g_8569_(_4933_, _5294_, _5297_);
  and g_8570_(_5293_, _5297_, _5298_);
  xor g_8571_(_5293_, _5297_, _5299_);
  and g_8572_(_5292_, _5299_, _5300_);
  xor g_8573_(_5292_, _5299_, _5301_);
  and g_8574_(_5291_, _5301_, _5302_);
  xor g_8575_(_5291_, _5301_, _5303_);
  and g_8576_(_5284_, _5303_, _5304_);
  xor g_8577_(_5284_, _5303_, _5305_);
  and g_8578_(_5283_, _5305_, _5306_);
  xor g_8579_(_5283_, _5305_, _5307_);
  and g_8580_(_5270_, _5307_, _5308_);
  xor g_8581_(_5270_, _5307_, _5309_);
  and g_8582_(_5269_, _5309_, _5310_);
  xor g_8583_(_5269_, _5309_, _5311_);
  and g_8584_(_5257_, _5311_, _5312_);
  xor g_8585_(_5257_, _5311_, _5313_);
  and g_8586_(_5202_, _5313_, _5314_);
  xor g_8587_(_5202_, _5313_, _5315_);
  and g_8588_(_5256_, _5315_, _5316_);
  xor g_8589_(_5256_, _5315_, _5317_);
  and g_8590_(_5187_, _5251_, _5318_);
  or g_8591_(_5250_, _5318_, _5319_);
  xor g_8592_(_5317_, _5319_, _5320_);
  and g_8593_(_5255_, _5320_, _5321_);
  xor g_8594_(_5255_, _5320_, _5322_);
  and g_8595_(_5254_, _5322_, _5323_);
  xor g_8596_(_5254_, _5322_, G14[11]);
  or g_8597_(_5321_, _5323_, _5324_);
  and g_8598_(_5317_, _5318_, _5325_);
  and g_8599_(_5250_, _5317_, _5326_);
  or g_8600_(_5312_, _5314_, _5327_);
  or g_8601_(_5308_, _5310_, _5328_);
  and g_8602_(G11[0], G12[12], _5329_);
  or g_8603_(_5261_, _5263_, _5330_);
  and g_8604_(G11[1], G12[11], _5331_);
  and g_8605_(G11[3], G12[9], _5332_);
  and g_8606_(G11[3], G12[10], _5333_);
  and g_8607_(_5260_, _5332_, _5334_);
  xor g_8608_(_5260_, _5332_, _5335_);
  and g_8609_(_5331_, _5335_, _5336_);
  xor g_8610_(_5331_, _5335_, _5337_);
  and g_8611_(_5330_, _5337_, _5338_);
  xor g_8612_(_5330_, _5337_, _5339_);
  and g_8613_(_5329_, _5339_, _5340_);
  xor g_8614_(_5329_, _5339_, _5341_);
  or g_8615_(_5280_, _5282_, _5342_);
  and g_8616_(_5341_, _5342_, _5343_);
  xor g_8617_(_5341_, _5342_, _5344_);
  and g_8618_(_5265_, _5344_, _5345_);
  xor g_8619_(_5265_, _5344_, _5346_);
  or g_8620_(_5304_, _5306_, _5347_);
  or g_8621_(_5275_, _5277_, _5348_);
  and g_8622_(G11[4], G12[8], _5349_);
  and g_8623_(G11[6], G12[6], _5350_);
  and g_8624_(G11[6], G12[7], _5351_);
  and g_8625_(_5274_, _5350_, _5352_);
  xor g_8626_(_5274_, _5350_, _5353_);
  and g_8627_(_5349_, _5353_, _5354_);
  xor g_8628_(_5349_, _5353_, _5355_);
  or g_8629_(_5288_, _5290_, _5356_);
  and g_8630_(_5355_, _5356_, _5357_);
  xor g_8631_(_5355_, _5356_, _5358_);
  and g_8632_(_5348_, _5358_, _5359_);
  xor g_8633_(_5348_, _5358_, _5360_);
  or g_8634_(_5300_, _5302_, _5361_);
  and g_8635_(G12[5], G11[7], _5362_);
  and g_8636_(G12[2], G11[10], _5363_);
  and g_8637_(G12[4], G11[10], _5364_);
  and g_8638_(_5221_, _5363_, _5365_);
  xor g_8639_(_5221_, _5363_, _5366_);
  and g_8640_(_5362_, _5366_, _5367_);
  xor g_8641_(_5362_, _5366_, _5368_);
  or g_8642_(_5296_, _5298_, _5369_);
  and g_8643_(G12[1], G11[11], _5370_);
  and g_8644_(G12[0], G11[12], _5371_);
  and g_8645_(G12[3], G11[12], _5372_);
  and g_8646_(_5143_, _5371_, _5373_);
  xor g_8647_(_5143_, _5371_, _5374_);
  and g_8648_(_5370_, _5374_, _5375_);
  xor g_8649_(_5370_, _5374_, _5376_);
  and g_8650_(_5369_, _5376_, _5377_);
  xor g_8651_(_5369_, _5376_, _5378_);
  and g_8652_(_5368_, _5378_, _5379_);
  xor g_8653_(_5368_, _5378_, _5380_);
  and g_8654_(_5361_, _5380_, _5381_);
  xor g_8655_(_5361_, _5380_, _5382_);
  and g_8656_(_5360_, _5382_, _5383_);
  xor g_8657_(_5360_, _5382_, _5384_);
  and g_8658_(_5347_, _5384_, _5385_);
  xor g_8659_(_5347_, _5384_, _5386_);
  and g_8660_(_5346_, _5386_, _5387_);
  xor g_8661_(_5346_, _5386_, _5388_);
  and g_8662_(_5328_, _5388_, _5389_);
  xor g_8663_(_5328_, _5388_, _5390_);
  and g_8664_(_5268_, _5390_, _5391_);
  xor g_8665_(_5268_, _5390_, _5392_);
  and g_8666_(_5327_, _5392_, _5393_);
  xor g_8667_(_5327_, _5392_, _5394_);
  and g_8668_(_5316_, _5394_, _5395_);
  xor g_8669_(_5316_, _5394_, _5396_);
  and g_8670_(_5326_, _5396_, _5397_);
  xor g_8671_(_5326_, _5396_, _5398_);
  and g_8672_(_5325_, _5398_, _5399_);
  xor g_8673_(_5325_, _5398_, _5400_);
  and g_8674_(_5324_, _5400_, _5401_);
  xor g_8675_(_5324_, _5400_, G14[12]);
  or g_8676_(_5399_, _5401_, _5402_);
  or g_8677_(_5389_, _5391_, _5403_);
  or g_8678_(_5343_, _5345_, _5404_);
  or g_8679_(_5385_, _5387_, _5405_);
  or g_8680_(_5338_, _5340_, _5406_);
  and g_8681_(G11[0], G12[13], _5407_);
  and g_8682_(G11[1], G12[12], _5408_);
  and g_8683_(G11[1], G12[13], _5409_);
  and g_8684_(_5329_, _5409_, _5410_);
  xor g_8685_(_5407_, _5408_, _5411_);
  or g_8686_(_5334_, _5336_, _5412_);
  and g_8687_(G11[2], G12[11], _5413_);
  and g_8688_(G11[4], G12[9], _5414_);
  and g_8689_(G11[4], G12[10], _5415_);
  and g_8690_(_5333_, _5414_, _5416_);
  xor g_8691_(_5333_, _5414_, _5417_);
  and g_8692_(_5413_, _5417_, _5418_);
  xor g_8693_(_5413_, _5417_, _5419_);
  and g_8694_(_5412_, _5419_, _5420_);
  xor g_8695_(_5412_, _5419_, _5421_);
  and g_8696_(_5411_, _5421_, _5422_);
  xor g_8697_(_5411_, _5421_, _5423_);
  or g_8698_(_5357_, _5359_, _5424_);
  and g_8699_(_5423_, _5424_, _5425_);
  xor g_8700_(_5423_, _5424_, _5426_);
  and g_8701_(_5406_, _5426_, _5427_);
  xor g_8702_(_5406_, _5426_, _5428_);
  or g_8703_(_5381_, _5383_, _5429_);
  or g_8704_(_5352_, _5354_, _5430_);
  and g_8705_(G11[5], G12[8], _5431_);
  and g_8706_(G12[6], G11[7], _5432_);
  and g_8707_(G11[7], G12[7], _5433_);
  and g_8708_(_5351_, _5432_, _5434_);
  xor g_8709_(_5351_, _5432_, _5435_);
  and g_8710_(_5431_, _5435_, _5436_);
  xor g_8711_(_5431_, _5435_, _5437_);
  or g_8712_(_5365_, _5367_, _5438_);
  and g_8713_(_5437_, _5438_, _5439_);
  xor g_8714_(_5437_, _5438_, _5440_);
  and g_8715_(_5430_, _5440_, _5441_);
  xor g_8716_(_5430_, _5440_, _5442_);
  or g_8717_(_5377_, _5379_, _5443_);
  and g_8718_(G12[5], G11[8], _5444_);
  and g_8719_(G12[2], G11[11], _5445_);
  and g_8720_(G12[4], G11[11], _5446_);
  and g_8721_(_5287_, _5445_, _5447_);
  xor g_8722_(_5287_, _5445_, _5448_);
  and g_8723_(_5444_, _5448_, _5449_);
  xor g_8724_(_5444_, _5448_, _5450_);
  or g_8725_(_5373_, _5375_, _5451_);
  and g_8726_(G12[1], G11[12], _5452_);
  and g_8727_(G12[0], G11[13], _5453_);
  and g_8728_(G12[3], G11[13], _5454_);
  and g_8729_(_5229_, _5453_, _5455_);
  xor g_8730_(_5229_, _5453_, _5456_);
  and g_8731_(_5452_, _5456_, _5457_);
  xor g_8732_(_5452_, _5456_, _5458_);
  and g_8733_(_5451_, _5458_, _5459_);
  xor g_8734_(_5451_, _5458_, _5460_);
  and g_8735_(_5450_, _5460_, _5461_);
  xor g_8736_(_5450_, _5460_, _5462_);
  and g_8737_(_5443_, _5462_, _5463_);
  xor g_8738_(_5443_, _5462_, _5464_);
  and g_8739_(_5442_, _5464_, _5465_);
  xor g_8740_(_5442_, _5464_, _5466_);
  and g_8741_(_5429_, _5466_, _5467_);
  xor g_8742_(_5429_, _5466_, _5468_);
  and g_8743_(_5428_, _5468_, _5469_);
  xor g_8744_(_5428_, _5468_, _5470_);
  and g_8745_(_5405_, _5470_, _5471_);
  xor g_8746_(_5405_, _5470_, _5472_);
  and g_8747_(_5404_, _5472_, _5473_);
  xor g_8748_(_5404_, _5472_, _5474_);
  and g_8749_(_5403_, _5474_, _5475_);
  xor g_8750_(_5403_, _5474_, _5476_);
  and g_8751_(_5393_, _5476_, _5477_);
  xor g_8752_(_5393_, _5476_, _5478_);
  or g_8753_(_5395_, _5397_, _5479_);
  xor g_8754_(_5478_, _5479_, _5480_);
  and g_8755_(_5402_, _5480_, _5481_);
  xor g_8756_(_5402_, _5480_, G14[13]);
  and g_8757_(_5397_, _5478_, _5482_);
  or g_8758_(_5481_, _5482_, _5483_);
  or g_8759_(_5471_, _5473_, _5484_);
  or g_8760_(_5425_, _5427_, _5485_);
  and g_8761_(_5410_, _5485_, _5486_);
  xor g_8762_(_5410_, _5485_, _5487_);
  or g_8763_(_5467_, _5469_, _5488_);
  or g_8764_(_5420_, _5422_, _5489_);
  and g_8765_(G11[0], G12[14], _5490_);
  and g_8766_(G11[2], G12[12], _5491_);
  and g_8767_(G11[2], G12[13], _5492_);
  and g_8768_(_5409_, _5491_, _5493_);
  xor g_8769_(_5409_, _5491_, _5494_);
  and g_8770_(_5490_, _5494_, _5495_);
  xor g_8771_(_5490_, _5494_, _5496_);
  or g_8772_(_5416_, _5418_, _5497_);
  and g_8773_(G11[3], G12[11], _5498_);
  and g_8774_(G11[5], G12[9], _5499_);
  and g_8775_(G11[5], G12[10], _5500_);
  and g_8776_(_5415_, _5499_, _5501_);
  xor g_8777_(_5415_, _5499_, _5502_);
  and g_8778_(_5498_, _5502_, _5503_);
  xor g_8779_(_5498_, _5502_, _5504_);
  and g_8780_(_5497_, _5504_, _5505_);
  xor g_8781_(_5497_, _5504_, _5506_);
  and g_8782_(_5496_, _5506_, _5507_);
  xor g_8783_(_5496_, _5506_, _5508_);
  or g_8784_(_5439_, _5441_, _5509_);
  and g_8785_(_5508_, _5509_, _5510_);
  xor g_8786_(_5508_, _5509_, _5511_);
  and g_8787_(_5489_, _5511_, _5512_);
  xor g_8788_(_5489_, _5511_, _5513_);
  or g_8789_(_5463_, _5465_, _5514_);
  or g_8790_(_5434_, _5436_, _5515_);
  and g_8791_(G11[6], G12[8], _5516_);
  and g_8792_(G12[6], G11[8], _5517_);
  and g_8793_(G12[7], G11[8], _5518_);

endmodule
