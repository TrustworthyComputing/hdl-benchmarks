module c880(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G7, G8, G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878, G879, G880, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, G293, G295, G296, G343, G349, G350, G369, G812, G829, G830, G831, G832, G844, G849, G850, G851;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G7, G8, G9;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878, G879, G880;
  lut lut_gate1(0x7, G8, 455, G855);
  lut lut_gate2(0x8, G6, G16, 455);
  lut lut_gate3(0x7, G17, 456, G856);
  lut lut_gate4(0x8, G7, G6, 456);
  lut lut_gate5(0x7, G8, 456, G857);
  lut lut_gate6(0x7, G18, G19, G858);
  lut lut_gate7(0x7, 458, 457, G859);
  lut lut_gate8(0x8, G1, G2, 457);
  lut lut_gate9(0x8, G3, G4, 458);
  lut lut_gate10(0x8, 459, G857, G860);
  lut lut_gate11(0x8, 460, 458, 459);
  lut lut_gate12(0x8, G5, G1, 460);
  lut lut_gate13(0xb, G23, 296, G864);
  lut lut_gate14(0x1, G20, G21, 296);
  lut lut_gate15(0x4, 459, G857, G865);
  lut lut_gate16(0x7, G9, 460, G866);
  lut lut_gate17(0xb, G22, 296, G869);
  lut lut_gate18(0x4, 298, 307, 297);
  lut lut_gate19(0x1, 304, 299, 298);
  lut lut_gate20(0x4, G39, 300, 299);
  lut lut_gate21(0x4, G1, 301, 300);
  lut lut_gate22(0x8, G4, 302, 301);
  lut lut_gate23(0x1, 303, G866, 302);
  lut lut_gate24(0x8, G11, G40, 303);
  lut lut_gate25(0x4, G31, 418, 304);
  lut lut_gate26(0x8, G8, 306, 305);
  lut lut_gate27(0x8, G11, G16, 306);
  lut lut_gate28(0x8, 310, 308, 307);
  lut lut_gate29(0x4, 309, G866, 308);
  lut lut_gate30(0x8, G17, 455, 309);
  lut lut_gate31(0x4, G10, G60, 310);
  lut lut_gate32(0x8, G50, G30, 311);
  lut lut_gate33(0x8, 316, 313, 312);
  lut lut_gate34(0x8, G14, 314, 313);
  lut lut_gate35(0x8, 315, 457, 314);
  lut lut_gate36(0x8, G10, G3, 315);
  lut lut_gate37(0x8, 318, 317, 316);
  lut lut_gate38(0x8, G12, G11, 317);
  lut lut_gate39(0x8, G13, G8, 318);
  lut lut_gate40(0x8, G55, G59, 319);
  lut lut_gate41(0x8, G52, 321, 320);
  lut lut_gate42(0x9, G48, 297, 321);
  lut lut_gate43(0x8, G51, 323, 322);
  lut lut_gate44(0x6, G58, 321, 323);
  lut lut_gate45(0x8, G51, 325, 324);
  lut lut_gate46(0x9, 334, 419, 325);
  lut lut_gate47(0x4, 328, 327, 326);
  lut lut_gate48(0x4, G37, 300, 327);
  lut lut_gate49(0x1, 307, 329, 328);
  lut lut_gate50(0x4, G30, 418, 329);
  lut lut_gate51(0x4, 332, 331, 330);
  lut lut_gate52(0x4, G36, 300, 331);
  lut lut_gate53(0x1, 307, 333, 332);
  lut lut_gate54(0x4, G29, 418, 333);
  lut lut_gate55(0x9, G45, 335, 334);
  lut lut_gate56(0x4, 337, 336, 335);
  lut lut_gate57(0x4, G35, 300, 336);
  lut lut_gate58(0x1, 307, 338, 337);
  lut lut_gate59(0x4, G28, 418, 338);
  lut lut_gate60(0x8, G27, G50, 339);
  lut lut_gate61(0x8, G52, 334, 340);
  lut lut_gate62(0x8, G51, 342, 341);
  lut lut_gate63(0x9, 343, 420, 342);
  lut lut_gate64(0x9, G46, 330, 343);
  lut lut_gate65(0x8, G28, G50, 344);
  lut lut_gate66(0x8, G56, G55, 345);
  lut lut_gate67(0x8, G52, 343, 346);
  lut lut_gate68(0x4, G51, 348, 347);
  lut lut_gate69(0x9, 349, 421, 348);
  lut lut_gate70(0x9, G47, 326, 349);
  lut lut_gate71(0x1, 352, 351, 350);
  lut lut_gate72(0x8, G29, G50, 351);
  lut lut_gate73(0x8, G57, G55, 352);
  lut lut_gate74(0x8, G52, 349, 353);
  lut lut_gate75(0x4, 355, 362, 354);
  lut lut_gate76(0x4, 358, 356, 355);
  lut lut_gate77(0x8, G39, 357, 356);
  lut lut_gate78(0x8, G10, 302, 357);
  lut lut_gate79(0x1, 361, 359, 358);
  lut lut_gate80(0x8, 360, 308, 359);
  lut lut_gate81(0x4, G4, G60, 360);
  lut lut_gate82(0x8, G38, G34, 361);
  lut lut_gate83(0x4, G27, 418, 362);
  lut lut_gate84(0x8, G37, 357, 363);
  lut lut_gate85(0x8, G36, 357, 364);
  lut lut_gate86(0x4, G25, 418, 365);
  lut lut_gate87(0x4, 367, 371, 366);
  lut lut_gate88(0x4, 369, 368, 367);
  lut lut_gate89(0x8, G35, 357, 368);
  lut lut_gate90(0x1, 370, 359, 369);
  lut lut_gate91(0x8, G34, G2, 370);
  lut lut_gate92(0x4, G24, 418, 371);
  lut lut_gate93(0x4, G51, 373, 372);
  lut lut_gate94(0x6, 374, 429, 373);
  lut lut_gate95(0x9, G44, 354, 374);
  lut lut_gate96(0x8, G26, G50, 375);
  lut lut_gate97(0x8, G52, 374, 376);
  lut lut_gate98(0x8, G51, 378, 377);
  lut lut_gate99(0x9, 379, 426, 378);
  lut lut_gate100(0x9, G41, 366, 379);
  lut lut_gate101(0x8, G60, G50, 380);
  lut lut_gate102(0x8, G52, 379, 381);
  lut lut_gate103(0x8, G51, 383, 382);
  lut lut_gate104(0x9, 384, 427, 383);
  lut lut_gate105(0x9, G42, 436, 384);
  lut lut_gate106(0x8, G24, G50, 385);
  lut lut_gate107(0x8, G52, 384, 386);
  lut lut_gate108(0x8, G51, 388, 387);
  lut lut_gate109(0x9, 389, 428, 388);
  lut lut_gate110(0x9, G43, 433, 389);
  lut lut_gate111(0x8, G25, G50, 390);
  lut lut_gate112(0x8, G52, 389, 391);
  lut lut_gate113(0x8, G17, 306, G861);
  lut lut_gate114(0x8, G17, 392, G862);
  lut lut_gate115(0x8, G11, G7, 392);
  lut lut_gate116(0x8, G8, 392, G863);
  lut lut_gate117(0x7, 393, 314, G867);
  lut lut_gate118(0x8, G12, G6, 393);
  lut lut_gate119(0x7, 394, 314, G868);
  lut lut_gate120(0x8, G15, 317, 394);
  lut lut_gate121(0x6, 400, 395, G870);
  lut lut_gate122(0x9, 398, 396, 395);
  lut lut_gate123(0x9, G25, 397, 396);
  lut lut_gate124(0x6, G32, G26, 397);
  lut lut_gate125(0x6, G28, 399, 398);
  lut lut_gate126(0x6, G33, G29, 399);
  lut lut_gate127(0x9, 402, 401, 400);
  lut lut_gate128(0x9, G31, G30, 401);
  lut lut_gate129(0x9, G24, G27, 402);
  lut lut_gate130(0x6, 409, 403, G871);
  lut lut_gate131(0x9, 407, 404, 403);
  lut lut_gate132(0x9, 406, 405, 404);
  lut lut_gate133(0x9, G45, G48, 405);
  lut lut_gate134(0x9, G42, G41, 406);
  lut lut_gate135(0x9, G46, 408, 407);
  lut lut_gate136(0x6, G49, G47, 408);
  lut lut_gate137(0x6, G43, 410, 409);
  lut lut_gate138(0x6, G32, G44, 410);
  lut lut_gate139(0xf8, G54, G48, G53, 411);
  lut lut_gate140(0x01, 320, 319, 311, 412);
  lut lut_gate141(0x4, 412, 322, 413);
  lut lut_gate142(0xb0, 413, 411, 297, 414);
  lut lut_gate143(0x70, 414, G48, 312, G872);
  lut lut_gate144(0x4, 303, G866, 415);
  lut lut_gate145(0x9f, 415, G4, G8, 416);
  lut lut_gate146(0x40, G9, 457, 305, 417);
  lut lut_gate147(0x70, 416, G4, 417, 418);
  lut lut_gate148(0x10, 448, 340, 324, G873);
  lut lut_gate149(0x4, 330, 420, G46, 419);
  lut lut_gate150(0x71, 326, 421, G47, 420);
  lut lut_gate151(0xb2, G58, 297, G48, 421);
  lut lut_gate152(0xf8, G54, G46, G53, 422);
  lut lut_gate153(0x01, 346, 345, 344, 423);
  lut lut_gate154(0x4, 423, 341, 424);
  lut lut_gate155(0x70, 424, G46, 312, 425);
  lut lut_gate156(0xb0, 425, 422, 330, G874);
  lut lut_gate157(0x10, 451, 353, 347, G875);
  lut lut_gate158(0x4, 366, 426, G41, G876);
  lut lut_gate159(0x4, 436, 427, G42, 426);
  lut lut_gate160(0x4, 433, 428, G43, 427);
  lut lut_gate161(0x4, 354, 429, G44, 428);
  lut lut_gate162(0x4, 419, 335, G45, 429);
  lut lut_gate163(0x1, 363, 359, 430);
  lut lut_gate164(0x8f, 416, 417, G4, 431);
  lut lut_gate165(0x70, 430, G26, 431, 432);
  lut lut_gate166(0x70, 432, G4, G34, 433);
  lut lut_gate167(0x7f, 360, 309, 460, 434);
  lut lut_gate168(0x4f, G9, 434, G34, 435);
  lut lut_gate169(0x10, 435, 365, 364, 436);
  lut lut_gate170(0xf8, G54, G44, G53, 437);
  lut lut_gate171(0x01, 376, 375, 372, 438);
  lut lut_gate172(0x70, 438, G44, 312, 439);
  lut lut_gate173(0xb0, 439, 437, 354, G877);
  lut lut_gate174(0x10, 454, 381, 377, G878);
  lut lut_gate175(0xf8, G54, G42, G53, 440);
  lut lut_gate176(0x01, 386, 385, 382, 441);
  lut lut_gate177(0x70, 441, G42, 312, 442);
  lut lut_gate178(0xb0, 442, 440, 436, G879);
  lut lut_gate179(0xf8, G54, G43, G53, 443);
  lut lut_gate180(0x01, 391, 390, 387, 444);
  lut lut_gate181(0x70, 444, G43, 312, 445);
  lut lut_gate182(0xb0, 445, 443, 433, G880);
  lut lut_gate183(0xf8, G54, G45, G53, 446);
  lut lut_gate184(0x07, 339, G45, 312, 447);
  lut lut_gate185(0xb0, 447, 446, 335, 448);
  lut lut_gate186(0xf8, G54, G47, G53, 449);
  lut lut_gate187(0x70, 350, G47, 312, 450);
  lut lut_gate188(0xb0, 450, 449, 326, 451);
  lut lut_gate189(0xf8, G54, G41, G53, 452);
  lut lut_gate190(0x07, 380, G41, 312, 453);
  lut lut_gate191(0xb0, 453, 452, 366, 454);

endmodule
