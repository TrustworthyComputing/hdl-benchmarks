module c3540(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, G1022, G2943, G2974, G2985, G3005, G3030, G3100, G3135, G3195, G3202, G3226, G3257, G3265, G3266, G3267, G3275, G3281, G3294, G3300, G3301, G3311, G3312, G3320, G3332, G3341, G3342, G3343, G3345, G3373, G3376, G3379, G3394, G3515, G3516, G722, G723, G724, G725, G731, G734, G735, G736, G739, G742, G745, G749, G781, G786, G791, G792, G793, G794, G795, G796, G797, G798, G799, G816, G831, G882, G883, G890, G891, G892, G893, G894, G897, G898, G901, G904, G907, G910, G913, G916, G919, G922, G925;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540;
  lut lut_gate1(0x50cf, 0928, 0935, 0943, 0944, 0927);
  lut lut_gate2(0x0c05, G14, 0932, 0929, 0934, 0928);
  lut lut_gate3(0x0, 0931, 0930, G3, 0929);
  lut lut_gate4(0x07ff, G1, G2, G4, G3, 0930);
  lut lut_gate5(0x1513, G1, G3, G4, G2, 0931);
  lut lut_gate6(0xc500, 0933, G4, G39, G12, 0932);
  lut lut_gate7(0x40, G2, G1, G3, 0933);
  lut lut_gate8(0x40, G3, G2, G1, 0934);
  lut lut_gate9(0x0e, 0936, 0939, 0937, 0935);
  lut lut_gate10(0x40, G38, 0938, G5, 0936);
  lut lut_gate11(0x7000, G1, G2, G4, G5, 0937);
  lut lut_gate12(0x1, G6, G1, 0938);
  lut lut_gate13(0x0007, 0940, 0942, 0941, G35, 0939);
  lut lut_gate14(0xfe00, G37, G1, G5, G6, 0940);
  lut lut_gate15(0x1, G49, G4, 0941);
  lut lut_gate16(0xca, G4, G36, G41, 0942);
  lut lut_gate17(0x1, G24, G23, 0943);
  lut lut_gate18(0x1, G26, G25, 0944);
  lut lut_gate19(0x4, 0946, 0928, 0945);
  lut lut_gate20(0x8, 0949, 0947, 0946);
  lut lut_gate21(0x4, 0948, G2, 0947);
  lut lut_gate22(0x1, G3, G1, 0948);
  lut lut_gate23(0x8, G48, G27, 0949);
  lut lut_gate24(0x4, 0687, G3, 0686);
  lut lut_gate25(0x4, G4, G2, 0687);
  lut lut_gate26(0xf4, 0689, 0701, G41, 0688);
  lut lut_gate27(0x80, 0699, 0697, 0690, 0689);
  lut lut_gate28(0x0e00, 0691, 0694, 0696, G7, 0690);
  lut lut_gate29(0xeee0, G13, 0692, G8, 0693, 0691);
  lut lut_gate30(0x4000, G26, G25, G3, G24, 0692);
  lut lut_gate31(0x001f, G26, G3, G25, G24, 0693);
  lut lut_gate32(0x1, G12, 0695, 0694);
  lut lut_gate33(0x01ff, G3, G25, G24, G26, 0695);
  lut lut_gate34(0x1f00, G26, G3, G25, G24, 0696);
  lut lut_gate35(0xeee0, G9, 0692, G11, 0698, 0697);
  lut lut_gate36(0x1000, G26, G3, G25, G24, 0698);
  lut lut_gate37(0x00f4, G4, 0700, G10, G22, 0699);
  lut lut_gate38(0x1000, G3, G25, G26, G24, 0700);
  lut lut_gate39(0x000, 0704, 0702, 0693, G44, 0701);
  lut lut_gate40(0x0, 0703, 0696, G45, 0702);
  lut lut_gate41(0x0e, 0692, G39, G43, 0703);
  lut lut_gate42(0xf100, G4, 0700, G46, G42, 0704);
  lut lut_gate43(0x4, 0706, G6, 0705);
  lut lut_gate44(0x8, G5, 0947, 0706);
  lut lut_gate45(0xe1, 0740, 0751, 0708, 0707);
  lut lut_gate46(0x00ef, 0946, 0737, 0709, 0739, 0708);
  lut lut_gate47(0x8000, 0729, 0721, 0711, 0710, 0709);
  lut lut_gate48(0x10, 0935, 0943, 0928, 0710);
  lut lut_gate49(0xc5, 0712, 0720, 0715, 0711);
  lut lut_gate50(0x0305, G13, 0713, 0931, 0714, 0712);
  lut lut_gate51(0xc500, 0933, G4, G14, G11, 0713);
  lut lut_gate52(0xf800, G3, G2, G4, G1, 0714);
  lut lut_gate53(0x01, 0943, 0716, 0936, 0715);
  lut lut_gate54(0x00ef, 0937, 0718, 0719, 0717, 0716);
  lut lut_gate55(0xfe00, G36, G6, G5, G1, 0717);
  lut lut_gate56(0x35, G4, G35, G40, 0718);
  lut lut_gate57(0x10, G34, G49, G4, 0719);
  lut lut_gate58(0x01, 0944, 0716, 0936, 0720);
  lut lut_gate59(0xc5, 0722, 0728, 0723, 0721);
  lut lut_gate60(0x0503, G12, 0891, 0934, 0931, 0722);
  lut lut_gate61(0x01, 0943, 0724, 0936, 0723);
  lut lut_gate62(0x00fe, 0937, 0726, 0725, 0727, 0724);
  lut lut_gate63(0xfe00, G35, G6, G5, G1, 0725);
  lut lut_gate64(0x10, G33, G49, G4, 0726);
  lut lut_gate65(0xca, G4, G34, G39, 0727);
  lut lut_gate66(0x01, 0944, 0724, 0936, 0728);
  lut lut_gate67(0x05fc, 0733, 0730, 0943, 0944, 0729);
  lut lut_gate68(0x008f, 0937, 0731, G32, 0941, 0730);
  lut lut_gate69(0x3500, 0732, 0938, G38, G34, 0731);
  lut lut_gate70(0x53, G4, G14, G33, 0732);
  lut lut_gate71(0x0503, G11, 0734, 0934, 0931, 0733);
  lut lut_gate72(0x0, 0930, 0735, 0736, 0734);
  lut lut_gate73(0xfe00, G3, G11, G12, G13, 0735);
  lut lut_gate74(0xfcfa, G4, G3, G12, G9, 0736);
  lut lut_gate75(0x5c, 0729, 0733, 0738, 0737);
  lut lut_gate76(0x4, 0723, 0722, 0738);
  lut lut_gate77(0x4000, 0715, 0721, 0729, 0712, 0739);
  lut lut_gate78(0x50cf, 0741, 0745, 0943, 0944, 0740);
  lut lut_gate79(0x000e, 0743, 0742, 0930, 0744, 0741);
  lut lut_gate80(0xbc00, G10, G3, 0930, G1, 0742);
  lut lut_gate81(0x4, 0934, G10, 0743);
  lut lut_gate82(0xfcfa, G4, G3, G11, G8, 0744);
  lut lut_gate83(0x0e, 0746, 0748, 0937, 0745);
  lut lut_gate84(0x8, G38, 0747, 0746);
  lut lut_gate85(0x0e, G1, G5, G6, 0747);
  lut lut_gate86(0x0007, 0749, 0750, 0941, G31, 0748);
  lut lut_gate87(0xf100, G33, G1, G6, G5, 0749);
  lut lut_gate88(0xca, G4, G32, G13, 0750);
  lut lut_gate89(0x4, 0946, 0741, 0751);
  lut lut_gate90(0xa300, G47, 0946, 0893, 0753, 0752);
  lut lut_gate91(0x8000, 0729, 0721, 0711, 0927, 0753);
  lut lut_gate92(0x9, 0751, 0740, 0754);
  lut lut_gate93(0x0, 0756, 0867, 0693, G40, 0755);
  lut lut_gate94(0xe0ee, G41, 0696, G13, 0698, 0756);
  lut lut_gate95(0xb0bb, G21, 0692, G19, 0696, 0757);
  lut lut_gate96(0xffe0, 0771, 0767, 0777, 0758, G3531);
  lut lut_gate97(0x008f, 0706, 0708, 0765, 0759, 0758);
  lut lut_gate98(0x6, 0761, G3526, 0759);
  lut lut_gate99(0x6000, G47, 0760, 0945, 0927, G3526);
  lut lut_gate100(0x553c, 0712, 0715, 0946, 0720, 0760);
  lut lut_gate101(0x0, 0764, 0762, 0763, 0760, 0761);
  lut lut_gate102(0x10, 0715, 0712, 0946, 0762);
  lut lut_gate103(0x0100, 0935, 0943, 0946, 0928, 0763);
  lut lut_gate104(0x553c, 0722, 0723, 0946, 0728, 0764);
  lut lut_gate105(0x827, 0766, 0945, 0927, G47, 0765);
  lut lut_gate106(0x9, 0763, 0760, 0766);
  lut lut_gate107(0x5ca3, 0768, 0769, 0770, G3526, 0767);
  lut lut_gate108(0xb4, 0729, 0946, 0733, 0768);
  lut lut_gate109(0xf400, 0764, 0762, 0760, 0763, 0769);
  lut lut_gate110(0x4, 0738, 0946, 0770);
  lut lut_gate111(0x70, 0898, 0768, 0686, 0771);
  lut lut_gate112(0xb0bb, G21, 0693, G20, 0696, 0772);
  lut lut_gate113(0x00f4, G4, 0700, G7, G19, 0773);
  lut lut_gate114(0xf100, G4, 0700, G43, G39, 0774);
  lut lut_gate115(0xe0ee, G41, 0693, G13, 0695, 0775);
  lut lut_gate116(0xe0ee, G42, 0696, 0698, G14, 0776);
  lut lut_gate117(0xff10, G1, G6, G3, G2, 0777);
  lut lut_gate118(0x7557, 0708, 0765, 0706, 0778, G3532);
  lut lut_gate119(0x07, 0902, 0765, 0777, 0778);
  lut lut_gate120(0x0e00, 0780, G4, 0692, G12, 0779);
  lut lut_gate121(0xeee0, G8, 0692, 0698, G10, 0780);
  lut lut_gate122(0xe0ee, G22, 0696, 0700, 0782, 0781);
  lut lut_gate123(0x4, G9, G21, 0782);
  lut lut_gate124(0x40, 0787, 0784, G40, 0783);
  lut lut_gate125(0x0, 0785, 0786, 0695, G39, 0784);
  lut lut_gate126(0xb0bb, G43, 0693, G44, 0696, 0785);
  lut lut_gate127(0x0b, 0692, G14, G42, 0786);
  lut lut_gate128(0xf100, G4, 0700, G45, G41, 0787);
  lut lut_gate129(0x0, 0790, 0789, 0693, G42, 0788);
  lut lut_gate130(0x0, 0692, G41, G13, 0789);
  lut lut_gate131(0xe0ee, G43, 0696, 0695, G14, 0790);
  lut lut_gate132(0x0b, 0700, G8, G20, 0791);
  lut lut_gate133(0xe0ee, G22, 0693, 0698, G9, 0792);
  lut lut_gate134(0xb, 0793, 0837, G3534);
  lut lut_gate135(0xfc45, 0833, 0794, 0706, 0777, 0793);
  lut lut_gate136(0x0bb0, 0830, 0828, 0826, 0795, 0794);
  lut lut_gate137(0xe0, 0910, 0708, 0825, 0795);
  lut lut_gate138(0x50cf, 0797, 0802, 0943, 0944, 0796);
  lut lut_gate139(0x000e, 0800, 0798, 0930, 0801, 0797);
  lut lut_gate140(0xac, G8, 0934, 0799, 0798);
  lut lut_gate141(0x0733, G1, G2, G3, G4, 0799);
  lut lut_gate142(0x1400, G3, G8, G9, 0930, 0800);
  lut lut_gate143(0xfcf5, G4, G3, G9, G22, 0801);
  lut lut_gate144(0x0e, 0746, 0803, 0937, 0802);
  lut lut_gate145(0x0700, 0805, 0804, 0941, G29, 0803);
  lut lut_gate146(0xf100, G31, G1, G6, G5, 0804);
  lut lut_gate147(0x35, G4, G30, G11, 0805);
  lut lut_gate148(0x50cf, 0807, 0811, 0943, 0944, 0806);
  lut lut_gate149(0x0503, G7, 0808, 0934, 0799, 0807);
  lut lut_gate150(0x0, 0930, 0809, 0810, 0808);
  lut lut_gate151(0xfe00, G3, G9, G7, G8, 0809);
  lut lut_gate152(0xfcf5, G4, G3, G8, G21, 0810);
  lut lut_gate153(0x00f4, 0746, 0937, 0812, 0813, 0811);
  lut lut_gate154(0x0bbb, G28, 0941, G30, 0747, 0812);
  lut lut_gate155(0xca, G4, G29, G10, 0813);
  lut lut_gate156(0x50cf, 0815, 0818, 0943, 0944, 0814);
  lut lut_gate157(0x0e, 0816, 0930, 0817, 0815);
  lut lut_gate158(0xac, G9, 0714, 0799, 0816);
  lut lut_gate159(0xf3f5, G4, G3, G10, G7, 0817);
  lut lut_gate160(0x0e, 0746, 0819, 0937, 0818);
  lut lut_gate161(0x0700, 0821, 0820, 0941, G30, 0819);
  lut lut_gate162(0xf100, G32, G1, G6, G5, 0820);
  lut lut_gate163(0x35, G4, G31, G12, 0821);
  lut lut_gate164(0x10, 0818, 0943, 0815, 0822);
  lut lut_gate165(0x10, 0802, 0943, 0797, 0823);
  lut lut_gate166(0x10, 0745, 0943, 0741, 0824);
  lut lut_gate167(0x8000, 0814, 0806, 0796, 0740, 0825);
  lut lut_gate168(0x8, G47, 0827, 0826);
  lut lut_gate169(0x050c, 0946, 0825, 0893, 0753, 0827);
  lut lut_gate170(0x0e, 0829, 0708, 0754, 0828);
  lut lut_gate171(0x4, 0824, 0946, 0829);
  lut lut_gate172(0x78, 0832, G47, 0831, 0830);
  lut lut_gate173(0x050c, 0946, 0754, 0893, 0753, 0831);
  lut lut_gate174(0xb4, 0814, 0946, 0815, 0832);
  lut lut_gate175(0x807f, 0834, G47, 0832, 0831, 0833);
  lut lut_gate176(0xf40b, 0835, 0822, 0832, 0829, 0834);
  lut lut_gate177(0x4b, 0796, 0836, 0797, 0835);
  lut lut_gate178(0x8, G27, 0947, 0836);
  lut lut_gate179(0x0, 0705, 0838, 0835, 0687, 0837);
  lut lut_gate180(0xe, 0839, 0842, 0838);
  lut lut_gate181(0x3a00, 0840, 0693, G39, G14, 0839);
  lut lut_gate182(0xe000, 0841, 0697, 0692, G13, 0840);
  lut lut_gate183(0xf400, G4, 0700, G12, G40, 0841);
  lut lut_gate184(0x4000, 0846, 0845, 0843, 0844, 0842);
  lut lut_gate185(0x00f1, G4, 0700, G16, G20, 0843);
  lut lut_gate186(0x0b, 0692, G7, G19, 0844);
  lut lut_gate187(0xb0bb, G18, 0693, G17, 0696, 0845);
  lut lut_gate188(0xb0bb, G22, 0695, G21, 0698, 0846);
  lut lut_gate189(0x4100, 0826, 0830, 0828, 0795, 0847);
  lut lut_gate190(0x000, G12, 0849, 0696, G40, 0848);
  lut lut_gate191(0x0, 0850, 0693, G39, 0849);
  lut lut_gate192(0x07, 0692, G14, G10, 0850);
  lut lut_gate193(0x0b, 0692, G8, G20, 0851);
  lut lut_gate194(0xb0bb, G19, 0693, G18, 0696, 0852);
  lut lut_gate195(0xe, 0860, 0853, G3535);
  lut lut_gate196(0xf400, 0855, 0777, 0854, 0847, 0853);
  lut lut_gate197(0x00bf, 0706, 0826, 0833, 0795, 0854);
  lut lut_gate198(0x78, 0857, G47, 0856, 0855);
  lut lut_gate199(0x40, 0831, 0832, 0835, 0856);
  lut lut_gate200(0xf40b, 0859, 0858, 0823, 0836, 0857);
  lut lut_gate201(0x00f4, 0835, 0822, 0832, 0829, 0858);
  lut lut_gate202(0x4b, 0806, 0836, 0807, 0859);
  lut lut_gate203(0x0, 0705, 0861, 0859, 0687, 0860);
  lut lut_gate204(0xf8, 0866, 0869, 0862, 0861);
  lut lut_gate205(0x40, 0865, 0863, G20, 0862);
  lut lut_gate206(0x00f1, 0864, 0692, G18, G22, 0863);
  lut lut_gate207(0x0e, 0700, G19, G15, 0864);
  lut lut_gate208(0x000, G4, G5, 0693, G17, 0865);
  lut lut_gate209(0x40, 0779, 0868, 0867, 0866);
  lut lut_gate210(0x0, 0700, G39, G11, 0867);
  lut lut_gate211(0xeee0, G13, 0693, 0696, G14, 0868);
  lut lut_gate212(0xb0bb, G16, 0696, G21, 0695, 0869);
  lut lut_gate213(0x14eb, 0871, G50, 0870, 0949, G3539);
  lut lut_gate214(0x03a9, 0837, 0860, 0853, 0793, 0870);
  lut lut_gate215(0x96, G3529, 0872, G3536, 0871);
  lut lut_gate216(0x9669, G3528, G3533, G3532, G3531, 0872);
  lut lut_gate217(0x1f, G11, G13, G12, G3520);
  lut lut_gate218(0xb0bb, G32, G9, G33, G10, 0873);
  lut lut_gate219(0x4, G31, G8, 0874);
  lut lut_gate220(0xb0bb, G35, G12, G30, G7, 0875);
  lut lut_gate221(0x0e, G7, G9, G8, 0876);
  lut lut_gate222(0x6, 0878, 0877, G3523);
  lut lut_gate223(0x6996, G8, G10, G9, G7, 0877);
  lut lut_gate224(0x6996, G13, G11, G12, G14, 0878);
  lut lut_gate225(0xb, 0910, 0879, G3525);
  lut lut_gate226(0xef00, 0825, 0737, 0709, 0739, 0879);
  lut lut_gate227(0x7, 0881, 0880, G3537);
  lut lut_gate228(0x0100, 0793, 0860, 0837, 0853, 0880);
  lut lut_gate229(0x1000, 0882, 0883, G3529, G3536, 0881);
  lut lut_gate230(0x1, G3528, G3532, 0882);
  lut lut_gate231(0x1, G3533, G3531, 0883);
  lut lut_gate232(0xe0ff, G27, 0880, G48, 0881, G3538);
  lut lut_gate233(0x0001, G8, G10, G9, G7, G3519);
  lut lut_gate234(0x9, 0885, 0884, G3522);
  lut lut_gate235(0x9669, G30, G31, G33, G32, 0884);
  lut lut_gate236(0x6996, G34, G36, G35, G37, 0885);
  lut lut_gate237(0x4f44, 0708, G1, 0876, 0706, G3527);
  lut lut_gate238(0x728, 0887, 0827, 0856, G47, 0886);
  lut lut_gate239(0x1e, 0795, 0858, 0823, 0887);
  lut lut_gate240(0xef54, G9, G8, G10, G7, 0888);
  lut lut_gate241(0x6, 0871, 0870, G3540);
  lut lut_gate242(0x8, 0825, 0753, G3524);
  lut lut_gate243(0x53fc, 0927, 0705, 0945, 0686, 0889);
  lut lut_gate244(0x5c03, 0889, 0705, G47, 0688, G3528);
  lut lut_gate245(0xaac3, 0705, 0752, 0707, 0923, G3529);
  lut lut_gate246(0xccca, G4, G3, G13, G10, 0890);
  lut lut_gate247(0x0708, 0890, 0930, G12, G3, 0891);
  lut lut_gate248(0xea03, G24, 0724, 0716, 0936, 0892);
  lut lut_gate249(0xe7ff, 0892, 0935, 0730, G24, 0893);
  lut lut_gate250(0x80, 0776, 0775, 0774, 0894);
  lut lut_gate251(0x0bff, 0894, 0692, G12, G40, 0895);
  lut lut_gate252(0x80, 0773, 0772, G8, 0896);
  lut lut_gate253(0x0bff, 0896, 0692, G10, G22, 0897);
  lut lut_gate254(0x80, 0705, 0897, 0895, 0898);
  lut lut_gate255(0xffe0, G26, G3, G25, G24, 0899);
  lut lut_gate256(0xb0ff, 0899, G7, G3, G11, 0900);
  lut lut_gate257(0x0b00, 0705, 0783, 0686, 0760, 0901);
  lut lut_gate258(0x7f00, 0901, 0781, 0779, 0900, 0902);
  lut lut_gate259(0x0b00, 0908, G6, 0686, 0764, 0903);
  lut lut_gate260(0x0f44, 0706, 0903, 0765, 0708, 0904);
  lut lut_gate261(0xb0ef, 0904, 0759, 0706, 0777, G3533);
  lut lut_gate262(0x00f1, G39, 0700, G44, G40, 0905);
  lut lut_gate263(0x0b00, 0792, 0791, G21, 0696, 0906);
  lut lut_gate264(0xf800, 0906, 0692, G7, G11, 0907);
  lut lut_gate265(0x770f, G4, 0907, 0788, 0905, 0908);
  lut lut_gate266(0x07ff, 0796, 0822, 0824, 0814, 0909);
  lut lut_gate267(0x44f0, 0806, 0807, 0909, 0823, 0910);
  lut lut_gate268(0x4f44, 0832, G2, 0848, 0789, 0911);
  lut lut_gate269(0x700, 0926, 0830, 0828, 0777, 0912);
  lut lut_gate270(0x01ff, 0912, 0847, 0794, 0706, G3536);
  lut lut_gate271(0x0, 0875, 0874, G14, G37, 0913);
  lut lut_gate272(0xfacf, G36, 0948, G35, G13, 0914);
  lut lut_gate273(0xccb0, 0948, 0873, G34, G11, 0915);
  lut lut_gate274(0xe000, 0914, 0915, 0913, 0948, 0916);
  lut lut_gate275(0x53cc, 0948, G2, 0916, 0876, G3521);
  lut lut_gate276(0x1c, G2, G1, G3, 0917);
  lut lut_gate277(0x41, G13, G12, G14, 0918);
  lut lut_gate278(0xca, G2, 0918, 0888, 0919);
  lut lut_gate279(0xb217, 0919, 0917, 0886, G2, G3530);
  lut lut_gate280(0xbbb0, 0754, G2, 0755, 0786, 0920);
  lut lut_gate281(0xb000, G9, G7, G20, 0693, 0921);
  lut lut_gate282(0xf100, 0757, 0700, G22, G18, 0922);
  lut lut_gate283(0xf077, G4, 0920, 0922, 0921, 0923);
  lut lut_gate284(0xf100, 0852, 0700, G21, G17, 0924);
  lut lut_gate285(0x0b00, 0924, 0851, G22, 0698, 0925);
  lut lut_gate286(0xcaff, 0705, G4, 0911, 0925, 0926);

endmodule
