module c432(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G426, G427, G428, G429, G430, G431, G432, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, G203, G213, G308, G318, G358;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G5, G6, G7, G8, G9;
  output G426, G427, G428, G429, G430, G431, G432;
  lut lut_gate1(0xbf, 207, 227, 236, G427);
  lut lut_gate2(0x8, 223, 208, 207);
  lut lut_gate3(0x0b, 209, 222, G19, 208);
  lut lut_gate4(0x4, 210, G31, 209);
  lut lut_gate5(0x70, G30, G426, G28, 210);
  lut lut_gate6(0xbf, 211, 216, 221, G426);
  lut lut_gate7(0x8, 214, 212, 211);
  lut lut_gate8(0x0, 213, G1, G2, 212);
  lut lut_gate9(0x4, G6, G4, 213);
  lut lut_gate10(0x0b, 215, G22, G20, 214);
  lut lut_gate11(0x4, G26, G24, 215);
  lut lut_gate12(0x10, 217, 220, 219, 216);
  lut lut_gate13(0x0b, 218, G18, G16, 217);
  lut lut_gate14(0x4, G30, G28, 218);
  lut lut_gate15(0x4, G10, G8, 219);
  lut lut_gate16(0x4, G14, G12, 220);
  lut lut_gate17(0x4, G34, G32, 221);
  lut lut_gate18(0x70, G18, G426, G16, 222);
  lut lut_gate19(0x0b, 224, 226, G15, 223);
  lut lut_gate20(0x4, 225, G11, 224);
  lut lut_gate21(0x70, G10, G426, G8, 225);
  lut lut_gate22(0x70, G14, G426, G12, 226);
  lut lut_gate23(0x8, 232, 228, 227);
  lut lut_gate24(0x0b, 229, 231, G23, 228);
  lut lut_gate25(0x4, 230, G7, 229);
  lut lut_gate26(0x70, G6, G426, G4, 230);
  lut lut_gate27(0x70, G22, G426, G20, 231);
  lut lut_gate28(0x0b, 233, 235, G3, 232);
  lut lut_gate29(0x4, 234, G27, 233);
  lut lut_gate30(0x70, G26, G426, G24, 234);
  lut lut_gate31(0x70, G2, G426, G1, 235);
  lut lut_gate32(0x4, 237, G35, 236);
  lut lut_gate33(0x4, G34, 238, 237);
  lut lut_gate34(0x70, G32, 211, 216, 238);
  lut lut_gate35(0x7f, 250, 246, 239, G428);
  lut lut_gate36(0x01, 244, 242, 240, 239);
  lut lut_gate37(0x4, 241, G17, 240);
  lut lut_gate38(0x70, 226, G427, G15, 241);
  lut lut_gate39(0x4, 243, G13, 242);
  lut lut_gate40(0x70, 225, G427, G11, 243);
  lut lut_gate41(0x4, 245, G9, 244);
  lut lut_gate42(0x70, 230, G427, G7, 245);
  lut lut_gate43(0x0b, 247, 249, G21, 246);
  lut lut_gate44(0x4, 248, G29, 247);
  lut lut_gate45(0x70, 234, G427, G27, 248);
  lut lut_gate46(0x70, 222, G427, G19, 249);
  lut lut_gate47(0x10, 253, 257, 251, 250);
  lut lut_gate48(0x4, 252, G33, 251);
  lut lut_gate49(0x70, 210, G427, G31, 252);
  lut lut_gate50(0x0b, 255, 254, G5, 253);
  lut lut_gate51(0x70, 235, G427, G3, 254);
  lut lut_gate52(0x10, 237, G36, 256, 255);
  lut lut_gate53(0x70, G35, 207, 227, 256);
  lut lut_gate54(0x4, 258, G25, 257);
  lut lut_gate55(0x70, 231, G427, G23, 258);
  lut lut_gate56(0x0, 203, G430, 198, G429);
  lut lut_gate57(0xb, 193, 197, G430);
  lut lut_gate58(0x10, 195, 196, 194, 193);
  lut lut_gate59(0x70, 241, G428, G17, 194);
  lut lut_gate60(0x8f, 249, G21, G428, 195);
  lut lut_gate61(0x70, 243, G428, G13, 196);
  lut lut_gate62(0x70, 245, G428, G9, 197);
  lut lut_gate63(0x4, 199, 202, 198);
  lut lut_gate64(0x01, G34, 201, 200, 199);
  lut lut_gate65(0x70, 252, G428, G33, 200);
  lut lut_gate66(0x70, 248, G428, G29, 201);
  lut lut_gate67(0x70, 258, G428, G25, 202);
  lut lut_gate68(0x70, 254, G428, G5, 203);
  lut lut_gate69(0xef, 204, 196, 205, G431);
  lut lut_gate70(0x07, 197, 193, 202, 204);
  lut lut_gate71(0x40, 201, 195, 194, 205);
  lut lut_gate72(0x1f, 204, 196, 206, G432);
  lut lut_gate73(0x0b, 194, 200, 201, 206);

endmodule
