module c880(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G7, G8, G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878, G879, G880, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, G293, G295, G296, G343, G349, G350, G369, G812, G829, G830, G831, G832, G844, G849, G850, G851;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G7, G8, G9;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878, G879, G880;
  lut lut_gate1(0x7f, G6, G16, G8, G855);
  lut lut_gate2(0x7f, G7, G17, G6, G856);
  lut lut_gate3(0x7f, G7, G6, G8, G857);
  lut lut_gate4(0x7, G18, G19, G858);
  lut lut_gate5(0x7, G3, 411, G859);
  lut lut_gate6(0x80, G1, G2, G4, 411);
  lut lut_gate7(0x8, G857, 412, G860);
  lut lut_gate8(0x8, G3, 413, 412);
  lut lut_gate9(0x80, G5, G1, G4, 413);
  lut lut_gate10(0x1f, G23, G21, G20, G864);
  lut lut_gate11(0x4, 412, G857, G865);
  lut lut_gate12(0x7f, G9, G5, G1, G866);
  lut lut_gate13(0x1f, G22, G21, G20, G869);
  lut lut_gate14(0x4, 296, 321, G872);
  lut lut_gate15(0x70, 297, 320, G52, 296);
  lut lut_gate16(0x8, 313, 298, 297);
  lut lut_gate17(0x0e, 311, 299, 312, 298);
  lut lut_gate18(0x01, 309, 306, 300, 299);
  lut lut_gate19(0xe0, G31, 301, 304, 300);
  lut lut_gate20(0x10, 303, 302, G866, 301);
  lut lut_gate21(0x9, G4, G8, 302);
  lut lut_gate22(0x8, G11, G40, 303);
  lut lut_gate23(0x40, G9, 411, 305, 304);
  lut lut_gate24(0x80, G11, G16, G8, 305);
  lut lut_gate25(0x40, 307, G10, G60, 306);
  lut lut_gate26(0x4, 308, G866, 307);
  lut lut_gate27(0x80, G17, G6, G16, 308);
  lut lut_gate28(0x0, G39, 310, G1, 309);
  lut lut_gate29(0x10, G4, 303, G866, 310);
  lut lut_gate30(0x8, G50, G30, 311);
  lut lut_gate31(0x07, G54, G48, G53, 312);
  lut lut_gate32(0x07, 319, 314, G48, 313);
  lut lut_gate33(0x80, 318, 317, 315, 314);
  lut lut_gate34(0x80, G10, G3, 316, 315);
  lut lut_gate35(0x8, G1, G2, 316);
  lut lut_gate36(0x8, G12, G11, 317);
  lut lut_gate37(0x80, G14, G13, G8, 318);
  lut lut_gate38(0x8, G55, G59, 319);
  lut lut_gate39(0x9, G48, 299, 320);
  lut lut_gate40(0x60, G51, G58, 320, 321);
  lut lut_gate41(0x40, 338, 336, 322, G873);
  lut lut_gate42(0x90, G51, 333, 323, 322);
  lut lut_gate43(0xb2, 329, G46, 324, 323);
  lut lut_gate44(0x71, 326, G47, 325, 324);
  lut lut_gate45(0x4, G58, G48, 299, 325);
  lut lut_gate46(0x01, 328, 327, 306, 326);
  lut lut_gate47(0x0, G37, 310, G1, 327);
  lut lut_gate48(0xe0, G30, 301, 304, 328);
  lut lut_gate49(0x0, 330, 332, G36, 329);
  lut lut_gate50(0x0, 306, 331, G29, 330);
  lut lut_gate51(0x1, 304, 301, 331);
  lut lut_gate52(0x4, G1, 310, 332);
  lut lut_gate53(0x9, G45, 334, 333);
  lut lut_gate54(0x0, 335, 332, G35, 334);
  lut lut_gate55(0x0, 306, 331, G28, 335);
  lut lut_gate56(0x07, 337, 333, G52, 336);
  lut lut_gate57(0x4, G54, 334, 337);
  lut lut_gate58(0x0, 340, 339, G45, 338);
  lut lut_gate59(0x0, 314, 334, G53, 339);
  lut lut_gate60(0x8, G27, G50, 340);
  lut lut_gate61(0x10, 343, 348, 341, G874);
  lut lut_gate62(0x90, G51, 342, 324, 341);
  lut lut_gate63(0x9, G46, 329, 342);
  lut lut_gate64(0x70, 344, 342, G52, 343);
  lut lut_gate65(0x0, 345, 329, G54, 344);
  lut lut_gate66(0x70, 346, 314, G46, 345);
  lut lut_gate67(0x07, 347, G55, G56, 346);
  lut lut_gate68(0x8, G28, G50, 347);
  lut lut_gate69(0x40, G46, G53, 329, 348);
  lut lut_gate70(0x8, G52, 350, 349);
  lut lut_gate71(0x9, G47, 326, 350);
  lut lut_gate72(0x70, 352, 314, G47, 351);
  lut lut_gate73(0x07, 353, G50, G29, 352);
  lut lut_gate74(0x8, G57, G55, 353);
  lut lut_gate75(0x60, G51, 350, 325, 354);
  lut lut_gate76(0xb2, 370, G41, 355, G876);
  lut lut_gate77(0xb2, 367, G42, 356, 355);
  lut lut_gate78(0xb2, 364, G43, 357, 356);
  lut lut_gate79(0xb2, 359, G44, 358, 357);
  lut lut_gate80(0xb2, 334, G45, 323, 358);
  lut lut_gate81(0x0, 360, 331, G27, 359);
  lut lut_gate82(0x70, 361, 363, G39, 360);
  lut lut_gate83(0x07, 362, G34, G38, 361);
  lut lut_gate84(0x40, 307, G4, G60, 362);
  lut lut_gate85(0x10, G10, 303, G866, 363);
  lut lut_gate86(0x0, 365, 331, G26, 364);
  lut lut_gate87(0x70, 366, 363, G37, 365);
  lut lut_gate88(0x07, 362, G4, G34, 366);
  lut lut_gate89(0x0, 368, 331, G25, 367);
  lut lut_gate90(0x70, 369, 363, G36, 368);
  lut lut_gate91(0x07, 362, G9, G34, 369);
  lut lut_gate92(0x0, 371, 331, G24, 370);
  lut lut_gate93(0x70, 372, 363, G35, 371);
  lut lut_gate94(0x07, 362, G2, G34, 372);
  lut lut_gate95(0x90, G51, 374, 358, 373);
  lut lut_gate96(0x9, G44, 359, 374);
  lut lut_gate97(0x8, G52, 374, 375);
  lut lut_gate98(0x8, G26, G50, 376);
  lut lut_gate99(0x4, 379, 377, G878);
  lut lut_gate100(0x90, G51, 378, 355, 377);
  lut lut_gate101(0x9, G41, 370, 378);
  lut lut_gate102(0x70, 410, 378, G52, 379);
  lut lut_gate103(0x07, 381, 314, G41, 380);
  lut lut_gate104(0x8, G60, G50, 381);
  lut lut_gate105(0x4, 384, 382, G879);
  lut lut_gate106(0x90, G51, 383, 356, 382);
  lut lut_gate107(0x9, G42, 367, 383);
  lut lut_gate108(0x70, 385, 383, G52, 384);
  lut lut_gate109(0x70, 386, 314, G42, 385);
  lut lut_gate110(0x0e, 387, 367, 388, 386);
  lut lut_gate111(0x8, G24, G50, 387);
  lut lut_gate112(0x07, G54, G53, G42, 388);
  lut lut_gate113(0x4, 391, 389, G880);
  lut lut_gate114(0x90, G51, 390, 357, 389);
  lut lut_gate115(0x9, G43, 364, 390);
  lut lut_gate116(0x70, 392, 390, G52, 391);
  lut lut_gate117(0x70, 393, 314, G43, 392);
  lut lut_gate118(0x0e, 394, 364, 395, 393);
  lut lut_gate119(0x8, G25, G50, 394);
  lut lut_gate120(0x07, G54, G53, G43, 395);
  lut lut_gate121(0x80, G11, G17, G16, G861);
  lut lut_gate122(0x80, G11, G7, G17, G862);
  lut lut_gate123(0x80, G11, G7, G8, G863);
  lut lut_gate124(0x7f, G12, G6, 315, G867);
  lut lut_gate125(0x7f, G15, 317, 315, G868);
  lut lut_gate126(0x69, 399, 398, 396, G870);
  lut lut_gate127(0x96, G31, G30, 397, 396);
  lut lut_gate128(0x9, G24, G27, 397);
  lut lut_gate129(0x69, G32, G26, G25, 398);
  lut lut_gate130(0x96, G33, G29, G28, 399);
  lut lut_gate131(0x69, 403, 402, 400, G871);
  lut lut_gate132(0x96, G45, G48, 401, 400);
  lut lut_gate133(0x9, G42, G41, 401);
  lut lut_gate134(0x96, G32, G44, G43, 402);
  lut lut_gate135(0x69, G49, G47, G46, 403);
  lut lut_gate136(0xf8, G54, G47, G53, 404);
  lut lut_gate137(0xb0, 351, 404, 326, 405);
  lut lut_gate138(0x10, 405, 354, 349, G875);
  lut lut_gate139(0xf8, G54, G44, G53, 406);
  lut lut_gate140(0x01, 376, 375, 373, 407);
  lut lut_gate141(0x70, 407, G44, 314, 408);
  lut lut_gate142(0xb0, 408, 406, 359, G877);
  lut lut_gate143(0xf8, G54, G41, G53, 409);
  lut lut_gate144(0xb0, 380, 409, 370, 410);

endmodule
