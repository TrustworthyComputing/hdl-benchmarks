module c3540(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, 0950, 0951, 0952, 0953, 0954, 0955, 0956, 0957, 0958, 0959, 0960, 0961, 0962, 0963, 0964, 0965, 0966, 0967, 0968, 0969, 0970, 0971, 0972, 0973, 0974, 0975, 0976, 0977, 0978, 0979, 0980, 0981, 0982, 0983, 0984, 0985, 0986, 0987, 0988, 0989, 0990, 0991, 0992, 0993, 0994, 0995, 0996, 0997, 0998, 0999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165, 1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 1178, 1179, G1022, G2943, G2974, G2985, G3005, G3030, G3100, G3135, G3195, G3202, G3226, G3257, G3265, G3266, G3267, G3275, G3281, G3294, G3300, G3301, G3311, G3312, G3320, G3332, G3341, G3342, G3343, G3345, G3373, G3376, G3379, G3394, G3515, G3516, G722, G723, G724, G725, G731, G734, G735, G736, G739, G742, G745, G749, G781, G786, G791, G792, G793, G794, G795, G796, G797, G798, G799, G816, G831, G882, G883, G890, G891, G892, G893, G894, G897, G898, G901, G904, G907, G910, G913, G916, G919, G922, G925;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540;
  lut lut_gate1(0x9, 0742, 1002, 0997);
  lut lut_gate2(0x4, 0694, 1005, 1013);
  lut lut_gate3(0x1, 1130, 1007, 1042);
  lut lut_gate4(0x1, 1088, 1070, 1063);
  lut lut_gate5(0x8, G4, 1078, 1070);
  lut lut_gate6(0x8, G3, G1, 1078);
  lut lut_gate7(0x8, G1, G2, 1088);
  lut lut_gate8(0x8, G3, 1113, 1104);
  lut lut_gate9(0x4, G2, G1, 1113);
  lut lut_gate10(0x4, G3, 1063, 1130);
  lut lut_gate11(0x4, 1088, G3, 1173);
  lut lut_gate12(0x4, 1010, 0739, 0694);
  lut lut_gate13(0x4, G37, 0732, 0731);
  lut lut_gate14(0x4, 0733, G5, 0732);
  lut lut_gate15(0x1, G6, G1, 0733);
  lut lut_gate16(0x8, G35, 0735, 0734);
  lut lut_gate17(0x1, G49, G4, 0735);
  lut lut_gate18(0x4, 1088, 0737, 0736);
  lut lut_gate19(0x8, G5, G4, 0737);
  lut lut_gate20(0x8, 0732, G38, 0738);
  lut lut_gate21(0x1, G24, G23, 0739);
  lut lut_gate22(0x4, 1010, 0741, 0740);
  lut lut_gate23(0x1, G26, G25, 0741);
  lut lut_gate24(0x4, 0743, 1005, 0742);
  lut lut_gate25(0x8, 0746, 0744, 0743);
  lut lut_gate26(0x4, 0745, G3, 0744);
  lut lut_gate27(0x1, G1, G2, 0745);
  lut lut_gate28(0x8, G48, G27, 0746);
  lut lut_gate29(0x4, 0748, G6, 0747);
  lut lut_gate30(0x8, G5, 0744, 0748);
  lut lut_gate31(0x4, 0750, G2, 0749);
  lut lut_gate32(0x4, G4, G3, 0750);
  lut lut_gate33(0x1, G13, 0752, 0751);
  lut lut_gate34(0x8, G25, 0753, 0752);
  lut lut_gate35(0x4, 0754, G24, 0753);
  lut lut_gate36(0x8, G26, G3, 0754);
  lut lut_gate37(0x4, 1017, G26, 0755);
  lut lut_gate38(0x8, G25, G3, 0756);
  lut lut_gate39(0x1, G7, 0758, 0757);
  lut lut_gate40(0x8, G26, 1017, 0758);
  lut lut_gate41(0x4, 1017, 0754, 0759);
  lut lut_gate42(0x1, 0763, 0761, 0760);
  lut lut_gate43(0x1, G11, 0762, 0761);
  lut lut_gate44(0x4, 0753, G25, 0762);
  lut lut_gate45(0x1, G9, 0752, 0763);
  lut lut_gate46(0x8, 0765, 0756, 0764);
  lut lut_gate47(0x1, G26, G24, 0765);
  lut lut_gate48(0x4, G41, 0762, 0766);
  lut lut_gate49(0x1, 0768, 0752, 0767);
  lut lut_gate50(0x1, G43, G39, 0768);
  lut lut_gate51(0x4, G44, 0755, 0769);
  lut lut_gate52(0x1, G46, G42, 0770);
  lut lut_gate53(0x1, 0794, 0772, 0771);
  lut lut_gate54(0x1, 0743, 1174, 0772);
  lut lut_gate55(0x8, 1048, 0774, 0773);
  lut lut_gate56(0x8, 0782, 1027, 0774);
  lut lut_gate57(0x4, 0778, 1032, 0775);
  lut lut_gate58(0x1, G10, G4, 0776);
  lut lut_gate59(0x6, G13, G12, 0777);
  lut lut_gate60(0x4, 0779, 0739, 0778);
  lut lut_gate61(0x1, 0738, 1035, 0779);
  lut lut_gate62(0x4, G35, 0732, 0780);
  lut lut_gate63(0x4, 0779, 0741, 0781);
  lut lut_gate64(0x1, 0786, 0783, 0782);
  lut lut_gate65(0x4, 0785, 1043, 0783);
  lut lut_gate66(0x1, G13, G12, 0784);
  lut lut_gate67(0x1, 0739, 1047, 0785);
  lut lut_gate68(0x4, 1043, 0787, 0786);
  lut lut_gate69(0x1, 0741, 1047, 0787);
  lut lut_gate70(0x4, 0789, 1054, 0788);
  lut lut_gate71(0x4, 0790, 0739, 0789);
  lut lut_gate72(0x1, 0738, 1051, 0790);
  lut lut_gate73(0x4, G36, 0732, 0791);
  lut lut_gate74(0x1, G2, 1070, 0792);
  lut lut_gate75(0x4, 0790, 0741, 0793);
  lut lut_gate76(0x9, 0804, 1057, 0794);
  lut lut_gate77(0x4, 0798, 1061, 0795);
  lut lut_gate78(0x4, 1063, 0797, 0796);
  lut lut_gate79(0x4, G3, G1, 0797);
  lut lut_gate80(0x4, 1065, 0739, 0798);
  lut lut_gate81(0x4, G33, 0800, 0799);
  lut lut_gate82(0x1, 0732, G1, 0800);
  lut lut_gate83(0x8, G31, 0735, 0801);
  lut lut_gate84(0x8, 0800, G38, 0802);
  lut lut_gate85(0x4, 1065, 0741, 0803);
  lut lut_gate86(0x4, 0743, 1061, 0804);
  lut lut_gate87(0x4, G47, 1066, 0805);
  lut lut_gate88(0x8, 1002, 0773, 0806);
  lut lut_gate89(0x4, G4, G2, 0807);
  lut lut_gate90(0x1, 0809, 0752, 0808);
  lut lut_gate91(0x4, G11, G39, 0809);
  lut lut_gate92(0x1, G13, 0762, 0810);
  lut lut_gate93(0x4, G14, G42, 0811);
  lut lut_gate94(0x4, G20, 0755, 0812);
  lut lut_gate95(0x1, G18, G22, 0813);
  lut lut_gate96(0x1, G7, 0762, 0814);
  lut lut_gate97(0x9, 0816, 1048, 0815);
  lut lut_gate98(0x4, 0743, 1054, 0816);
  lut lut_gate99(0x8, G47, 0997, 0817);
  lut lut_gate100(0x6, G3526, 0819, 0818);
  lut lut_gate101(0x9, 0820, 1079, 0819);
  lut lut_gate102(0x9, 0821, 1027, 0820);
  lut lut_gate103(0x4, 0743, 1032, 0821);
  lut lut_gate104(0x8, 0815, 0822, G3526);
  lut lut_gate105(0x4, G47, 0997, 0822);
  lut lut_gate106(0x4, 0824, 0797, 0823);
  lut lut_gate107(0x1, 0733, 1113, 0824);
  lut lut_gate108(0x4, 0775, 0743, 0825);
  lut lut_gate109(0x6, 0827, 0782, 0826);
  lut lut_gate110(0x4, 0743, 1043, 0827);
  lut lut_gate111(0x8, 0749, 0826, 0828);
  lut lut_gate112(0x4, G21, 0755, 0829);
  lut lut_gate113(0x1, 0832, 0831, 0830);
  lut lut_gate114(0x1, G8, 0762, 0831);
  lut lut_gate115(0x1, 0833, 0752, 0832);
  lut lut_gate116(0x4, G10, G22, 0833);
  lut lut_gate117(0x1, 0835, 0764, 0834);
  lut lut_gate118(0x4, G7, G19, 0835);
  lut lut_gate119(0x1, 0768, 0764, 0836);
  lut lut_gate120(0x1, 0839, 0838, 0837);
  lut lut_gate121(0x1, G14, 0762, 0838);
  lut lut_gate122(0x4, G42, 0758, 0839);
  lut lut_gate123(0x1, 0841, 0752, 0840);
  lut lut_gate124(0x4, G12, G40, 0841);
  lut lut_gate125(0x4, 0691, 0772, 0842);
  lut lut_gate126(0x4, 0749, 0815, 0843);
  lut lut_gate127(0x1, G11, 0759, 0844);
  lut lut_gate128(0x1, 0847, 0846, 0845);
  lut lut_gate129(0x4, G22, 0758, 0846);
  lut lut_gate130(0x1, 0848, 0764, 0847);
  lut lut_gate131(0x4, G9, G21, 0848);
  lut lut_gate132(0x1, G10, 0762, 0849);
  lut lut_gate133(0x4, G44, 0758, 0850);
  lut lut_gate134(0x1, 0853, 0852, 0851);
  lut lut_gate135(0x4, G39, 0759, 0852);
  lut lut_gate136(0x1, 0811, 0752, 0853);
  lut lut_gate137(0x4, 0856, 0855, 0854);
  lut lut_gate138(0x4, G40, 0762, 0855);
  lut lut_gate139(0x4, G4, 0857, 0856);
  lut lut_gate140(0x1, 0858, 0764, 0857);
  lut lut_gate141(0x1, G45, G41, 0858);
  lut lut_gate142(0x4, 0749, 0820, 0859);
  lut lut_gate143(0x1, G9, 0762, 0860);
  lut lut_gate144(0x1, G10, 0759, 0861);
  lut lut_gate145(0x1, 0864, 0863, 0862);
  lut lut_gate146(0x4, G21, 0758, 0863);
  lut lut_gate147(0x1, 0865, 0764, 0864);
  lut lut_gate148(0x4, G8, G20, 0865);
  lut lut_gate149(0x1, 0867, 0752, 0866);
  lut lut_gate150(0x4, G13, G41, 0867);
  lut lut_gate151(0x1, 0870, 0869, 0868);
  lut lut_gate152(0x1, G14, 0759, 0869);
  lut lut_gate153(0x4, G43, 0758, 0870);
  lut lut_gate154(0x4, 0873, 0872, 0871);
  lut lut_gate155(0x4, G39, 0762, 0872);
  lut lut_gate156(0x4, G4, 0874, 0873);
  lut lut_gate157(0x1, 0875, 0764, 0874);
  lut lut_gate158(0x1, G44, G40, 0875);
  lut lut_gate159(0x1, 0726, 0877, 0876);
  lut lut_gate160(0x9, 0886, 0878, 0877);
  lut lut_gate161(0x6, 0881, 0879, 0878);
  lut lut_gate162(0x8, G47, 0880, 0879);
  lut lut_gate163(0x4, 1066, 0794, 0880);
  lut lut_gate164(0x6, 0885, 1109, 0881);
  lut lut_gate165(0x4, 0883, 1116, 0882);
  lut lut_gate166(0x4, 1111, 0739, 0883);
  lut lut_gate167(0x4, 1111, 0741, 0884);
  lut lut_gate168(0x4, 0743, 1116, 0885);
  lut lut_gate169(0x1, 0887, 0771, 0886);
  lut lut_gate170(0x4, 0795, 0743, 0887);
  lut lut_gate171(0x4, 0708, 0889, 0888);
  lut lut_gate172(0x1, 0890, 0772, 0889);
  lut lut_gate173(0x8, 1057, 0891, 0890);
  lut lut_gate174(0x8, 1109, 0892, 0891);
  lut lut_gate175(0x8, 0898, 1119, 0892);
  lut lut_gate176(0x4, 0894, 1125, 0893);
  lut lut_gate177(0x4, 1128, 0739, 0894);
  lut lut_gate178(0x4, G31, 0800, 0895);
  lut lut_gate179(0x8, G29, 0735, 0896);
  lut lut_gate180(0x4, 1128, 0741, 0897);
  lut lut_gate181(0x1, 0902, 0899, 0898);
  lut lut_gate182(0x4, 0901, 0706, 0899);
  lut lut_gate183(0x1, G8, G9, 0900);
  lut lut_gate184(0x4, 1133, 0739, 0901);
  lut lut_gate185(0x4, 0706, 0903, 0902);
  lut lut_gate186(0x4, 1133, 0741, 0903);
  lut lut_gate187(0x9, 0906, 0905, 0904);
  lut lut_gate188(0x8, 0881, 0879, 0905);
  lut lut_gate189(0x6, 0909, 0907, 0906);
  lut lut_gate190(0x1, 0882, 0908, 0907);
  lut lut_gate191(0x4, 0881, 0887, 0908);
  lut lut_gate192(0x9, 0910, 1119, 0909);
  lut lut_gate193(0x4, 0911, 1125, 0910);
  lut lut_gate194(0x8, G27, 0744, 0911);
  lut lut_gate195(0x4, 0807, 0909, 0912);
  lut lut_gate196(0x1, G14, 0755, 0913);
  lut lut_gate197(0x1, 0916, 0915, 0914);
  lut lut_gate198(0x1, 0835, 0752, 0915);
  lut lut_gate199(0x4, G21, 0762, 0916);
  lut lut_gate200(0x1, G16, G20, 0917);
  lut lut_gate201(0x8, 0807, 0881, 0918);
  lut lut_gate202(0x4, G18, 0758, 0919);
  lut lut_gate203(0x1, G17, G21, 0920);
  lut lut_gate204(0x4, G22, 0762, 0921);
  lut lut_gate205(0x1, 0865, 0752, 0922);
  lut lut_gate206(0x8, 0927, 0924, 0923);
  lut lut_gate207(0x1, 0926, 0925, 0924);
  lut lut_gate208(0x4, G40, 0758, 0925);
  lut lut_gate209(0x1, G12, 0762, 0926);
  lut lut_gate210(0x1, 0929, 0928, 0927);
  lut lut_gate211(0x4, G39, 0755, 0928);
  lut lut_gate212(0x1, 0930, 0752, 0929);
  lut lut_gate213(0x8, G10, G14, 0930);
  lut lut_gate214(0x6, 0935, 0932, 0931);
  lut lut_gate215(0x8, G47, 0933, 0932);
  lut lut_gate216(0x8, 0934, 0880, 0933);
  lut lut_gate217(0x4, 0881, 0909, 0934);
  lut lut_gate218(0x6, 0939, 0936, 0935);
  lut lut_gate219(0x1, 0938, 0937, 0936);
  lut lut_gate220(0x1, 0909, 0907, 0937);
  lut lut_gate221(0x4, 0893, 0911, 0938);
  lut lut_gate222(0x9, 0940, 0898, 0939);
  lut lut_gate223(0x4, 0911, 0706, 0940);
  lut lut_gate224(0x1, 0813, 0752, 0941);
  lut lut_gate225(0x4, G20, 0762, 0942);
  lut lut_gate226(0x1, 0944, 0764, 0943);
  lut lut_gate227(0x1, G15, G19, 0944);
  lut lut_gate228(0x4, G5, 0946, 0945);
  lut lut_gate229(0x1, 0809, 0764, 0946);
  lut lut_gate230(0x1, G14, 0758, 0947);
  lut lut_gate231(0x9, 0951, 0948, G3539);
  lut lut_gate232(0x4, 0949, 0746, 0948);
  lut lut_gate233(0x6, G50, 0950, 0949);
  lut lut_gate234(0x6, G3534, G3535, 0950);
  lut lut_gate235(0x6, 0953, 0952, 0951);
  lut lut_gate236(0x6, G3529, G3536, 0952);
  lut lut_gate237(0x9, 0955, 0954, 0953);
  lut lut_gate238(0x6, G3533, G3531, 0954);
  lut lut_gate239(0x6, G3528, G3532, 0955);
  lut lut_gate240(0xb, G11, 0784, G3520);
  lut lut_gate241(0x8, 0960, 0957, 0956);
  lut lut_gate242(0x1, 0959, 0958, 0957);
  lut lut_gate243(0x4, G32, G9, 0958);
  lut lut_gate244(0x4, G33, G10, 0959);
  lut lut_gate245(0x1, 0962, 0961, 0960);
  lut lut_gate246(0x4, G36, G13, 0961);
  lut lut_gate247(0x4, G31, G8, 0962);
  lut lut_gate248(0x1, 0965, 0964, 0963);
  lut lut_gate249(0x4, G35, G12, 0964);
  lut lut_gate250(0x4, G30, G7, 0965);
  lut lut_gate251(0x4, G37, G14, 0966);
  lut lut_gate252(0x1, G3, G1, 0967);
  lut lut_gate253(0x8, 0970, 0969, 0968);
  lut lut_gate254(0x4, 1113, G3, 0969);
  lut lut_gate255(0x1, G7, 0900, 0970);
  lut lut_gate256(0x1, G36, G35, 0971);
  lut lut_gate257(0x6, 0975, 0972, G3523);
  lut lut_gate258(0x9, 0974, 0973, 0972);
  lut lut_gate259(0x6, G10, G9, 0973);
  lut lut_gate260(0x9, G8, G7, 0974);
  lut lut_gate261(0x9, 0977, 0976, 0975);
  lut lut_gate262(0x9, G12, G14, 0976);
  lut lut_gate263(0x6, G13, G11, 0977);
  lut lut_gate264(0xb, 0708, 0978, G3525);
  lut lut_gate265(0x4, 0890, 1174, 0978);
  lut lut_gate266(0x7, 0980, 0979, G3537);
  lut lut_gate267(0x1, G3534, G3535, 0979);
  lut lut_gate268(0x8, 0982, 0981, 0980);
  lut lut_gate269(0x1, G3529, G3536, 0981);
  lut lut_gate270(0x8, 0984, 0983, 0982);
  lut lut_gate271(0x1, G3533, G3531, 0983);
  lut lut_gate272(0x1, G3528, G3532, 0984);
  lut lut_gate273(0xb, G27, 0985, G3538);
  lut lut_gate274(0x4, 0979, 0986, 0985);
  lut lut_gate275(0x1, G48, 0980, 0986);
  lut lut_gate276(0x8, 0987, 0900, G3519);
  lut lut_gate277(0x1, G10, G7, 0987);
  lut lut_gate278(0x9, 0991, 0988, G3522);
  lut lut_gate279(0x6, 0990, 0989, 0988);
  lut lut_gate280(0x6, G30, G31, 0989);
  lut lut_gate281(0x9, G33, G32, 0990);
  lut lut_gate282(0x9, 0993, 0992, 0991);
  lut lut_gate283(0x6, G34, G36, 0992);
  lut lut_gate284(0x9, G35, G37, 0993);
  lut lut_gate285(0xe, 0995, 0994, G3527);
  lut lut_gate286(0x4, 0772, G1, 0994);
  lut lut_gate287(0x4, 0970, 0748, 0995);
  lut lut_gate288(0x9, 0936, 0888, 0996);
  lut lut_gate289(0x4, 0999, 0777, 0998);
  lut lut_gate290(0x4, 0969, G14, 0999);
  lut lut_gate291(0x6, 0951, 0950, G3540);
  lut lut_gate292(0x8, 0890, 0806, G3524);
  lut lut_gate293(0xac, 0747, G47, 0749, 1000);
  lut lut_gate294(0x9e, 1000, 0747, 0997, 1001);
  lut lut_gate295(0xb0, 1001, 0747, 1016, G3528);
  lut lut_gate296(0xc5, 1005, 0740, 0694, 1002);
  lut lut_gate297(0xc5, G14, 1042, 1104, 1003);
  lut lut_gate298(0xc5, G4, G39, G12, 1004);
  lut lut_gate299(0x70, 1003, 1004, 1173, 1005);
  lut lut_gate300(0x4f, G4, G1, 1078, 1006);
  lut lut_gate301(0x10, 1006, 1104, 1088, 1007);
  lut lut_gate302(0x35, G4, G36, G41, 1008);
  lut lut_gate303(0xef, 1008, 0734, 0731, 1009);
  lut lut_gate304(0x0b, 0738, 1009, 0736, 1010);
  lut lut_gate305(0x4, 1021, 0769, 1011);
  lut lut_gate306(0xca, G4, 1011, 1171, 1012);
  lut lut_gate307(0x4, G10, G22, 1014);
  lut lut_gate308(0x35, G4, 0770, 1014, 1015);
  lut lut_gate309(0x4f, 1012, 1015, 0764, 1016);
  lut lut_gate310(0x1f, G3, G25, G24, 1017);
  lut lut_gate311(0x8f, G45, 1017, G26, 1018);
  lut lut_gate312(0x4f, G40, 1017, 0754, 1019);
  lut lut_gate313(0x1, 0767, 0766, 1020);
  lut lut_gate314(0x80, 1020, 1019, 1018, 1021);
  lut lut_gate315(0xc5, 0747, 0807, 0772, 1022);
  lut lut_gate316(0xca, 0747, 1071, 0805, 1023);
  lut lut_gate317(0x43, 1023, 0747, 1022, 1024);
  lut lut_gate318(0x4b, 1057, 1022, 0804, 1025);
  lut lut_gate319(0xca, 1025, 1024, 1023, G3529);
  lut lut_gate320(0xf8, 0788, 1013, 1048, 1026);
  lut lut_gate321(0xc5, 1032, 0781, 0778, 1027);
  lut lut_gate322(0xc5, G13, G3, 0750, 1028);
  lut lut_gate323(0xc5, G3, G12, 0776, 1029);
  lut lut_gate324(0x68, G13, 1029, 1028, 1030);
  lut lut_gate325(0x35, G12, 1007, 1104, 1031);
  lut lut_gate326(0xb0, 1031, 1030, 1063, 1032);
  lut lut_gate327(0x0, G39, G49, G33, 1033);
  lut lut_gate328(0x3a, G4, G34, 1033, 1034);
  lut lut_gate329(0x0b, 0736, 1034, 0780, 1035);
  lut lut_gate330(0xca, G4, G12, G9, 1036);
  lut lut_gate331(0x3a, G11, 1007, 0784, 1037);
  lut lut_gate332(0xc5, G11, 1037, 1104, 1038);
  lut lut_gate333(0xe0, 1038, 1036, 1063, 1039);
  lut lut_gate334(0x4, 1037, 1063, G11, 1040);
  lut lut_gate335(0x0, 1040, G11, 1104, 1041);
  lut lut_gate336(0xca, G3, 1041, 1039, 1043);
  lut lut_gate337(0x0, G14, G49, G32, 1044);
  lut lut_gate338(0x5c, G4, 1044, G33, 1045);
  lut lut_gate339(0x35, 0733, G38, G34, 1046);
  lut lut_gate340(0x07, 0736, 1045, 1046, 1047);
  lut lut_gate341(0xa3, 1054, 0789, 0793, 1048);
  lut lut_gate342(0x0, G40, G49, G34, 1049);
  lut lut_gate343(0x3a, G4, G35, 1049, 1050);
  lut lut_gate344(0x0b, 0736, 1050, 0791, 1051);
  lut lut_gate345(0x4, G3, 0792, 1052);
  lut lut_gate346(0x53, G13, 1052, 1007, 1053);
  lut lut_gate347(0x4, 1053, 1056, 1054);
  lut lut_gate348(0xc5, G4, G14, G11, 1055);
  lut lut_gate349(0x8, 1173, 1055, 1056);
  lut lut_gate350(0xc5, 1061, 0803, 0798, 1057);
  lut lut_gate351(0xca, G4, G11, G8, 1058);
  lut lut_gate352(0xc5, G3, G10, 1058, 1059);
  lut lut_gate353(0x35, G10, 0796, 1104, 1060);
  lut lut_gate354(0xb0, 1060, 1059, 1063, 1061);
  lut lut_gate355(0x35, G4, G32, G13, 1062);
  lut lut_gate356(0xef, 1062, 0801, 0799, 1064);
  lut lut_gate357(0x0b, 0802, 1064, 0736, 1065);
  lut lut_gate358(0x3a, 0743, 0806, 1068, 1066);
  lut lut_gate359(0x18, 1010, 1047, G24, 1067);
  lut lut_gate360(0x7, 1067, 1176, 1068);
  lut lut_gate361(0x35, G4, 0811, 0813, 1069);
  lut lut_gate362(0x4f, 0689, 1069, 0764, 1071);
  lut lut_gate363(0x0, 0825, 1079, 0820, 1072);
  lut lut_gate364(0x78, 0826, G3526, 0820, 1073);
  lut lut_gate365(0xeb, 1073, 1072, 1076, 1074);
  lut lut_gate366(0xb, 1074, 1082, G3531);
  lut lut_gate367(0x8f, 0772, 0818, 0691, 1075);
  lut lut_gate368(0x0, 0823, 0748, 1075, 1076);
  lut lut_gate369(0x4f, 0815, 1013, 0743, 1077);
  lut lut_gate370(0x0, 1077, 0743, 0788, 1079);
  lut lut_gate371(0x40, 1085, 0837, 0840, 1080);
  lut lut_gate372(0x35, G4, 1080, 0696, 1081);
  lut lut_gate373(0x40, 1081, 0747, 0828, 1082);
  lut lut_gate374(0x4f, G41, 1017, G26, 1083);
  lut lut_gate375(0xf4, G13, 1017, 0754, 1084);
  lut lut_gate376(0x40, 1083, 1084, 0836, 1085);
  lut lut_gate377(0x10, 1094, 0843, G6, 1086);
  lut lut_gate378(0x3a, 0748, 1086, 0772, 1087);
  lut lut_gate379(0x87, 1087, 0691, 0748, 1089);
  lut lut_gate380(0xbc, 0691, 1089, 0823, G3532);
  lut lut_gate381(0x40, 0698, 0845, 0844, 1090);
  lut lut_gate382(0x1f, 1090, G7, 0755, 1091);
  lut lut_gate383(0x40, 0854, 0851, 0850, 1092);
  lut lut_gate384(0x4f, 1092, G43, 0755, 1093);
  lut lut_gate385(0x8, 1093, 1091, 1094);
  lut lut_gate386(0x10, 1102, 0859, G6, 1095);
  lut lut_gate387(0x3a, 0748, 1095, 0842, 1096);
  lut lut_gate388(0x87, 1096, 0818, 0748, 1097);
  lut lut_gate389(0xbc, 1097, 0818, 0823, G3533);
  lut lut_gate390(0x10, 1105, 0861, 0860, 1098);
  lut lut_gate391(0x4f, 1098, G22, 0755, 1099);
  lut lut_gate392(0x40, 0871, 0868, 0866, 1100);
  lut lut_gate393(0x4f, 1100, G42, 0755, 1101);
  lut lut_gate394(0x8, 1101, 1099, 1102);
  lut lut_gate395(0xf8, 0752, G7, G11, 1103);
  lut lut_gate396(0x40, 0862, 1103, G4, 1105);
  lut lut_gate397(0x10, 1139, 0912, G6, 1106);
  lut lut_gate398(0x3a, 0748, 1106, 0876, 1107);
  lut lut_gate399(0x4b, 1107, 0748, 0904, 1108);
  lut lut_gate400(0xe3, 1108, 0904, 0823, G3534);
  lut lut_gate401(0xa3, 1116, 0883, 0884, 1109);
  lut lut_gate402(0x35, 0800, G38, G32, 1110);
  lut lut_gate403(0xac, 0701, 1110, 0736, 1111);
  lut lut_gate404(0x4, G30, G49, 1112);
  lut lut_gate405(0x4, G3, 0792, 1114);
  lut lut_gate406(0x53, G9, 1114, 0796, 1115);
  lut lut_gate407(0x4, 1115, 1118, 1116);
  lut lut_gate408(0xca, G4, G10, G7, 1117);
  lut lut_gate409(0x10, 1117, 1063, G3, 1118);
  lut lut_gate410(0xc5, 1125, 0897, 0894, 1119);
  lut lut_gate411(0x4, G22, G4, 1120);
  lut lut_gate412(0xc5, G3, G8, 1120, 1121);
  lut lut_gate413(0x1e, 1121, G9, G3, 1122);
  lut lut_gate414(0xe3, 1122, G9, 0750, 1123);
  lut lut_gate415(0x35, G8, 0796, 1104, 1124);
  lut lut_gate416(0xb0, 1124, 1123, 1063, 1125);
  lut lut_gate417(0x35, G4, G30, G11, 1126);
  lut lut_gate418(0xef, 1126, 0896, 0895, 1127);
  lut lut_gate419(0x0b, 0802, 1127, 0736, 1128);
  lut lut_gate420(0xc5, G4, G8, G21, 1129);
  lut lut_gate421(0x35, 0800, G38, G30, 1131);
  lut lut_gate422(0x35, 1131, 1136, 0800, 1132);
  lut lut_gate423(0xac, 1132, 1131, 0736, 1133);
  lut lut_gate424(0x4, G28, G49, 1134);
  lut lut_gate425(0xf4, 0776, G4, G29, 1135);
  lut lut_gate426(0x0, 1135, G4, 1134, 1136);
  lut lut_gate427(0xf8, 0882, 1109, 0795, 1137);
  lut lut_gate428(0x35, G4, 0841, 0917, 1138);
  lut lut_gate429(0x4f, 0713, 1138, 0764, 1139);
  lut lut_gate430(0x4f, G18, 1017, G26, 1140);
  lut lut_gate431(0x4f, G22, 1017, 0754, 1141);
  lut lut_gate432(0x80, 0914, 1141, 1140, 1142);
  lut lut_gate433(0x10, 1149, 0918, G6, 1143);
  lut lut_gate434(0x3a, 0748, 1143, 0726, 1144);
  lut lut_gate435(0x4b, 1144, 0748, 0877, 1145);
  lut lut_gate436(0xe3, 1145, 0877, 0823, G3536);
  lut lut_gate437(0x4, 0923, 0844, 1146);
  lut lut_gate438(0xca, G4, 1146, 0717, 1147);
  lut lut_gate439(0x35, G4, 0867, 0920, 1148);
  lut lut_gate440(0x4f, 1147, 1148, 0764, 1149);
  lut lut_gate441(0x1f, 0726, 0904, 0877, 1150);
  lut lut_gate442(0xf4, 0823, 1150, 0748, 1151);
  lut lut_gate443(0xf8, 1155, 1151, 0931, G3535);
  lut lut_gate444(0x10, G5, 0943, 0942, 1152);
  lut lut_gate445(0x1f, 0721, 0939, G2, 1153);
  lut lut_gate446(0x07, 1160, 1153, G4, 1154);
  lut lut_gate447(0x8, 0747, 1154, 1155);
  lut lut_gate448(0x8f, G16, 1017, G26, 1156);
  lut lut_gate449(0xf4, G13, 1017, G26, 1157);
  lut lut_gate450(0xf4, G9, 1017, 0754, 1158);
  lut lut_gate451(0x40, 0698, 0945, 0947, 1159);
  lut lut_gate452(0x80, 1159, 1158, 1157, 1160);
  lut lut_gate453(0x40, 0956, 0963, 0966, 1161);
  lut lut_gate454(0x4f, 1161, G34, G11, 1162);
  lut lut_gate455(0x4, 0744, 0971, 1163);
  lut lut_gate456(0x07, 0968, G34, 1163, 1164);
  lut lut_gate457(0xb0, 1164, 1162, 0967, G3521);
  lut lut_gate458(0xc5, 0745, 1167, 0724, 1165);
  lut lut_gate459(0xb, 1165, 0998, G3530);
  lut lut_gate460(0x6f, 0987, G8, G9, 1166);
  lut lut_gate461(0xb0, 1166, G7, G9, 1167);
  lut lut_gate462(0xf4, G12, 1017, 0754, 1168);
  lut lut_gate463(0xf4, G8, 1017, G26, 1169);
  lut lut_gate464(0x10, 0760, 0757, 0751, 1170);
  lut lut_gate465(0x80, 1170, 1169, 1168, 1171);
  lut lut_gate466(0xf8, 0775, 1027, 1026, 1172);
  lut lut_gate467(0x0b, 0783, 1172, 0786, 1174);
  lut lut_gate468(0x2b, 1051, 1035, G24, 1175);
  lut lut_gate469(0xbc, 1175, G24, 0738, 1176);
  lut lut_gate470(0x4f, G40, 1017, G26, 1177);
  lut lut_gate471(0x8f, G19, 1017, G26, 1178);
  lut lut_gate472(0xf4, G8, 1017, 0754, 1179);
  lut lut_gate473(0xf4, 0752, G9, G21, 0686);
  lut lut_gate474(0x40, 1179, 1178, 0812, 0687);
  lut lut_gate475(0x40, 0686, 0687, 0814, 0688);
  lut lut_gate476(0xca, G4, 0730, 0688, 0689);
  lut lut_gate477(0xa3, 0743, 1013, 1054, 0690);
  lut lut_gate478(0x96, 1048, 0817, 0690, 0691);
  lut lut_gate479(0x8f, G20, 1017, G26, 0692);
  lut lut_gate480(0xf4, G9, 1017, 0754, 0693);
  lut lut_gate481(0x10, 0830, 0834, 0829, 0695);
  lut lut_gate482(0x80, 0695, 0693, 0692, 0696);
  lut lut_gate483(0xf8, 0752, G12, G8, 0697);
  lut lut_gate484(0x10, 0697, 0849, G4, 0698);
  lut lut_gate485(0x1, 1112, G12, 0699);
  lut lut_gate486(0xc5, G4, G31, 0699, 0700);
  lut lut_gate487(0xc5, 1110, 0700, 0800, 0701);
  lut lut_gate488(0xac, 1063, G3, 0797, 0702);
  lut lut_gate489(0xc5, G7, 0702, 1104, 0703);
  lut lut_gate490(0xb4, 0703, G7, 1063, 0704);
  lut lut_gate491(0xca, 0702, 0900, 1129, 0705);
  lut lut_gate492(0xe0, 0704, 1063, 0705, 0706);
  lut lut_gate493(0xf8, 0893, 1137, 1119, 0707);
  lut lut_gate494(0x0b, 0899, 0707, 0902, 0708);
  lut lut_gate495(0x01, 0913, 0861, 0751, 0709);
  lut lut_gate496(0x8, 0760, 0709, 0710);
  lut lut_gate497(0xca, G4, 0710, 1142, 0711);
  lut lut_gate498(0xca, G4, G39, G17, 0712);
  lut lut_gate499(0xb0, 0711, 0712, 0758, 0713);
  lut lut_gate500(0x4f, G19, 1017, G26, 0714);
  lut lut_gate501(0xf4, G7, 1017, 0754, 0715);
  lut lut_gate502(0x01, 0922, 0921, 0919, 0716);
  lut lut_gate503(0x80, 0716, 0715, 0714, 0717);
  lut lut_gate504(0x4f, G17, 1017, G26, 0718);
  lut lut_gate505(0x4f, G21, 1017, 0754, 0719);
  lut lut_gate506(0x40, 1156, 1152, 0941, 0720);
  lut lut_gate507(0x7f, 0720, 0719, 0718, 0721);
  lut lut_gate508(0x4b, 0890, 0934, 0794, 0722);
  lut lut_gate509(0x80, 1066, 0722, G47, 0723);
  lut lut_gate510(0x41, 0996, 0723, 0967, 0724);
  lut lut_gate511(0x07, 0890, 0772, 0708, 0725);
  lut lut_gate512(0x80, 1066, 0725, G47, 0726);
  lut lut_gate513(0xf4, G12, 1017, 0754, 0727);
  lut lut_gate514(0x8f, G41, 1017, G26, 0728);
  lut lut_gate515(0x10, 1177, 0810, 0808, 0729);
  lut lut_gate516(0x80, 0729, 0728, 0727, 0730);

endmodule
