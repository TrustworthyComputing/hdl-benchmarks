module c432(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G426, G427, G428, G429, G430, G431, G432, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, G203, G213, G308, G318, G358;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G5, G6, G7, G8, G9;
  output G426, G427, G428, G429, G430, G431, G432;
  lut lut_gate1(0xb, 196, 215, G427);
  lut lut_gate2(0x8000, 212, 209, 206, 197, 196);
  lut lut_gate3(0xb0bb, 198, G19, 205, G31, 197);
  lut lut_gate4(0x4f00, G18, G16, 199, 204, 198);
  lut lut_gate5(0x8000, 203, 202, 201, 200, 199);
  lut lut_gate6(0xb0bb, G14, G12, G26, G24, 200);
  lut lut_gate7(0xb0bb, G10, G8, G22, G20, 201);
  lut lut_gate8(0xb0bb, G2, G1, G6, G4, 202);
  lut lut_gate9(0xb0bb, G18, G16, G30, G28, 203);
  lut lut_gate10(0x4, G34, G32, 204);
  lut lut_gate11(0x4f00, G30, G28, 199, 204, 205);
  lut lut_gate12(0xb0bb, 207, G15, 208, G11, 206);
  lut lut_gate13(0x4f00, G14, G12, 199, 204, 207);
  lut lut_gate14(0x4f00, G10, G8, 199, 204, 208);
  lut lut_gate15(0xb0bb, 210, G23, 211, G7, 209);
  lut lut_gate16(0x4f00, G22, G20, 199, 204, 210);
  lut lut_gate17(0x4f00, G6, G4, 199, 204, 211);
  lut lut_gate18(0xb0bb, 213, G3, 214, G27, 212);
  lut lut_gate19(0x4f00, G2, G1, 199, 204, 213);
  lut lut_gate20(0x4f00, G26, G24, 199, 204, 214);
  lut lut_gate21(0x4, 216, G35, 215);
  lut lut_gate22(0x0, G34, 199, G32, 216);
  lut lut_gate23(0x7, 223, 217, G428);
  lut lut_gate24(0x0001, 221, 220, 219, 218, 217);
  lut lut_gate25(0x0700, 205, G33, G427, G31, 218);
  lut lut_gate26(0x0700, 198, G21, G427, G19, 219);
  lut lut_gate27(0x0700, 213, G5, G427, G3, 220);
  lut lut_gate28(0x1, G36, 222, 221);
  lut lut_gate29(0x4f, 216, G35, 196, 222);
  lut lut_gate30(0x0100, 227, 226, 225, 224, 223);
  lut lut_gate31(0x0700, 207, G17, G427, G15, 224);
  lut lut_gate32(0x0700, 208, G13, G427, G11, 225);
  lut lut_gate33(0x0700, 211, G9, G427, G7, 226);
  lut lut_gate34(0xb0bb, 228, G29, 229, G25, 227);
  lut lut_gate35(0x4f00, 214, G27, 196, 215, 228);
  lut lut_gate36(0x4f00, 210, G23, 196, 215, 229);
  lut lut_gate37(0xb, 199, 204, G426);
  lut lut_gate38(0x00bf, 244, 238, 240, G430, G429);
  lut lut_gate39(0xfeff, 232, 236, 234, 230, G430);
  lut lut_gate40(0x8f00, 231, G17, 217, 223, 230);
  lut lut_gate41(0x70, 207, G427, G15, 231);
  lut lut_gate42(0x70ff, 233, G21, 217, 223, 232);
  lut lut_gate43(0x70, 198, G427, G19, 233);
  lut lut_gate44(0x8f00, 235, G13, 217, 223, 234);
  lut lut_gate45(0x70, 208, G427, G11, 235);
  lut lut_gate46(0x8f00, 237, G9, 217, 223, 236);
  lut lut_gate47(0x70, 211, G427, G7, 237);
  lut lut_gate48(0x4, 222, 239, 238);
  lut lut_gate49(0x8f00, 229, G25, 217, 223, 239);
  lut lut_gate50(0x1, 243, 241, 240);
  lut lut_gate51(0xb0, 242, G33, 217, 241);
  lut lut_gate52(0x70, 205, G427, G31, 242);
  lut lut_gate53(0xb0, 228, G29, 217, 243);
  lut lut_gate54(0x70, 245, G428, G5, 244);
  lut lut_gate55(0x70, 213, G427, G3, 245);
  lut lut_gate56(0xf2ff, 194, 193, G430, 243, G431);
  lut lut_gate57(0x1000, 239, 232, 234, 230, 193);
  lut lut_gate58(0x1, 236, 234, 194);
  lut lut_gate59(0xfe, 236, 195, 193, G432);
  lut lut_gate60(0x00f4, 234, 230, 241, 243, 195);

endmodule
