module c5315(G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G16, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G17, G170, G171, G172, G173, G174, G175, G176, G177, G178, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G5193, G5194, G5195, G5196, G5197, G5198, G5199, G52, G5200, G5201, G5202, G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212, G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222, G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232, G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242, G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252, G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262, G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272, G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282, G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292, G5293, G5294, G5295, G5296, G5297, G5298, G5299, G53, G5300, G5301, G5302, G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312, G5313, G5314, G5315, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, 0950, 0951, 0952, 0953, 0954, 0955, 0956, 0957, 0958, 0959, 0960, 0961, 0962, 0963, 0964, 0965, 0966, 0967, 0968, 0969, 0970, 0971, 0972, 0973, 0974, 0975, 0976, 0977, 0978, 0979, 0980, 0981, 0982, 0983, 0984, 0985, 0986, 0987, 0988, 0989, 0990, 0991, 0992, 0993, 0994, 0995, 0996, 0997, 0998, 0999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165, 1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187, 1188, 1189, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198, 1199, 1200, 1201, 1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209, 1210, 1211, 1212, 1213, 1214, 1215, 1216, 1217, 1218, 1219, 1220, 1221, 1222, 1223, 1224, 1225, 1226, 1227, 1228, 1229, 1230, 1231, 1232, 1233, 1234, 1235, 1236, 1237, 1238, 1239, 1240, 1241, 1242, 1243, 1244, 1245, 1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264, 1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 1274, 1275, 1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 1286, 1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297, 1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308, 1309, 1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319, 1320, 1321, 1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361, 1362, 1363, 1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371, 1372, 1373, 1374, 1375, 1376, 1377, 1378, 1379, 1380, 1381, 1382, 1383, 1384, 1385, 1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 1394, 1395, 1396, 1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 1418, 1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429, 1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440, 1441, 1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451, 1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495, 1496, 1497, 1498, 1499, 1500, 1501, 1502, 1503, 1504, 1505, 1506, 1507, 1508, 1509, 1510, 1511, 1512, 1513, 1514, 1515, 1516, 1517, 1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550, 1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561, 1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572, 1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1601, 1602, 1603, 1604, 1605, 1606, 1607, 1608, 1609, 1610, 1611, 1612, 1613, 1614, 1615, 1616, 1617, 1618, 1619, 1620, 1621, 1622, 1623, 1624, 1625, 1626, 1627, 1628, 1629, 1630, 1631, 1632, 1633, 1634, 1635, 1636, 1637, 1638, 1639, 1640, 1641, 1642, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1651, 1652, 1653, 1654, 1655, 1656, 1657, 1658, 1659, 1660, 1661, 1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 1670, 1671, 1672, 1673, 1674, 1675, 1676, G1099, G1425, G1501, G1502, G1503, G1504, G1505, G1506, G1507, G1508, G1509, G1510, G1511, G1512, G1513, G1514, G1515, G1516, G1517, G1518, G1519, G1520, G1526, G1537, G1548, G1554, G1565, G1577, G1582, G1583, G1584, G1585, G1586, G1587, G1588, G1589, G1590, G1591, G1592, G1593, G1594, G1595, G1601, G1612, G1623, G1629, G1640, G1652, G1663, G1674, G1685, G1696, G1697, G1698, G1699, G1700, G1701, G1702, G1703, G1712, G1713, G1714, G1715, G1716, G1717, G1718, G1719, G1728, G1734, G1750, G1755, G1764, G1774, G1775, G1776, G1777, G1778, G1779, G1786, G1787, G1788, G1789, G1790, G1791, G1799, G1800, G1801, G1802, G1803, G1804, G1805, G1806, G1815, G1821, G1837, G1846, G1847, G1848, G1849, G1850, G1851, G1860, G1861, G1862, G1863, G1864, G1865, G1872, G1873, G1876, G1879, G1880, G1883, G1888, G1889, G1890, G1891, G1892, G1893, G1894, G1895, G1904, G1905, G1906, G1907, G1908, G1911, G1914, G1925, G1936, G1941, G1948, G1959, G1970, G1981, G1992, G2003, G2014, G2015, G2016, G2017, G2018, G2019, G2020, G2031, G2042, G2053, G2064, G2067, G2068, G2069, G2070, G2071, G2072, G2073, G2076, G3688, G4264, G4377, G4716, G4776, G4777, G685, G993;
  input G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G16, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G17, G170, G171, G172, G173, G174, G175, G176, G177, G178, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202, G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212, G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222, G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232, G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242, G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252, G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262, G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272, G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282, G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292, G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302, G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312, G5313, G5314, G5315;
  lut lut_gate1(0x9, 1250, 1249, G5251);
  lut lut_gate2(0xca, G123, G115, G116, 1249);
  lut lut_gate3(0x53, G123, G114, G113, 1250);
  lut lut_gate4(0xb, G11, G164, G5212);
  lut lut_gate5(0x7, G136, G154, G5213);
  lut lut_gate6(0xb, G65, G5221, G5220);
  lut lut_gate7(0x7, G12, G11, G5221);
  lut lut_gate8(0xe, 1251, G5221, G5228);
  lut lut_gate9(0x53, G163, G33, G34, 1251);
  lut lut_gate10(0xe, 1252, G5221, G5229);
  lut lut_gate11(0x35, G163, G13, G35, 1252);
  lut lut_gate12(0xb, G32, G5221, G5231);
  lut lut_gate13(0x07, 1253, 1258, G60, G5248);
  lut lut_gate14(0xe0, 1256, 1254, G176, 1253);
  lut lut_gate15(0x6, G21, 1255, 1254);
  lut lut_gate16(0x35, G123, G130, G131, 1255);
  lut lut_gate17(0x70, G177, 1257, G176, 1256);
  lut lut_gate18(0x35, G130, G101, G100, 1257);
  lut lut_gate19(0x4, G176, G177, 1258);
  lut lut_gate20(0x07, 1259, 1258, G58, G5249);
  lut lut_gate21(0xb0, 1263, 1260, G176, 1259);
  lut lut_gate22(0x6, 1255, 1261, 1260);
  lut lut_gate23(0x9, G150, 1262, 1261);
  lut lut_gate24(0x35, G123, G128, G129, 1262);
  lut lut_gate25(0x0, G177, 1264, G176, 1263);
  lut lut_gate26(0xca, G150, 1265, 1266, 1264);
  lut lut_gate27(0xca, G128, G168, G169, 1265);
  lut lut_gate28(0x35, G128, G167, G166, 1266);
  lut lut_gate29(0x07, 1267, 1258, G48, G5250);
  lut lut_gate30(0xe0, 1271, 1268, G176, 1267);
  lut lut_gate31(0x6, G2, 1269, 1268);
  lut lut_gate32(0x9, G135, 1270, 1269);
  lut lut_gate33(0x35, G124, G109, G110, 1270);
  lut lut_gate34(0x0, G177, 1272, G176, 1271);
  lut lut_gate35(0xca, G135, 1273, 1274, 1272);
  lut lut_gate36(0xac, G109, G169, G168, 1273);
  lut lut_gate37(0x53, G109, G166, G167, 1274);
  lut lut_gate38(0x0, 1287, 1275, G177, G5253);
  lut lut_gate39(0x53, G176, 1276, 1284, 1275);
  lut lut_gate40(0x6, 1282, 1277, 1276);
  lut lut_gate41(0xb2, 1281, G148, 1278, 1277);
  lut lut_gate42(0xb2, 1280, G149, 1279, 1278);
  lut lut_gate43(0x71, 1262, G150, 1255, 1279);
  lut lut_gate44(0x35, G123, G126, G127, 1280);
  lut lut_gate45(0x1, G125, G123, 1281);
  lut lut_gate46(0x6, G147, 1283, 1282);
  lut lut_gate47(0xca, G123, G121, G122, 1283);
  lut lut_gate48(0xca, G147, 1285, 1286, 1284);
  lut lut_gate49(0xca, G121, G168, G169, 1285);
  lut lut_gate50(0x35, G121, G167, G166, 1286);
  lut lut_gate51(0x8, G19, 1258, 1287);
  lut lut_gate52(0x07, 1288, 1258, G59, G5254);
  lut lut_gate53(0xb0, 1290, 1289, G176, 1288);
  lut lut_gate54(0x96, G148, 1281, 1278, 1289);
  lut lut_gate55(0x70, G177, 1291, G176, 1290);
  lut lut_gate56(0x3a, G148, G169, G166, 1291);
  lut lut_gate57(0x07, 1292, 1258, G50, G5255);
  lut lut_gate58(0xe0, 1295, 1293, G176, 1292);
  lut lut_gate59(0x6, 1294, 1279, 1293);
  lut lut_gate60(0x9, G149, 1280, 1294);
  lut lut_gate61(0x0, G177, 1296, G176, 1295);
  lut lut_gate62(0xca, G149, 1297, 1298, 1296);
  lut lut_gate63(0xca, G126, G168, G169, 1297);
  lut lut_gate64(0x35, G126, G167, G166, 1298);
  lut lut_gate65(0x0, 1319, 1299, 1315, G5257);
  lut lut_gate66(0x14, 1313, 1300, G176, 1299);
  lut lut_gate67(0x71, G137, 1312, 1301, 1300);
  lut lut_gate68(0x70, 1302, 1311, G2, 1301);
  lut lut_gate69(0x4, 1309, 1303, 1302);
  lut lut_gate70(0x80, 1307, 1305, 1304, 1303);
  lut lut_gate71(0x4, G135, 1270, 1304);
  lut lut_gate72(0x9, G138, 1306, 1305);
  lut lut_gate73(0x35, G124, G105, G106, 1306);
  lut lut_gate74(0x9, G139, 1308, 1307);
  lut lut_gate75(0x35, G124, G107, G108, 1308);
  lut lut_gate76(0x71, 1306, G138, 1310, 1309);
  lut lut_gate77(0x4, G139, 1308, 1310);
  lut lut_gate78(0x80, 1307, 1305, 1269, 1311);
  lut lut_gate79(0x35, G124, G103, G104, 1312);
  lut lut_gate80(0x9, G141, 1314, 1313);
  lut lut_gate81(0x35, G124, G96, G97, 1314);
  lut lut_gate82(0x0, G177, 1316, G176, 1315);
  lut lut_gate83(0xca, G141, 1317, 1318, 1316);
  lut lut_gate84(0xac, G96, G169, G168, 1317);
  lut lut_gate85(0x53, G96, G166, G167, 1318);
  lut lut_gate86(0x8, G53, 1258, 1319);
  lut lut_gate87(0x07, 1320, 1258, G57, G5258);
  lut lut_gate88(0xe0, 1323, 1321, G176, 1320);
  lut lut_gate89(0x6, 1322, 1301, 1321);
  lut lut_gate90(0x9, G137, 1312, 1322);
  lut lut_gate91(0x0, G177, 1324, G176, 1323);
  lut lut_gate92(0xca, G137, 1325, 1326, 1324);
  lut lut_gate93(0xac, G103, G169, G168, 1325);
  lut lut_gate94(0x53, G103, G166, G167, 1326);
  lut lut_gate95(0x07, 1327, 1258, G56, G5259);
  lut lut_gate96(0xb0, 1331, 1328, G176, 1327);
  lut lut_gate97(0x1e, 1305, 1310, 1329, 1328);
  lut lut_gate98(0xe0, 1307, 1330, 1304, 1329);
  lut lut_gate99(0x8, G2, 1269, 1330);
  lut lut_gate100(0x0, G177, 1332, G176, 1331);
  lut lut_gate101(0xca, G138, 1333, 1334, 1332);
  lut lut_gate102(0xac, G105, G169, G168, 1333);
  lut lut_gate103(0x53, G105, G166, G167, 1334);
  lut lut_gate104(0x07, 1335, 1258, G55, G5260);
  lut lut_gate105(0xb0, 1337, 1336, G176, 1335);
  lut lut_gate106(0x1e, 1307, 1304, 1330, 1336);
  lut lut_gate107(0x0, G177, 1338, G176, 1337);
  lut lut_gate108(0xca, G139, 1339, 1340, 1338);
  lut lut_gate109(0xac, G107, G169, G168, 1339);
  lut lut_gate110(0x53, G107, G166, G167, 1340);
  lut lut_gate111(0x07, 1341, 1258, G54, G5285);
  lut lut_gate112(0xb0, 1342, G5251, G176, 1341);
  lut lut_gate113(0x70, G177, 1343, G176, 1342);
  lut lut_gate114(0x35, G113, G102, G98, 1343);
  lut lut_gate115(0x0, 1354, 1344, 1355, G5286);
  lut lut_gate116(0x14, 1249, 1345, G176, 1344);
  lut lut_gate117(0x70, 1347, 1346, 1351, 1345);
  lut lut_gate118(0x4, G147, 1283, 1277, 1346);
  lut lut_gate119(0x71, 1350, G145, 1348, 1347);
  lut lut_gate120(0x4, G146, 1349, 1348);
  lut lut_gate121(0x35, G123, G119, G120, 1349);
  lut lut_gate122(0x35, G123, G117, G118, 1350);
  lut lut_gate123(0x8, 1353, 1352, 1351);
  lut lut_gate124(0x9, G145, 1350, 1352);
  lut lut_gate125(0x9, G146, 1349, 1353);
  lut lut_gate126(0x8, G52, 1258, 1354);
  lut lut_gate127(0x70, G177, 1356, G176, 1355);
  lut lut_gate128(0x35, G115, G101, G100, 1356);
  lut lut_gate129(0x07, 1357, 1258, G47, G5287);
  lut lut_gate130(0xb0, 1360, 1358, G176, 1357);
  lut lut_gate131(0x9, 1352, 1359, 1358);
  lut lut_gate132(0x18, G146, 1349, 1346, 1359);
  lut lut_gate133(0x0, G177, 1361, G176, 1360);
  lut lut_gate134(0xca, G145, 1362, 1363, 1361);
  lut lut_gate135(0xca, G117, G101, G100, 1362);
  lut lut_gate136(0x35, G117, G102, G98, 1363);
  lut lut_gate137(0x07, 1364, 1258, G43, G5288);
  lut lut_gate138(0xe0, 1366, 1365, G176, 1364);
  lut lut_gate139(0x6, 1353, 1346, 1365);
  lut lut_gate140(0x0, G177, 1367, G176, 1366);
  lut lut_gate141(0xca, G146, 1368, 1369, 1367);
  lut lut_gate142(0xca, G119, G101, G100, 1368);
  lut lut_gate143(0x35, G119, G102, G98, 1369);
  lut lut_gate144(0x07, 1370, 1258, G46, G5290);
  lut lut_gate145(0xb0, 1398, 1371, G176, 1370);
  lut lut_gate146(0x9, 1396, 1372, 1371);
  lut lut_gate147(0x0, 1385, 1373, 1391, 1372);
  lut lut_gate148(0x70, 1374, 1383, G2, 1373);
  lut lut_gate149(0x01, 1382, 1378, 1375, 1374);
  lut lut_gate150(0x8, 1377, 1376, 1375);
  lut lut_gate151(0x8, 1307, 1304, 1376);
  lut lut_gate152(0x80, 1322, 1305, 1313, 1377);
  lut lut_gate153(0xb0, 1379, 1309, 1381, 1378);
  lut lut_gate154(0x4, 1313, 1380, 1379);
  lut lut_gate155(0x4, 1312, G137, 1380);
  lut lut_gate156(0x4, G137, 1312, 1381);
  lut lut_gate157(0x4, G141, 1314, 1382);
  lut lut_gate158(0x8, 1313, 1384, 1383);
  lut lut_gate159(0x8, 1322, 1311, 1384);
  lut lut_gate160(0xb2, 1390, G143, 1386, 1385);
  lut lut_gate161(0x71, 1389, G144, 1387, 1386);
  lut lut_gate162(0x4, G140, 1388, 1387);
  lut lut_gate163(0x35, G124, G94, G95, 1388);
  lut lut_gate164(0x35, G124, G92, G93, 1389);
  lut lut_gate165(0x35, G124, G90, G91, 1390);
  lut lut_gate166(0x8, 1395, 1392, 1391);
  lut lut_gate167(0x8, 1394, 1393, 1392);
  lut lut_gate168(0x9, G144, 1389, 1393);
  lut lut_gate169(0x9, G140, 1388, 1394);
  lut lut_gate170(0x9, G143, 1390, 1395);
  lut lut_gate171(0x9, G142, 1397, 1396);
  lut lut_gate172(0x35, G124, G88, G89, 1397);
  lut lut_gate173(0x0, G177, 1399, G176, 1398);
  lut lut_gate174(0xca, G142, 1400, 1401, 1399);
  lut lut_gate175(0xca, G88, G100, G101, 1400);
  lut lut_gate176(0x35, G88, G98, G102, 1401);
  lut lut_gate177(0x0, 1408, 1402, 1404, G5291);
  lut lut_gate178(0x41, 1403, 1395, G176, 1402);
  lut lut_gate179(0x0, 1386, 1373, 1392, 1403);
  lut lut_gate180(0x0, G177, 1405, G176, 1404);
  lut lut_gate181(0xca, G143, 1406, 1407, 1405);
  lut lut_gate182(0xac, G90, G169, G168, 1406);
  lut lut_gate183(0x53, G90, G166, G167, 1407);
  lut lut_gate184(0x8, G45, 1258, 1408);
  lut lut_gate185(0x0, 1415, 1409, 1411, G5292);
  lut lut_gate186(0x14, 1393, 1410, G176, 1409);
  lut lut_gate187(0xe7, 1388, G140, 1373, 1410);
  lut lut_gate188(0x0, G177, 1412, G176, 1411);
  lut lut_gate189(0xca, G144, 1413, 1414, 1412);
  lut lut_gate190(0xac, G92, G169, G168, 1413);
  lut lut_gate191(0x53, G92, G166, G167, 1414);
  lut lut_gate192(0x8, G20, 1258, 1415);
  lut lut_gate193(0x0, 1421, 1416, G177, G5293);
  lut lut_gate194(0x5c, G176, 1417, 1418, 1416);
  lut lut_gate195(0x6, 1394, 1373, 1417);
  lut lut_gate196(0xca, G140, 1419, 1420, 1418);
  lut lut_gate197(0xac, G94, G169, G168, 1419);
  lut lut_gate198(0x53, G94, G166, G167, 1420);
  lut lut_gate199(0x8, G44, 1258, 1421);
  lut lut_gate200(0x0e, 1244, G177, G38, 1422);
  lut lut_gate201(0x53, 1394, 1424, 1427, 1423);
  lut lut_gate202(0xb4, 1425, 1385, 1391, 1424);
  lut lut_gate203(0x18, 1389, G144, 1426, 1425);
  lut lut_gate204(0x4, 1388, G140, 1426);
  lut lut_gate205(0x18, 1390, G143, 1386, 1427);
  lut lut_gate206(0x69, 1393, 1395, 1396, 1428);
  lut lut_gate207(0x96, 1394, 1428, 1424, 1429);
  lut lut_gate208(0x69, 1434, 1433, 1431, 1430);
  lut lut_gate209(0x0e, 1384, 1432, 1380, 1431);
  lut lut_gate210(0x10, 1309, 1381, 1303, 1432);
  lut lut_gate211(0x6, 1307, 1269, 1433);
  lut lut_gate212(0x6, 1305, 1313, 1434);
  lut lut_gate213(0xe7, 1308, G139, 1436, 1435);
  lut lut_gate214(0x4, 1270, G135, 1436);
  lut lut_gate215(0xe1, 1438, 1380, 1432, 1437);
  lut lut_gate216(0x1e, 1433, 1310, 1376, 1438);
  lut lut_gate217(0xbc, 1304, 1309, 1303, 1439);
  lut lut_gate218(0x69, 1448, 1445, 1441, 1440);
  lut lut_gate219(0x6, 1442, 1399, 1441);
  lut lut_gate220(0xca, G143, 1443, 1444, 1442);
  lut lut_gate221(0xac, G90, G100, G101, 1443);
  lut lut_gate222(0x53, G90, G98, G102, 1444);
  lut lut_gate223(0xca, G140, 1446, 1447, 1445);
  lut lut_gate224(0xac, G94, G100, G101, 1446);
  lut lut_gate225(0x53, G94, G98, G102, 1447);
  lut lut_gate226(0xca, G144, 1449, 1450, 1448);
  lut lut_gate227(0xac, G92, G100, G101, 1449);
  lut lut_gate228(0x53, G92, G98, G102, 1450);
  lut lut_gate229(0x96, 1465, 1462, 1452, 1451);
  lut lut_gate230(0x96, 1459, 1456, 1453, 1452);
  lut lut_gate231(0xca, G141, 1454, 1455, 1453);
  lut lut_gate232(0xac, G96, G100, G101, 1454);
  lut lut_gate233(0x35, G96, G102, G98, 1455);
  lut lut_gate234(0xca, G135, 1457, 1458, 1456);
  lut lut_gate235(0xac, G109, G100, G101, 1457);
  lut lut_gate236(0x35, G109, G102, G98, 1458);
  lut lut_gate237(0xca, G137, 1460, 1461, 1459);
  lut lut_gate238(0xac, G103, G100, G101, 1460);
  lut lut_gate239(0x35, G103, G102, G98, 1461);
  lut lut_gate240(0xca, G138, 1463, 1464, 1462);
  lut lut_gate241(0xac, G105, G100, G101, 1463);
  lut lut_gate242(0x35, G105, G102, G98, 1464);
  lut lut_gate243(0xca, G139, 1466, 1467, 1465);
  lut lut_gate244(0xac, G107, G100, G101, 1466);
  lut lut_gate245(0x35, G107, G102, G98, 1467);
  lut lut_gate246(0x0e, 1606, G177, G37, 1468);
  lut lut_gate247(0x18, 1350, G145, 1470, 1469);
  lut lut_gate248(0x4, 1349, G146, 1470);
  lut lut_gate249(0x69, G5251, 1277, 1472, 1471);
  lut lut_gate250(0x96, 1476, 1278, 1473, 1472);
  lut lut_gate251(0x69, 1294, 1475, 1474, 1473);
  lut lut_gate252(0x69, G148, 1281, 1282, 1474);
  lut lut_gate253(0x1e, 1261, G162, 1255, 1475);
  lut lut_gate254(0x18, G150, 1262, 1255, 1476);
  lut lut_gate255(0x90, G176, 1490, 1478, 1477);
  lut lut_gate256(0x69, 1487, 1484, 1479, 1478);
  lut lut_gate257(0x96, 1483, 1257, 1480, 1479);
  lut lut_gate258(0xca, G150, 1481, 1482, 1480);
  lut lut_gate259(0xca, G128, G101, G100, 1481);
  lut lut_gate260(0x35, G128, G102, G98, 1482);
  lut lut_gate261(0x3a, G148, G100, G98, 1483);
  lut lut_gate262(0xca, G147, 1485, 1486, 1484);
  lut lut_gate263(0xca, G121, G101, G100, 1485);
  lut lut_gate264(0x35, G121, G102, G98, 1486);
  lut lut_gate265(0xca, G149, 1488, 1489, 1487);
  lut lut_gate266(0xca, G126, G101, G100, 1488);
  lut lut_gate267(0x35, G126, G102, G98, 1489);
  lut lut_gate268(0x96, 1491, 1367, 1361, 1490);
  lut lut_gate269(0x9, 1356, 1343, 1491);
  lut lut_gate270(0x8, G134, G1, G5210);
  lut lut_gate271(0x6, 1494, 1492, G5242);
  lut lut_gate272(0x69, G115, G119, 1493, 1492);
  lut lut_gate273(0x9, G117, G113, 1493);
  lut lut_gate274(0x96, G128, G126, 1495, 1494);
  lut lut_gate275(0x69, G132, G130, G121, 1495);
  lut lut_gate276(0x6, 1499, 1496, G5243);
  lut lut_gate277(0x96, G90, G88, 1497, 1496);
  lut lut_gate278(0x69, G107, G105, 1498, 1497);
  lut lut_gate279(0x6, G94, G92, 1498);
  lut lut_gate280(0x69, G111, G103, 1500, 1499);
  lut lut_gate281(0x9, G96, G109, 1500);
  lut lut_gate282(0x69, 1504, G5251, 1501, G5261);
  lut lut_gate283(0x69, 1255, 1503, 1502, 1501);
  lut lut_gate284(0x9, 1281, 1283, 1502);
  lut lut_gate285(0x6, 1349, 1350, 1503);
  lut lut_gate286(0x69, 1505, 1280, 1262, 1504);
  lut lut_gate287(0x35, G123, G132, G133, 1505);
  lut lut_gate288(0x9, 1508, 1506, G5262);
  lut lut_gate289(0x96, 1308, 1306, 1507, 1506);
  lut lut_gate290(0x9, 1312, 1270, 1507);
  lut lut_gate291(0x69, 1388, 1510, 1509, 1508);
  lut lut_gate292(0x6, 1389, 1390, 1509);
  lut lut_gate293(0x96, 1511, 1397, 1314, 1510);
  lut lut_gate294(0x35, G124, G111, G112, 1511);
  lut lut_gate295(0x8, G156, G153, G5199);
  lut lut_gate296(0x8, G67, G66, G5205);
  lut lut_gate297(0x4, G63, G165, G5211);
  lut lut_gate298(0x8, 1515, 1512, G5236);
  lut lut_gate299(0x40, 1514, 1513, 1264, 1512);
  lut lut_gate300(0x40, 1291, 1257, 1296, 1513);
  lut lut_gate301(0x4, 1356, 1343, 1514);
  lut lut_gate302(0x01, 1367, 1361, 1284, 1515);
  lut lut_gate303(0x80, 1519, 1518, 1516, G5237);
  lut lut_gate304(0x10, 1517, 1332, 1324, 1516);
  lut lut_gate305(0x1, 1399, 1338, 1517);
  lut lut_gate306(0x01, 1418, 1412, 1405, 1518);
  lut lut_gate307(0x1, 1316, 1272, 1519);
  lut lut_gate308(0x80, 1396, 1391, 1383, G5238);
  lut lut_gate309(0x80, 1523, 1522, 1520, G5239);
  lut lut_gate310(0x8, 1521, 1351, 1520);
  lut lut_gate311(0x90, 1282, G148, 1281, 1521);
  lut lut_gate312(0x8, 1255, 1261, 1522);
  lut lut_gate313(0x40, 1250, 1294, 1249, 1523);
  lut lut_gate314(0x7, 1250, 1249, G5245);
  lut lut_gate315(0x8f, 1524, G22, 1528, G5252);
  lut lut_gate316(0x07, 1525, 1527, G3, 1524);
  lut lut_gate317(0xb0, 1526, G5250, G173, 1525);
  lut lut_gate318(0x70, G172, G5248, G173, 1526);
  lut lut_gate319(0x4, G173, G172, 1527);
  lut lut_gate320(0x1, G173, G172, 1528);
  lut lut_gate321(0x8f, 1529, G3, 1533, G5256);
  lut lut_gate322(0x07, 1530, 1532, G22, 1529);
  lut lut_gate323(0xb0, 1531, G5250, G174, 1530);
  lut lut_gate324(0x70, G175, G5248, G174, 1531);
  lut lut_gate325(0x1, G174, G175, 1532);
  lut lut_gate326(0x4, G174, G175, 1533);
  lut lut_gate327(0x80, 1371, 1536, 1534, G5263);
  lut lut_gate328(0x41, 1395, 1403, 1535, 1534);
  lut lut_gate329(0x9, 1393, 1410, 1535);
  lut lut_gate330(0x80, 1539, 1417, 1537, 1536);
  lut lut_gate331(0x60, 1538, 1313, 1300, 1537);
  lut lut_gate332(0x4, 1336, 1321, 1538);
  lut lut_gate333(0x4, 1328, 1268, 1539);
  lut lut_gate334(0x8, 1358, 1540, G5264);
  lut lut_gate335(0x60, 1541, 1249, 1345, 1540);
  lut lut_gate336(0x10, 1542, 1276, 1365, 1541);
  lut lut_gate337(0x40, 1289, 1543, 1293, 1542);
  lut lut_gate338(0x40, 1260, G5251, 1254, 1543);
  lut lut_gate339(0x8f, 1544, G14, 1528, G5267);
  lut lut_gate340(0x07, 1545, 1527, G16, 1544);
  lut lut_gate341(0xb0, 1546, G5257, G173, 1545);
  lut lut_gate342(0x70, G172, G5253, G173, 1546);
  lut lut_gate343(0x8f, 1547, G26, 1527, G5269);
  lut lut_gate344(0x07, 1548, 1528, G5, 1547);
  lut lut_gate345(0xb0, 1549, G5259, G173, 1548);
  lut lut_gate346(0x70, G172, G5255, G173, 1549);
  lut lut_gate347(0x8f, 1550, G24, 1527, G5270);
  lut lut_gate348(0x07, 1551, 1528, G25, 1550);
  lut lut_gate349(0xb0, 1552, G5260, G173, 1551);
  lut lut_gate350(0x70, G172, G5249, G173, 1552);
  lut lut_gate351(0x8f, 1553, G14, 1532, G5271);
  lut lut_gate352(0x07, 1554, 1533, G16, 1553);
  lut lut_gate353(0x70, 1555, G5253, G174, 1554);
  lut lut_gate354(0xb0, G175, G5257, G174, 1555);
  lut lut_gate355(0x8f, 1556, G26, 1533, G5273);
  lut lut_gate356(0x07, 1557, 1532, G5, 1556);
  lut lut_gate357(0xb0, 1558, G5259, G174, 1557);
  lut lut_gate358(0x70, G175, G5255, G174, 1558);
  lut lut_gate359(0x8f, 1559, G24, 1533, G5274);
  lut lut_gate360(0x07, 1560, 1532, G25, 1559);
  lut lut_gate361(0xb0, 1561, G5260, G174, 1560);
  lut lut_gate362(0x70, G175, G5249, G174, 1561);
  lut lut_gate363(0x4, G64, 1562, G5281);
  lut lut_gate364(0xca, G161, 1563, 1564, 1562);
  lut lut_gate365(0xac, G160, G5259, G5255, 1563);
  lut lut_gate366(0x35, G160, G71, G70, 1564);
  lut lut_gate367(0x0, 1567, 1565, G171, G5283);
  lut lut_gate368(0x3a, G170, G5251, 1566, 1565);
  lut lut_gate369(0x9, G61, 1250, 1566);
  lut lut_gate370(0x0e, 1569, 1568, G171, 1567);
  lut lut_gate371(0xa3, G170, 1343, G54, 1568);
  lut lut_gate372(0x8, G62, G178, 1569);
  lut lut_gate373(0x9, 1566, G5251, G5284);
  lut lut_gate374(0x8, G5262, 1570, G5289);
  lut lut_gate375(0x80, 1571, G5261, G5243, 1570);
  lut lut_gate376(0x80, G5199, 1572, G5242, 1571);
  lut lut_gate377(0x40, G155, G99, G5213, 1572);
  lut lut_gate378(0x8f, 1573, G18, 1528, G5296);
  lut lut_gate379(0x07, 1574, 1527, G17, 1573);
  lut lut_gate380(0xb0, 1575, G5291, G173, 1574);
  lut lut_gate381(0x70, G172, G5286, G173, 1575);
  lut lut_gate382(0x8f, 1576, G40, 1528, G5297);
  lut lut_gate383(0x07, 1577, 1527, G39, 1576);
  lut lut_gate384(0x70, 1578, G5287, G173, 1577);
  lut lut_gate385(0xb0, G172, G5292, G173, 1578);
  lut lut_gate386(0x8f, 1579, G15, 1528, G5298);
  lut lut_gate387(0x07, 1580, 1527, G36, 1579);
  lut lut_gate388(0xb0, 1581, G5293, G173, 1580);
  lut lut_gate389(0x70, G172, G5288, G173, 1581);
  lut lut_gate390(0x8f, 1582, G17, 1533, G5299);
  lut lut_gate391(0x07, 1583, 1532, G18, 1582);
  lut lut_gate392(0xb0, 1584, G5291, G174, 1583);
  lut lut_gate393(0x70, G175, G5286, G174, 1584);
  lut lut_gate394(0x8f, 1585, G40, 1532, G5300);
  lut lut_gate395(0x07, 1586, 1533, G39, 1585);
  lut lut_gate396(0x70, 1587, G5287, G174, 1586);
  lut lut_gate397(0xb0, G175, G5292, G174, 1587);
  lut lut_gate398(0x8f, 1588, G15, 1532, G5301);
  lut lut_gate399(0x07, 1589, 1533, G36, 1588);
  lut lut_gate400(0xb0, 1590, G5293, G174, 1589);
  lut lut_gate401(0x70, G175, G5288, G174, 1590);
  lut lut_gate402(0x4, G64, 1591, G5308);
  lut lut_gate403(0xca, G161, 1592, 1593, 1591);
  lut lut_gate404(0xac, G160, G5291, G5286, 1592);
  lut lut_gate405(0x35, G160, G84, G74, 1593);
  lut lut_gate406(0xe, 1594, 1606, G5310);
  lut lut_gate407(0x0b, G177, G176, G51, 1594);
  lut lut_gate408(0xe, 1595, 1244, G5311);
  lut lut_gate409(0x0b, G177, G176, G49, 1595);
  lut lut_gate410(0x1, G165, G5195);
  lut lut_gate411(0x1, G66, G5193);
  lut lut_gate412(0x1, G113, G5194);
  lut lut_gate413(0x1, G151, G5196);
  lut lut_gate414(0x1, G127, G5197);
  lut lut_gate415(0x1, G131, G5198);
  lut lut_gate416(0x1, G152, G5200);
  lut lut_gate417(0x1, G125, G5203);
  lut lut_gate418(0x1, G129, G5204);
  lut lut_gate419(0x1, G99, G5206);
  lut lut_gate420(0x1, G153, G5207);
  lut lut_gate421(0x1, G156, G5208);
  lut lut_gate422(0x1, G155, G5209);
  lut lut_gate423(0x1, G1, G5222);
  lut lut_gate424(0x1, G114, G5226);
  lut lut_gate425(0xca, G158, 1468, 1422, 1596);
  lut lut_gate426(0xca, G158, G78, G79, 1597);
  lut lut_gate427(0x3, G64, G159, 1597, 1598);
  lut lut_gate428(0x7c, 1598, G159, 1596, G5314);
  lut lut_gate429(0x6, 1428, 1423, 1599);
  lut lut_gate430(0xb4, 1435, 1302, 1311, 1600);
  lut lut_gate431(0x6, 1430, 1600, 1601);
  lut lut_gate432(0x96, 1439, 1437, 1434, 1602);
  lut lut_gate433(0x2c, 1353, 1352, 1346, 1603);
  lut lut_gate434(0x96, 1471, 1469, 1603, 1604);
  lut lut_gate435(0xbe, 1604, 1249, G176, 1605);
  lut lut_gate436(0x40, G177, 1605, 1477, 1606);
  lut lut_gate437(0xca, G160, G78, G79, 1607);
  lut lut_gate438(0x3, G64, G161, 1607, 1608);
  lut lut_gate439(0xca, G160, 1468, 1422, 1609);
  lut lut_gate440(0x7c, G161, 1608, 1609, G5315);
  lut lut_gate441(0x35, G163, G8, G9, 1610);
  lut lut_gate442(0xb0, G66, 1610, G5221, G5232);
  lut lut_gate443(0x35, G163, G10, G30, 1611);
  lut lut_gate444(0xb0, G66, 1611, G5221, G5233);
  lut lut_gate445(0x35, G163, G28, G7, 1612);
  lut lut_gate446(0xb0, G66, 1612, G5221, G5234);
  lut lut_gate447(0x35, G163, G31, G29, 1613);
  lut lut_gate448(0xb0, G66, 1613, G5221, G5235);
  lut lut_gate449(0x0, 1385, 1374, 1391, 1614);
  lut lut_gate450(0x2b, 1397, 1614, G142, G5244);
  lut lut_gate451(0xca, G158, G5248, G5250, 1615);
  lut lut_gate452(0xca, G158, G80, G81, 1616);
  lut lut_gate453(0x3a, G159, 1615, 1616, 1617);
  lut lut_gate454(0x8, G64, 1617, G5265);
  lut lut_gate455(0xca, G160, G5248, G5250, 1618);
  lut lut_gate456(0xca, G160, G80, G81, 1619);
  lut lut_gate457(0x3a, G161, 1618, 1619, 1620);
  lut lut_gate458(0x8, 1620, G64, G5266);
  lut lut_gate459(0xca, G173, G27, G6, 1621);
  lut lut_gate460(0xca, G174, G27, G6, 1622);
  lut lut_gate461(0xca, G158, G5253, G5257, 1623);
  lut lut_gate462(0xca, G158, G86, G76, 1624);
  lut lut_gate463(0x3a, G159, 1623, 1624, 1625);
  lut lut_gate464(0x8, G64, 1625, G5275);
  lut lut_gate465(0xca, G158, G5249, G5260, 1626);
  lut lut_gate466(0xca, G158, G82, G72, 1627);
  lut lut_gate467(0x3a, G159, 1626, 1627, 1628);
  lut lut_gate468(0x8, G64, 1628, G5276);
  lut lut_gate469(0xca, G158, G5255, G5259, 1629);
  lut lut_gate470(0xca, G158, G71, G70, 1630);
  lut lut_gate471(0x3a, G159, 1629, 1630, 1631);
  lut lut_gate472(0x8, G64, 1631, G5277);
  lut lut_gate473(0xca, G158, G5254, G5258, 1632);
  lut lut_gate474(0xca, G158, G69, G68, 1633);
  lut lut_gate475(0x3a, G159, 1632, 1633, 1634);
  lut lut_gate476(0x8, G64, 1634, G5278);
  lut lut_gate477(0xca, G160, G5253, G5257, 1635);
  lut lut_gate478(0xca, G160, G86, G76, 1636);
  lut lut_gate479(0x3a, G161, 1635, 1636, 1637);
  lut lut_gate480(0x8, 1637, G64, G5279);
  lut lut_gate481(0xca, G160, G5249, G5260, 1638);
  lut lut_gate482(0xca, G160, G82, G72, 1639);
  lut lut_gate483(0x3a, G161, 1638, 1639, 1640);
  lut lut_gate484(0x8, 1640, G64, G5280);
  lut lut_gate485(0xca, G160, G5254, G5258, 1641);
  lut lut_gate486(0xca, G160, G69, G68, 1642);
  lut lut_gate487(0x3a, G161, 1641, 1642, 1643);
  lut lut_gate488(0x8, 1643, G64, G5282);
  lut lut_gate489(0x35, G174, G5285, G5290, 1644);
  lut lut_gate490(0x35, G173, G5285, G5290, 1645);
  lut lut_gate491(0xca, G158, G5288, G5293, 1646);
  lut lut_gate492(0xca, G158, G87, G77, 1647);
  lut lut_gate493(0x3a, G159, 1646, 1647, 1648);
  lut lut_gate494(0x8, G64, 1648, G5302);
  lut lut_gate495(0xca, G158, G5287, G5292, 1649);
  lut lut_gate496(0xca, G158, G85, G75, 1650);
  lut lut_gate497(0x3a, G159, 1649, 1650, 1651);
  lut lut_gate498(0x8, G64, 1651, G5303);
  lut lut_gate499(0xca, G158, G5286, G5291, 1652);
  lut lut_gate500(0xca, G158, G84, G74, 1653);
  lut lut_gate501(0x3a, G159, 1652, 1653, 1654);
  lut lut_gate502(0x8, G64, 1654, G5304);
  lut lut_gate503(0xca, G158, G5285, G5290, 1655);
  lut lut_gate504(0xca, G158, G83, G73, 1656);
  lut lut_gate505(0x3a, G159, 1655, 1656, 1657);
  lut lut_gate506(0x8, G64, 1657, G5305);
  lut lut_gate507(0xca, G160, G5288, G5293, 1658);
  lut lut_gate508(0xca, G160, G87, G77, 1659);
  lut lut_gate509(0x3a, G161, 1658, 1659, 1660);
  lut lut_gate510(0x8, 1660, G64, G5306);
  lut lut_gate511(0xca, G160, G5287, G5292, 1661);
  lut lut_gate512(0xca, G160, G85, G75, 1662);
  lut lut_gate513(0x3a, G161, 1661, 1662, 1663);
  lut lut_gate514(0x8, 1663, G64, G5307);
  lut lut_gate515(0xca, G160, G5285, G5290, 1664);
  lut lut_gate516(0xca, G160, G83, G73, 1665);
  lut lut_gate517(0x3a, G161, 1664, 1665, 1666);
  lut lut_gate518(0x8, 1666, G64, G5309);
  lut lut_gate519(0x6, G173, G172, 1667);
  lut lut_gate520(0xca, G172, 1422, G4, 1668);
  lut lut_gate521(0xca, G172, 1468, G23, 1669);
  lut lut_gate522(0xca, 1667, 1668, 1669, G5312);
  lut lut_gate523(0x6, G174, G175, 1670);
  lut lut_gate524(0xca, G175, 1422, G4, 1671);
  lut lut_gate525(0xca, G175, 1468, G23, 1672);
  lut lut_gate526(0xca, 1670, 1671, 1672, G5313);
  lut lut_gate527(0x70, 1374, G157, 1383, 1673);
  lut lut_gate528(0xc5, 1673, 1599, 1429, 1674);
  lut lut_gate529(0x6, 1451, 1440, 1675);
  lut lut_gate530(0x70, G177, G176, 1675, 1676);
  lut lut_gate531(0xc5, G157, 1601, 1602, 1242);
  lut lut_gate532(0x96, 1674, 1322, 1242, 1243);
  lut lut_gate533(0xe0, 1676, G176, 1243, 1244);
  lut lut_gate534(0xca, G173, G5254, G5258, 1245);
  lut lut_gate535(0x3a, G172, 1245, 1621, G5268);
  lut lut_gate536(0xca, G174, G5254, G5258, 1246);
  lut lut_gate537(0x3a, G175, 1246, 1622, G5272);
  lut lut_gate538(0xca, G174, G42, G41, 1247);
  lut lut_gate539(0xca, G175, 1644, 1247, G5294);
  lut lut_gate540(0xca, G173, G42, G41, 1248);
  lut lut_gate541(0xca, G172, 1645, 1248, G5295);

endmodule
