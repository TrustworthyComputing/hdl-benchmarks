module mmult (a_0_0, b_0_0, a_0_1, b_0_1, a_0_2, b_0_2, a_0_3, b_0_3, a_0_4, b_0_4, a_0_5, b_0_5, a_0_6, b_0_6, a_0_7, b_0_7, a_0_8, b_0_8, a_0_9, b_0_9, a_0_10, b_0_10, a_0_11, b_0_11, a_0_12, b_0_12, a_0_13, b_0_13, a_0_14, b_0_14, a_1_0, b_1_0, a_1_1, b_1_1, a_1_2, b_1_2, a_1_3, b_1_3, a_1_4, b_1_4, a_1_5, b_1_5, a_1_6, b_1_6, a_1_7, b_1_7, a_1_8, b_1_8, a_1_9, b_1_9, a_1_10, b_1_10, a_1_11, b_1_11, a_1_12, b_1_12, a_1_13, b_1_13, a_1_14, b_1_14, a_2_0, b_2_0, a_2_1, b_2_1, a_2_2, b_2_2, a_2_3, b_2_3, a_2_4, b_2_4, a_2_5, b_2_5, a_2_6, b_2_6, a_2_7, b_2_7, a_2_8, b_2_8, a_2_9, b_2_9, a_2_10, b_2_10, a_2_11, b_2_11, a_2_12, b_2_12, a_2_13, b_2_13, a_2_14, b_2_14, a_3_0, b_3_0, a_3_1, b_3_1, a_3_2, b_3_2, a_3_3, b_3_3, a_3_4, b_3_4, a_3_5, b_3_5, a_3_6, b_3_6, a_3_7, b_3_7, a_3_8, b_3_8, a_3_9, b_3_9, a_3_10, b_3_10, a_3_11, b_3_11, a_3_12, b_3_12, a_3_13, b_3_13, a_3_14, b_3_14, a_4_0, b_4_0, a_4_1, b_4_1, a_4_2, b_4_2, a_4_3, b_4_3, a_4_4, b_4_4, a_4_5, b_4_5, a_4_6, b_4_6, a_4_7, b_4_7, a_4_8, b_4_8, a_4_9, b_4_9, a_4_10, b_4_10, a_4_11, b_4_11, a_4_12, b_4_12, a_4_13, b_4_13, a_4_14, b_4_14, a_5_0, b_5_0, a_5_1, b_5_1, a_5_2, b_5_2, a_5_3, b_5_3, a_5_4, b_5_4, a_5_5, b_5_5, a_5_6, b_5_6, a_5_7, b_5_7, a_5_8, b_5_8, a_5_9, b_5_9, a_5_10, b_5_10, a_5_11, b_5_11, a_5_12, b_5_12, a_5_13, b_5_13, a_5_14, b_5_14, a_6_0, b_6_0, a_6_1, b_6_1, a_6_2, b_6_2, a_6_3, b_6_3, a_6_4, b_6_4, a_6_5, b_6_5, a_6_6, b_6_6, a_6_7, b_6_7, a_6_8, b_6_8, a_6_9, b_6_9, a_6_10, b_6_10, a_6_11, b_6_11, a_6_12, b_6_12, a_6_13, b_6_13, a_6_14, b_6_14, a_7_0, b_7_0, a_7_1, b_7_1, a_7_2, b_7_2, a_7_3, b_7_3, a_7_4, b_7_4, a_7_5, b_7_5, a_7_6, b_7_6, a_7_7, b_7_7, a_7_8, b_7_8, a_7_9, b_7_9, a_7_10, b_7_10, a_7_11, b_7_11, a_7_12, b_7_12, a_7_13, b_7_13, a_7_14, b_7_14, a_8_0, b_8_0, a_8_1, b_8_1, a_8_2, b_8_2, a_8_3, b_8_3, a_8_4, b_8_4, a_8_5, b_8_5, a_8_6, b_8_6, a_8_7, b_8_7, a_8_8, b_8_8, a_8_9, b_8_9, a_8_10, b_8_10, a_8_11, b_8_11, a_8_12, b_8_12, a_8_13, b_8_13, a_8_14, b_8_14, a_9_0, b_9_0, a_9_1, b_9_1, a_9_2, b_9_2, a_9_3, b_9_3, a_9_4, b_9_4, a_9_5, b_9_5, a_9_6, b_9_6, a_9_7, b_9_7, a_9_8, b_9_8, a_9_9, b_9_9, a_9_10, b_9_10, a_9_11, b_9_11, a_9_12, b_9_12, a_9_13, b_9_13, a_9_14, b_9_14, a_10_0, b_10_0, a_10_1, b_10_1, a_10_2, b_10_2, a_10_3, b_10_3, a_10_4, b_10_4, a_10_5, b_10_5, a_10_6, b_10_6, a_10_7, b_10_7, a_10_8, b_10_8, a_10_9, b_10_9, a_10_10, b_10_10, a_10_11, b_10_11, a_10_12, b_10_12, a_10_13, b_10_13, a_10_14, b_10_14, a_11_0, b_11_0, a_11_1, b_11_1, a_11_2, b_11_2, a_11_3, b_11_3, a_11_4, b_11_4, a_11_5, b_11_5, a_11_6, b_11_6, a_11_7, b_11_7, a_11_8, b_11_8, a_11_9, b_11_9, a_11_10, b_11_10, a_11_11, b_11_11, a_11_12, b_11_12, a_11_13, b_11_13, a_11_14, b_11_14, a_12_0, b_12_0, a_12_1, b_12_1, a_12_2, b_12_2, a_12_3, b_12_3, a_12_4, b_12_4, a_12_5, b_12_5, a_12_6, b_12_6, a_12_7, b_12_7, a_12_8, b_12_8, a_12_9, b_12_9, a_12_10, b_12_10, a_12_11, b_12_11, a_12_12, b_12_12, a_12_13, b_12_13, a_12_14, b_12_14, a_13_0, b_13_0, a_13_1, b_13_1, a_13_2, b_13_2, a_13_3, b_13_3, a_13_4, b_13_4, a_13_5, b_13_5, a_13_6, b_13_6, a_13_7, b_13_7, a_13_8, b_13_8, a_13_9, b_13_9, a_13_10, b_13_10, a_13_11, b_13_11, a_13_12, b_13_12, a_13_13, b_13_13, a_13_14, b_13_14, a_14_0, b_14_0, a_14_1, b_14_1, a_14_2, b_14_2, a_14_3, b_14_3, a_14_4, b_14_4, a_14_5, b_14_5, a_14_6, b_14_6, a_14_7, b_14_7, a_14_8, b_14_8, a_14_9, b_14_9, a_14_10, b_14_10, a_14_11, b_14_11, a_14_12, b_14_12, a_14_13, b_14_13, a_14_14, b_14_14, c_0_0, c_0_1, c_0_2, c_0_3, c_0_4, c_0_5, c_0_6, c_0_7, c_0_8, c_0_9, c_0_10, c_0_11, c_0_12, c_0_13, c_0_14, c_1_0, c_1_1, c_1_2, c_1_3, c_1_4, c_1_5, c_1_6, c_1_7, c_1_8, c_1_9, c_1_10, c_1_11, c_1_12, c_1_13, c_1_14, c_2_0, c_2_1, c_2_2, c_2_3, c_2_4, c_2_5, c_2_6, c_2_7, c_2_8, c_2_9, c_2_10, c_2_11, c_2_12, c_2_13, c_2_14, c_3_0, c_3_1, c_3_2, c_3_3, c_3_4, c_3_5, c_3_6, c_3_7, c_3_8, c_3_9, c_3_10, c_3_11, c_3_12, c_3_13, c_3_14, c_4_0, c_4_1, c_4_2, c_4_3, c_4_4, c_4_5, c_4_6, c_4_7, c_4_8, c_4_9, c_4_10, c_4_11, c_4_12, c_4_13, c_4_14, c_5_0, c_5_1, c_5_2, c_5_3, c_5_4, c_5_5, c_5_6, c_5_7, c_5_8, c_5_9, c_5_10, c_5_11, c_5_12, c_5_13, c_5_14, c_6_0, c_6_1, c_6_2, c_6_3, c_6_4, c_6_5, c_6_6, c_6_7, c_6_8, c_6_9, c_6_10, c_6_11, c_6_12, c_6_13, c_6_14, c_7_0, c_7_1, c_7_2, c_7_3, c_7_4, c_7_5, c_7_6, c_7_7, c_7_8, c_7_9, c_7_10, c_7_11, c_7_12, c_7_13, c_7_14, c_8_0, c_8_1, c_8_2, c_8_3, c_8_4, c_8_5, c_8_6, c_8_7, c_8_8, c_8_9, c_8_10, c_8_11, c_8_12, c_8_13, c_8_14, c_9_0, c_9_1, c_9_2, c_9_3, c_9_4, c_9_5, c_9_6, c_9_7, c_9_8, c_9_9, c_9_10, c_9_11, c_9_12, c_9_13, c_9_14, c_10_0, c_10_1, c_10_2, c_10_3, c_10_4, c_10_5, c_10_6, c_10_7, c_10_8, c_10_9, c_10_10, c_10_11, c_10_12, c_10_13, c_10_14, c_11_0, c_11_1, c_11_2, c_11_3, c_11_4, c_11_5, c_11_6, c_11_7, c_11_8, c_11_9, c_11_10, c_11_11, c_11_12, c_11_13, c_11_14, c_12_0, c_12_1, c_12_2, c_12_3, c_12_4, c_12_5, c_12_6, c_12_7, c_12_8, c_12_9, c_12_10, c_12_11, c_12_12, c_12_13, c_12_14, c_13_0, c_13_1, c_13_2, c_13_3, c_13_4, c_13_5, c_13_6, c_13_7, c_13_8, c_13_9, c_13_10, c_13_11, c_13_12, c_13_13, c_13_14, c_14_0, c_14_1, c_14_2, c_14_3, c_14_4, c_14_5, c_14_6, c_14_7, c_14_8, c_14_9, c_14_10, c_14_11, c_14_12, c_14_13, c_14_14);

  input [15:0] a_0_0;
  input [15:0] b_0_0;
  input [15:0] a_0_1;
  input [15:0] b_0_1;
  input [15:0] a_0_2;
  input [15:0] b_0_2;
  input [15:0] a_0_3;
  input [15:0] b_0_3;
  input [15:0] a_0_4;
  input [15:0] b_0_4;
  input [15:0] a_0_5;
  input [15:0] b_0_5;
  input [15:0] a_0_6;
  input [15:0] b_0_6;
  input [15:0] a_0_7;
  input [15:0] b_0_7;
  input [15:0] a_0_8;
  input [15:0] b_0_8;
  input [15:0] a_0_9;
  input [15:0] b_0_9;
  input [15:0] a_0_10;
  input [15:0] b_0_10;
  input [15:0] a_0_11;
  input [15:0] b_0_11;
  input [15:0] a_0_12;
  input [15:0] b_0_12;
  input [15:0] a_0_13;
  input [15:0] b_0_13;
  input [15:0] a_0_14;
  input [15:0] b_0_14;
  input [15:0] a_1_0;
  input [15:0] b_1_0;
  input [15:0] a_1_1;
  input [15:0] b_1_1;
  input [15:0] a_1_2;
  input [15:0] b_1_2;
  input [15:0] a_1_3;
  input [15:0] b_1_3;
  input [15:0] a_1_4;
  input [15:0] b_1_4;
  input [15:0] a_1_5;
  input [15:0] b_1_5;
  input [15:0] a_1_6;
  input [15:0] b_1_6;
  input [15:0] a_1_7;
  input [15:0] b_1_7;
  input [15:0] a_1_8;
  input [15:0] b_1_8;
  input [15:0] a_1_9;
  input [15:0] b_1_9;
  input [15:0] a_1_10;
  input [15:0] b_1_10;
  input [15:0] a_1_11;
  input [15:0] b_1_11;
  input [15:0] a_1_12;
  input [15:0] b_1_12;
  input [15:0] a_1_13;
  input [15:0] b_1_13;
  input [15:0] a_1_14;
  input [15:0] b_1_14;
  input [15:0] a_2_0;
  input [15:0] b_2_0;
  input [15:0] a_2_1;
  input [15:0] b_2_1;
  input [15:0] a_2_2;
  input [15:0] b_2_2;
  input [15:0] a_2_3;
  input [15:0] b_2_3;
  input [15:0] a_2_4;
  input [15:0] b_2_4;
  input [15:0] a_2_5;
  input [15:0] b_2_5;
  input [15:0] a_2_6;
  input [15:0] b_2_6;
  input [15:0] a_2_7;
  input [15:0] b_2_7;
  input [15:0] a_2_8;
  input [15:0] b_2_8;
  input [15:0] a_2_9;
  input [15:0] b_2_9;
  input [15:0] a_2_10;
  input [15:0] b_2_10;
  input [15:0] a_2_11;
  input [15:0] b_2_11;
  input [15:0] a_2_12;
  input [15:0] b_2_12;
  input [15:0] a_2_13;
  input [15:0] b_2_13;
  input [15:0] a_2_14;
  input [15:0] b_2_14;
  input [15:0] a_3_0;
  input [15:0] b_3_0;
  input [15:0] a_3_1;
  input [15:0] b_3_1;
  input [15:0] a_3_2;
  input [15:0] b_3_2;
  input [15:0] a_3_3;
  input [15:0] b_3_3;
  input [15:0] a_3_4;
  input [15:0] b_3_4;
  input [15:0] a_3_5;
  input [15:0] b_3_5;
  input [15:0] a_3_6;
  input [15:0] b_3_6;
  input [15:0] a_3_7;
  input [15:0] b_3_7;
  input [15:0] a_3_8;
  input [15:0] b_3_8;
  input [15:0] a_3_9;
  input [15:0] b_3_9;
  input [15:0] a_3_10;
  input [15:0] b_3_10;
  input [15:0] a_3_11;
  input [15:0] b_3_11;
  input [15:0] a_3_12;
  input [15:0] b_3_12;
  input [15:0] a_3_13;
  input [15:0] b_3_13;
  input [15:0] a_3_14;
  input [15:0] b_3_14;
  input [15:0] a_4_0;
  input [15:0] b_4_0;
  input [15:0] a_4_1;
  input [15:0] b_4_1;
  input [15:0] a_4_2;
  input [15:0] b_4_2;
  input [15:0] a_4_3;
  input [15:0] b_4_3;
  input [15:0] a_4_4;
  input [15:0] b_4_4;
  input [15:0] a_4_5;
  input [15:0] b_4_5;
  input [15:0] a_4_6;
  input [15:0] b_4_6;
  input [15:0] a_4_7;
  input [15:0] b_4_7;
  input [15:0] a_4_8;
  input [15:0] b_4_8;
  input [15:0] a_4_9;
  input [15:0] b_4_9;
  input [15:0] a_4_10;
  input [15:0] b_4_10;
  input [15:0] a_4_11;
  input [15:0] b_4_11;
  input [15:0] a_4_12;
  input [15:0] b_4_12;
  input [15:0] a_4_13;
  input [15:0] b_4_13;
  input [15:0] a_4_14;
  input [15:0] b_4_14;
  input [15:0] a_5_0;
  input [15:0] b_5_0;
  input [15:0] a_5_1;
  input [15:0] b_5_1;
  input [15:0] a_5_2;
  input [15:0] b_5_2;
  input [15:0] a_5_3;
  input [15:0] b_5_3;
  input [15:0] a_5_4;
  input [15:0] b_5_4;
  input [15:0] a_5_5;
  input [15:0] b_5_5;
  input [15:0] a_5_6;
  input [15:0] b_5_6;
  input [15:0] a_5_7;
  input [15:0] b_5_7;
  input [15:0] a_5_8;
  input [15:0] b_5_8;
  input [15:0] a_5_9;
  input [15:0] b_5_9;
  input [15:0] a_5_10;
  input [15:0] b_5_10;
  input [15:0] a_5_11;
  input [15:0] b_5_11;
  input [15:0] a_5_12;
  input [15:0] b_5_12;
  input [15:0] a_5_13;
  input [15:0] b_5_13;
  input [15:0] a_5_14;
  input [15:0] b_5_14;
  input [15:0] a_6_0;
  input [15:0] b_6_0;
  input [15:0] a_6_1;
  input [15:0] b_6_1;
  input [15:0] a_6_2;
  input [15:0] b_6_2;
  input [15:0] a_6_3;
  input [15:0] b_6_3;
  input [15:0] a_6_4;
  input [15:0] b_6_4;
  input [15:0] a_6_5;
  input [15:0] b_6_5;
  input [15:0] a_6_6;
  input [15:0] b_6_6;
  input [15:0] a_6_7;
  input [15:0] b_6_7;
  input [15:0] a_6_8;
  input [15:0] b_6_8;
  input [15:0] a_6_9;
  input [15:0] b_6_9;
  input [15:0] a_6_10;
  input [15:0] b_6_10;
  input [15:0] a_6_11;
  input [15:0] b_6_11;
  input [15:0] a_6_12;
  input [15:0] b_6_12;
  input [15:0] a_6_13;
  input [15:0] b_6_13;
  input [15:0] a_6_14;
  input [15:0] b_6_14;
  input [15:0] a_7_0;
  input [15:0] b_7_0;
  input [15:0] a_7_1;
  input [15:0] b_7_1;
  input [15:0] a_7_2;
  input [15:0] b_7_2;
  input [15:0] a_7_3;
  input [15:0] b_7_3;
  input [15:0] a_7_4;
  input [15:0] b_7_4;
  input [15:0] a_7_5;
  input [15:0] b_7_5;
  input [15:0] a_7_6;
  input [15:0] b_7_6;
  input [15:0] a_7_7;
  input [15:0] b_7_7;
  input [15:0] a_7_8;
  input [15:0] b_7_8;
  input [15:0] a_7_9;
  input [15:0] b_7_9;
  input [15:0] a_7_10;
  input [15:0] b_7_10;
  input [15:0] a_7_11;
  input [15:0] b_7_11;
  input [15:0] a_7_12;
  input [15:0] b_7_12;
  input [15:0] a_7_13;
  input [15:0] b_7_13;
  input [15:0] a_7_14;
  input [15:0] b_7_14;
  input [15:0] a_8_0;
  input [15:0] b_8_0;
  input [15:0] a_8_1;
  input [15:0] b_8_1;
  input [15:0] a_8_2;
  input [15:0] b_8_2;
  input [15:0] a_8_3;
  input [15:0] b_8_3;
  input [15:0] a_8_4;
  input [15:0] b_8_4;
  input [15:0] a_8_5;
  input [15:0] b_8_5;
  input [15:0] a_8_6;
  input [15:0] b_8_6;
  input [15:0] a_8_7;
  input [15:0] b_8_7;
  input [15:0] a_8_8;
  input [15:0] b_8_8;
  input [15:0] a_8_9;
  input [15:0] b_8_9;
  input [15:0] a_8_10;
  input [15:0] b_8_10;
  input [15:0] a_8_11;
  input [15:0] b_8_11;
  input [15:0] a_8_12;
  input [15:0] b_8_12;
  input [15:0] a_8_13;
  input [15:0] b_8_13;
  input [15:0] a_8_14;
  input [15:0] b_8_14;
  input [15:0] a_9_0;
  input [15:0] b_9_0;
  input [15:0] a_9_1;
  input [15:0] b_9_1;
  input [15:0] a_9_2;
  input [15:0] b_9_2;
  input [15:0] a_9_3;
  input [15:0] b_9_3;
  input [15:0] a_9_4;
  input [15:0] b_9_4;
  input [15:0] a_9_5;
  input [15:0] b_9_5;
  input [15:0] a_9_6;
  input [15:0] b_9_6;
  input [15:0] a_9_7;
  input [15:0] b_9_7;
  input [15:0] a_9_8;
  input [15:0] b_9_8;
  input [15:0] a_9_9;
  input [15:0] b_9_9;
  input [15:0] a_9_10;
  input [15:0] b_9_10;
  input [15:0] a_9_11;
  input [15:0] b_9_11;
  input [15:0] a_9_12;
  input [15:0] b_9_12;
  input [15:0] a_9_13;
  input [15:0] b_9_13;
  input [15:0] a_9_14;
  input [15:0] b_9_14;
  input [15:0] a_10_0;
  input [15:0] b_10_0;
  input [15:0] a_10_1;
  input [15:0] b_10_1;
  input [15:0] a_10_2;
  input [15:0] b_10_2;
  input [15:0] a_10_3;
  input [15:0] b_10_3;
  input [15:0] a_10_4;
  input [15:0] b_10_4;
  input [15:0] a_10_5;
  input [15:0] b_10_5;
  input [15:0] a_10_6;
  input [15:0] b_10_6;
  input [15:0] a_10_7;
  input [15:0] b_10_7;
  input [15:0] a_10_8;
  input [15:0] b_10_8;
  input [15:0] a_10_9;
  input [15:0] b_10_9;
  input [15:0] a_10_10;
  input [15:0] b_10_10;
  input [15:0] a_10_11;
  input [15:0] b_10_11;
  input [15:0] a_10_12;
  input [15:0] b_10_12;
  input [15:0] a_10_13;
  input [15:0] b_10_13;
  input [15:0] a_10_14;
  input [15:0] b_10_14;
  input [15:0] a_11_0;
  input [15:0] b_11_0;
  input [15:0] a_11_1;
  input [15:0] b_11_1;
  input [15:0] a_11_2;
  input [15:0] b_11_2;
  input [15:0] a_11_3;
  input [15:0] b_11_3;
  input [15:0] a_11_4;
  input [15:0] b_11_4;
  input [15:0] a_11_5;
  input [15:0] b_11_5;
  input [15:0] a_11_6;
  input [15:0] b_11_6;
  input [15:0] a_11_7;
  input [15:0] b_11_7;
  input [15:0] a_11_8;
  input [15:0] b_11_8;
  input [15:0] a_11_9;
  input [15:0] b_11_9;
  input [15:0] a_11_10;
  input [15:0] b_11_10;
  input [15:0] a_11_11;
  input [15:0] b_11_11;
  input [15:0] a_11_12;
  input [15:0] b_11_12;
  input [15:0] a_11_13;
  input [15:0] b_11_13;
  input [15:0] a_11_14;
  input [15:0] b_11_14;
  input [15:0] a_12_0;
  input [15:0] b_12_0;
  input [15:0] a_12_1;
  input [15:0] b_12_1;
  input [15:0] a_12_2;
  input [15:0] b_12_2;
  input [15:0] a_12_3;
  input [15:0] b_12_3;
  input [15:0] a_12_4;
  input [15:0] b_12_4;
  input [15:0] a_12_5;
  input [15:0] b_12_5;
  input [15:0] a_12_6;
  input [15:0] b_12_6;
  input [15:0] a_12_7;
  input [15:0] b_12_7;
  input [15:0] a_12_8;
  input [15:0] b_12_8;
  input [15:0] a_12_9;
  input [15:0] b_12_9;
  input [15:0] a_12_10;
  input [15:0] b_12_10;
  input [15:0] a_12_11;
  input [15:0] b_12_11;
  input [15:0] a_12_12;
  input [15:0] b_12_12;
  input [15:0] a_12_13;
  input [15:0] b_12_13;
  input [15:0] a_12_14;
  input [15:0] b_12_14;
  input [15:0] a_13_0;
  input [15:0] b_13_0;
  input [15:0] a_13_1;
  input [15:0] b_13_1;
  input [15:0] a_13_2;
  input [15:0] b_13_2;
  input [15:0] a_13_3;
  input [15:0] b_13_3;
  input [15:0] a_13_4;
  input [15:0] b_13_4;
  input [15:0] a_13_5;
  input [15:0] b_13_5;
  input [15:0] a_13_6;
  input [15:0] b_13_6;
  input [15:0] a_13_7;
  input [15:0] b_13_7;
  input [15:0] a_13_8;
  input [15:0] b_13_8;
  input [15:0] a_13_9;
  input [15:0] b_13_9;
  input [15:0] a_13_10;
  input [15:0] b_13_10;
  input [15:0] a_13_11;
  input [15:0] b_13_11;
  input [15:0] a_13_12;
  input [15:0] b_13_12;
  input [15:0] a_13_13;
  input [15:0] b_13_13;
  input [15:0] a_13_14;
  input [15:0] b_13_14;
  input [15:0] a_14_0;
  input [15:0] b_14_0;
  input [15:0] a_14_1;
  input [15:0] b_14_1;
  input [15:0] a_14_2;
  input [15:0] b_14_2;
  input [15:0] a_14_3;
  input [15:0] b_14_3;
  input [15:0] a_14_4;
  input [15:0] b_14_4;
  input [15:0] a_14_5;
  input [15:0] b_14_5;
  input [15:0] a_14_6;
  input [15:0] b_14_6;
  input [15:0] a_14_7;
  input [15:0] b_14_7;
  input [15:0] a_14_8;
  input [15:0] b_14_8;
  input [15:0] a_14_9;
  input [15:0] b_14_9;
  input [15:0] a_14_10;
  input [15:0] b_14_10;
  input [15:0] a_14_11;
  input [15:0] b_14_11;
  input [15:0] a_14_12;
  input [15:0] b_14_12;
  input [15:0] a_14_13;
  input [15:0] b_14_13;
  input [15:0] a_14_14;
  input [15:0] b_14_14;

  output [15:0] c_0_0;
  output [15:0] c_0_1;
  output [15:0] c_0_2;
  output [15:0] c_0_3;
  output [15:0] c_0_4;
  output [15:0] c_0_5;
  output [15:0] c_0_6;
  output [15:0] c_0_7;
  output [15:0] c_0_8;
  output [15:0] c_0_9;
  output [15:0] c_0_10;
  output [15:0] c_0_11;
  output [15:0] c_0_12;
  output [15:0] c_0_13;
  output [15:0] c_0_14;
  output [15:0] c_1_0;
  output [15:0] c_1_1;
  output [15:0] c_1_2;
  output [15:0] c_1_3;
  output [15:0] c_1_4;
  output [15:0] c_1_5;
  output [15:0] c_1_6;
  output [15:0] c_1_7;
  output [15:0] c_1_8;
  output [15:0] c_1_9;
  output [15:0] c_1_10;
  output [15:0] c_1_11;
  output [15:0] c_1_12;
  output [15:0] c_1_13;
  output [15:0] c_1_14;
  output [15:0] c_2_0;
  output [15:0] c_2_1;
  output [15:0] c_2_2;
  output [15:0] c_2_3;
  output [15:0] c_2_4;
  output [15:0] c_2_5;
  output [15:0] c_2_6;
  output [15:0] c_2_7;
  output [15:0] c_2_8;
  output [15:0] c_2_9;
  output [15:0] c_2_10;
  output [15:0] c_2_11;
  output [15:0] c_2_12;
  output [15:0] c_2_13;
  output [15:0] c_2_14;
  output [15:0] c_3_0;
  output [15:0] c_3_1;
  output [15:0] c_3_2;
  output [15:0] c_3_3;
  output [15:0] c_3_4;
  output [15:0] c_3_5;
  output [15:0] c_3_6;
  output [15:0] c_3_7;
  output [15:0] c_3_8;
  output [15:0] c_3_9;
  output [15:0] c_3_10;
  output [15:0] c_3_11;
  output [15:0] c_3_12;
  output [15:0] c_3_13;
  output [15:0] c_3_14;
  output [15:0] c_4_0;
  output [15:0] c_4_1;
  output [15:0] c_4_2;
  output [15:0] c_4_3;
  output [15:0] c_4_4;
  output [15:0] c_4_5;
  output [15:0] c_4_6;
  output [15:0] c_4_7;
  output [15:0] c_4_8;
  output [15:0] c_4_9;
  output [15:0] c_4_10;
  output [15:0] c_4_11;
  output [15:0] c_4_12;
  output [15:0] c_4_13;
  output [15:0] c_4_14;
  output [15:0] c_5_0;
  output [15:0] c_5_1;
  output [15:0] c_5_2;
  output [15:0] c_5_3;
  output [15:0] c_5_4;
  output [15:0] c_5_5;
  output [15:0] c_5_6;
  output [15:0] c_5_7;
  output [15:0] c_5_8;
  output [15:0] c_5_9;
  output [15:0] c_5_10;
  output [15:0] c_5_11;
  output [15:0] c_5_12;
  output [15:0] c_5_13;
  output [15:0] c_5_14;
  output [15:0] c_6_0;
  output [15:0] c_6_1;
  output [15:0] c_6_2;
  output [15:0] c_6_3;
  output [15:0] c_6_4;
  output [15:0] c_6_5;
  output [15:0] c_6_6;
  output [15:0] c_6_7;
  output [15:0] c_6_8;
  output [15:0] c_6_9;
  output [15:0] c_6_10;
  output [15:0] c_6_11;
  output [15:0] c_6_12;
  output [15:0] c_6_13;
  output [15:0] c_6_14;
  output [15:0] c_7_0;
  output [15:0] c_7_1;
  output [15:0] c_7_2;
  output [15:0] c_7_3;
  output [15:0] c_7_4;
  output [15:0] c_7_5;
  output [15:0] c_7_6;
  output [15:0] c_7_7;
  output [15:0] c_7_8;
  output [15:0] c_7_9;
  output [15:0] c_7_10;
  output [15:0] c_7_11;
  output [15:0] c_7_12;
  output [15:0] c_7_13;
  output [15:0] c_7_14;
  output [15:0] c_8_0;
  output [15:0] c_8_1;
  output [15:0] c_8_2;
  output [15:0] c_8_3;
  output [15:0] c_8_4;
  output [15:0] c_8_5;
  output [15:0] c_8_6;
  output [15:0] c_8_7;
  output [15:0] c_8_8;
  output [15:0] c_8_9;
  output [15:0] c_8_10;
  output [15:0] c_8_11;
  output [15:0] c_8_12;
  output [15:0] c_8_13;
  output [15:0] c_8_14;
  output [15:0] c_9_0;
  output [15:0] c_9_1;
  output [15:0] c_9_2;
  output [15:0] c_9_3;
  output [15:0] c_9_4;
  output [15:0] c_9_5;
  output [15:0] c_9_6;
  output [15:0] c_9_7;
  output [15:0] c_9_8;
  output [15:0] c_9_9;
  output [15:0] c_9_10;
  output [15:0] c_9_11;
  output [15:0] c_9_12;
  output [15:0] c_9_13;
  output [15:0] c_9_14;
  output [15:0] c_10_0;
  output [15:0] c_10_1;
  output [15:0] c_10_2;
  output [15:0] c_10_3;
  output [15:0] c_10_4;
  output [15:0] c_10_5;
  output [15:0] c_10_6;
  output [15:0] c_10_7;
  output [15:0] c_10_8;
  output [15:0] c_10_9;
  output [15:0] c_10_10;
  output [15:0] c_10_11;
  output [15:0] c_10_12;
  output [15:0] c_10_13;
  output [15:0] c_10_14;
  output [15:0] c_11_0;
  output [15:0] c_11_1;
  output [15:0] c_11_2;
  output [15:0] c_11_3;
  output [15:0] c_11_4;
  output [15:0] c_11_5;
  output [15:0] c_11_6;
  output [15:0] c_11_7;
  output [15:0] c_11_8;
  output [15:0] c_11_9;
  output [15:0] c_11_10;
  output [15:0] c_11_11;
  output [15:0] c_11_12;
  output [15:0] c_11_13;
  output [15:0] c_11_14;
  output [15:0] c_12_0;
  output [15:0] c_12_1;
  output [15:0] c_12_2;
  output [15:0] c_12_3;
  output [15:0] c_12_4;
  output [15:0] c_12_5;
  output [15:0] c_12_6;
  output [15:0] c_12_7;
  output [15:0] c_12_8;
  output [15:0] c_12_9;
  output [15:0] c_12_10;
  output [15:0] c_12_11;
  output [15:0] c_12_12;
  output [15:0] c_12_13;
  output [15:0] c_12_14;
  output [15:0] c_13_0;
  output [15:0] c_13_1;
  output [15:0] c_13_2;
  output [15:0] c_13_3;
  output [15:0] c_13_4;
  output [15:0] c_13_5;
  output [15:0] c_13_6;
  output [15:0] c_13_7;
  output [15:0] c_13_8;
  output [15:0] c_13_9;
  output [15:0] c_13_10;
  output [15:0] c_13_11;
  output [15:0] c_13_12;
  output [15:0] c_13_13;
  output [15:0] c_13_14;
  output [15:0] c_14_0;
  output [15:0] c_14_1;
  output [15:0] c_14_2;
  output [15:0] c_14_3;
  output [15:0] c_14_4;
  output [15:0] c_14_5;
  output [15:0] c_14_6;
  output [15:0] c_14_7;
  output [15:0] c_14_8;
  output [15:0] c_14_9;
  output [15:0] c_14_10;
  output [15:0] c_14_11;
  output [15:0] c_14_12;
  output [15:0] c_14_13;
  output [15:0] c_14_14;

  wire [15:0] t0_r0_c0_rr0;
  wire [15:0] t0_r0_c0_rr1;
  wire [15:0] t0_r0_c0_rr2;
  wire [15:0] t0_r0_c0_rr3;
  wire [15:0] t0_r0_c0_rr4;
  wire [15:0] t0_r0_c0_rr5;
  wire [15:0] t0_r0_c0_rr6;
  wire [15:0] t0_r0_c0_rr7;
  wire [15:0] t0_r0_c0_rr8;
  wire [15:0] t0_r0_c0_rr9;
  wire [15:0] t0_r0_c0_rr10;
  wire [15:0] t0_r0_c0_rr11;
  wire [15:0] t0_r0_c0_rr12;
  wire [15:0] t0_r0_c0_rr13;
  wire [15:0] t0_r0_c0_rr14;
  wire [15:0] t1_r0_c0_rr0;
  wire [15:0] t1_r0_c0_rr1;
  wire [15:0] t1_r0_c0_rr2;
  wire [15:0] t1_r0_c0_rr3;
  wire [15:0] t1_r0_c0_rr4;
  wire [15:0] t1_r0_c0_rr5;
  wire [15:0] t1_r0_c0_rr6;
  wire [15:0] t1_r0_c0_rr7;
  wire [15:0] t2_r0_c0_rr0;
  wire [15:0] t2_r0_c0_rr1;
  wire [15:0] t2_r0_c0_rr2;
  wire [15:0] t2_r0_c0_rr3;
  wire [15:0] t3_r0_c0_rr0;
  wire [15:0] t3_r0_c0_rr1;
  wire [15:0] t4_r0_c0_rr0;
  wire [15:0] t0_r0_c1_rr0;
  wire [15:0] t0_r0_c1_rr1;
  wire [15:0] t0_r0_c1_rr2;
  wire [15:0] t0_r0_c1_rr3;
  wire [15:0] t0_r0_c1_rr4;
  wire [15:0] t0_r0_c1_rr5;
  wire [15:0] t0_r0_c1_rr6;
  wire [15:0] t0_r0_c1_rr7;
  wire [15:0] t0_r0_c1_rr8;
  wire [15:0] t0_r0_c1_rr9;
  wire [15:0] t0_r0_c1_rr10;
  wire [15:0] t0_r0_c1_rr11;
  wire [15:0] t0_r0_c1_rr12;
  wire [15:0] t0_r0_c1_rr13;
  wire [15:0] t0_r0_c1_rr14;
  wire [15:0] t1_r0_c1_rr0;
  wire [15:0] t1_r0_c1_rr1;
  wire [15:0] t1_r0_c1_rr2;
  wire [15:0] t1_r0_c1_rr3;
  wire [15:0] t1_r0_c1_rr4;
  wire [15:0] t1_r0_c1_rr5;
  wire [15:0] t1_r0_c1_rr6;
  wire [15:0] t1_r0_c1_rr7;
  wire [15:0] t2_r0_c1_rr0;
  wire [15:0] t2_r0_c1_rr1;
  wire [15:0] t2_r0_c1_rr2;
  wire [15:0] t2_r0_c1_rr3;
  wire [15:0] t3_r0_c1_rr0;
  wire [15:0] t3_r0_c1_rr1;
  wire [15:0] t4_r0_c1_rr0;
  wire [15:0] t0_r0_c2_rr0;
  wire [15:0] t0_r0_c2_rr1;
  wire [15:0] t0_r0_c2_rr2;
  wire [15:0] t0_r0_c2_rr3;
  wire [15:0] t0_r0_c2_rr4;
  wire [15:0] t0_r0_c2_rr5;
  wire [15:0] t0_r0_c2_rr6;
  wire [15:0] t0_r0_c2_rr7;
  wire [15:0] t0_r0_c2_rr8;
  wire [15:0] t0_r0_c2_rr9;
  wire [15:0] t0_r0_c2_rr10;
  wire [15:0] t0_r0_c2_rr11;
  wire [15:0] t0_r0_c2_rr12;
  wire [15:0] t0_r0_c2_rr13;
  wire [15:0] t0_r0_c2_rr14;
  wire [15:0] t1_r0_c2_rr0;
  wire [15:0] t1_r0_c2_rr1;
  wire [15:0] t1_r0_c2_rr2;
  wire [15:0] t1_r0_c2_rr3;
  wire [15:0] t1_r0_c2_rr4;
  wire [15:0] t1_r0_c2_rr5;
  wire [15:0] t1_r0_c2_rr6;
  wire [15:0] t1_r0_c2_rr7;
  wire [15:0] t2_r0_c2_rr0;
  wire [15:0] t2_r0_c2_rr1;
  wire [15:0] t2_r0_c2_rr2;
  wire [15:0] t2_r0_c2_rr3;
  wire [15:0] t3_r0_c2_rr0;
  wire [15:0] t3_r0_c2_rr1;
  wire [15:0] t4_r0_c2_rr0;
  wire [15:0] t0_r0_c3_rr0;
  wire [15:0] t0_r0_c3_rr1;
  wire [15:0] t0_r0_c3_rr2;
  wire [15:0] t0_r0_c3_rr3;
  wire [15:0] t0_r0_c3_rr4;
  wire [15:0] t0_r0_c3_rr5;
  wire [15:0] t0_r0_c3_rr6;
  wire [15:0] t0_r0_c3_rr7;
  wire [15:0] t0_r0_c3_rr8;
  wire [15:0] t0_r0_c3_rr9;
  wire [15:0] t0_r0_c3_rr10;
  wire [15:0] t0_r0_c3_rr11;
  wire [15:0] t0_r0_c3_rr12;
  wire [15:0] t0_r0_c3_rr13;
  wire [15:0] t0_r0_c3_rr14;
  wire [15:0] t1_r0_c3_rr0;
  wire [15:0] t1_r0_c3_rr1;
  wire [15:0] t1_r0_c3_rr2;
  wire [15:0] t1_r0_c3_rr3;
  wire [15:0] t1_r0_c3_rr4;
  wire [15:0] t1_r0_c3_rr5;
  wire [15:0] t1_r0_c3_rr6;
  wire [15:0] t1_r0_c3_rr7;
  wire [15:0] t2_r0_c3_rr0;
  wire [15:0] t2_r0_c3_rr1;
  wire [15:0] t2_r0_c3_rr2;
  wire [15:0] t2_r0_c3_rr3;
  wire [15:0] t3_r0_c3_rr0;
  wire [15:0] t3_r0_c3_rr1;
  wire [15:0] t4_r0_c3_rr0;
  wire [15:0] t0_r0_c4_rr0;
  wire [15:0] t0_r0_c4_rr1;
  wire [15:0] t0_r0_c4_rr2;
  wire [15:0] t0_r0_c4_rr3;
  wire [15:0] t0_r0_c4_rr4;
  wire [15:0] t0_r0_c4_rr5;
  wire [15:0] t0_r0_c4_rr6;
  wire [15:0] t0_r0_c4_rr7;
  wire [15:0] t0_r0_c4_rr8;
  wire [15:0] t0_r0_c4_rr9;
  wire [15:0] t0_r0_c4_rr10;
  wire [15:0] t0_r0_c4_rr11;
  wire [15:0] t0_r0_c4_rr12;
  wire [15:0] t0_r0_c4_rr13;
  wire [15:0] t0_r0_c4_rr14;
  wire [15:0] t1_r0_c4_rr0;
  wire [15:0] t1_r0_c4_rr1;
  wire [15:0] t1_r0_c4_rr2;
  wire [15:0] t1_r0_c4_rr3;
  wire [15:0] t1_r0_c4_rr4;
  wire [15:0] t1_r0_c4_rr5;
  wire [15:0] t1_r0_c4_rr6;
  wire [15:0] t1_r0_c4_rr7;
  wire [15:0] t2_r0_c4_rr0;
  wire [15:0] t2_r0_c4_rr1;
  wire [15:0] t2_r0_c4_rr2;
  wire [15:0] t2_r0_c4_rr3;
  wire [15:0] t3_r0_c4_rr0;
  wire [15:0] t3_r0_c4_rr1;
  wire [15:0] t4_r0_c4_rr0;
  wire [15:0] t0_r0_c5_rr0;
  wire [15:0] t0_r0_c5_rr1;
  wire [15:0] t0_r0_c5_rr2;
  wire [15:0] t0_r0_c5_rr3;
  wire [15:0] t0_r0_c5_rr4;
  wire [15:0] t0_r0_c5_rr5;
  wire [15:0] t0_r0_c5_rr6;
  wire [15:0] t0_r0_c5_rr7;
  wire [15:0] t0_r0_c5_rr8;
  wire [15:0] t0_r0_c5_rr9;
  wire [15:0] t0_r0_c5_rr10;
  wire [15:0] t0_r0_c5_rr11;
  wire [15:0] t0_r0_c5_rr12;
  wire [15:0] t0_r0_c5_rr13;
  wire [15:0] t0_r0_c5_rr14;
  wire [15:0] t1_r0_c5_rr0;
  wire [15:0] t1_r0_c5_rr1;
  wire [15:0] t1_r0_c5_rr2;
  wire [15:0] t1_r0_c5_rr3;
  wire [15:0] t1_r0_c5_rr4;
  wire [15:0] t1_r0_c5_rr5;
  wire [15:0] t1_r0_c5_rr6;
  wire [15:0] t1_r0_c5_rr7;
  wire [15:0] t2_r0_c5_rr0;
  wire [15:0] t2_r0_c5_rr1;
  wire [15:0] t2_r0_c5_rr2;
  wire [15:0] t2_r0_c5_rr3;
  wire [15:0] t3_r0_c5_rr0;
  wire [15:0] t3_r0_c5_rr1;
  wire [15:0] t4_r0_c5_rr0;
  wire [15:0] t0_r0_c6_rr0;
  wire [15:0] t0_r0_c6_rr1;
  wire [15:0] t0_r0_c6_rr2;
  wire [15:0] t0_r0_c6_rr3;
  wire [15:0] t0_r0_c6_rr4;
  wire [15:0] t0_r0_c6_rr5;
  wire [15:0] t0_r0_c6_rr6;
  wire [15:0] t0_r0_c6_rr7;
  wire [15:0] t0_r0_c6_rr8;
  wire [15:0] t0_r0_c6_rr9;
  wire [15:0] t0_r0_c6_rr10;
  wire [15:0] t0_r0_c6_rr11;
  wire [15:0] t0_r0_c6_rr12;
  wire [15:0] t0_r0_c6_rr13;
  wire [15:0] t0_r0_c6_rr14;
  wire [15:0] t1_r0_c6_rr0;
  wire [15:0] t1_r0_c6_rr1;
  wire [15:0] t1_r0_c6_rr2;
  wire [15:0] t1_r0_c6_rr3;
  wire [15:0] t1_r0_c6_rr4;
  wire [15:0] t1_r0_c6_rr5;
  wire [15:0] t1_r0_c6_rr6;
  wire [15:0] t1_r0_c6_rr7;
  wire [15:0] t2_r0_c6_rr0;
  wire [15:0] t2_r0_c6_rr1;
  wire [15:0] t2_r0_c6_rr2;
  wire [15:0] t2_r0_c6_rr3;
  wire [15:0] t3_r0_c6_rr0;
  wire [15:0] t3_r0_c6_rr1;
  wire [15:0] t4_r0_c6_rr0;
  wire [15:0] t0_r0_c7_rr0;
  wire [15:0] t0_r0_c7_rr1;
  wire [15:0] t0_r0_c7_rr2;
  wire [15:0] t0_r0_c7_rr3;
  wire [15:0] t0_r0_c7_rr4;
  wire [15:0] t0_r0_c7_rr5;
  wire [15:0] t0_r0_c7_rr6;
  wire [15:0] t0_r0_c7_rr7;
  wire [15:0] t0_r0_c7_rr8;
  wire [15:0] t0_r0_c7_rr9;
  wire [15:0] t0_r0_c7_rr10;
  wire [15:0] t0_r0_c7_rr11;
  wire [15:0] t0_r0_c7_rr12;
  wire [15:0] t0_r0_c7_rr13;
  wire [15:0] t0_r0_c7_rr14;
  wire [15:0] t1_r0_c7_rr0;
  wire [15:0] t1_r0_c7_rr1;
  wire [15:0] t1_r0_c7_rr2;
  wire [15:0] t1_r0_c7_rr3;
  wire [15:0] t1_r0_c7_rr4;
  wire [15:0] t1_r0_c7_rr5;
  wire [15:0] t1_r0_c7_rr6;
  wire [15:0] t1_r0_c7_rr7;
  wire [15:0] t2_r0_c7_rr0;
  wire [15:0] t2_r0_c7_rr1;
  wire [15:0] t2_r0_c7_rr2;
  wire [15:0] t2_r0_c7_rr3;
  wire [15:0] t3_r0_c7_rr0;
  wire [15:0] t3_r0_c7_rr1;
  wire [15:0] t4_r0_c7_rr0;
  wire [15:0] t0_r0_c8_rr0;
  wire [15:0] t0_r0_c8_rr1;
  wire [15:0] t0_r0_c8_rr2;
  wire [15:0] t0_r0_c8_rr3;
  wire [15:0] t0_r0_c8_rr4;
  wire [15:0] t0_r0_c8_rr5;
  wire [15:0] t0_r0_c8_rr6;
  wire [15:0] t0_r0_c8_rr7;
  wire [15:0] t0_r0_c8_rr8;
  wire [15:0] t0_r0_c8_rr9;
  wire [15:0] t0_r0_c8_rr10;
  wire [15:0] t0_r0_c8_rr11;
  wire [15:0] t0_r0_c8_rr12;
  wire [15:0] t0_r0_c8_rr13;
  wire [15:0] t0_r0_c8_rr14;
  wire [15:0] t1_r0_c8_rr0;
  wire [15:0] t1_r0_c8_rr1;
  wire [15:0] t1_r0_c8_rr2;
  wire [15:0] t1_r0_c8_rr3;
  wire [15:0] t1_r0_c8_rr4;
  wire [15:0] t1_r0_c8_rr5;
  wire [15:0] t1_r0_c8_rr6;
  wire [15:0] t1_r0_c8_rr7;
  wire [15:0] t2_r0_c8_rr0;
  wire [15:0] t2_r0_c8_rr1;
  wire [15:0] t2_r0_c8_rr2;
  wire [15:0] t2_r0_c8_rr3;
  wire [15:0] t3_r0_c8_rr0;
  wire [15:0] t3_r0_c8_rr1;
  wire [15:0] t4_r0_c8_rr0;
  wire [15:0] t0_r0_c9_rr0;
  wire [15:0] t0_r0_c9_rr1;
  wire [15:0] t0_r0_c9_rr2;
  wire [15:0] t0_r0_c9_rr3;
  wire [15:0] t0_r0_c9_rr4;
  wire [15:0] t0_r0_c9_rr5;
  wire [15:0] t0_r0_c9_rr6;
  wire [15:0] t0_r0_c9_rr7;
  wire [15:0] t0_r0_c9_rr8;
  wire [15:0] t0_r0_c9_rr9;
  wire [15:0] t0_r0_c9_rr10;
  wire [15:0] t0_r0_c9_rr11;
  wire [15:0] t0_r0_c9_rr12;
  wire [15:0] t0_r0_c9_rr13;
  wire [15:0] t0_r0_c9_rr14;
  wire [15:0] t1_r0_c9_rr0;
  wire [15:0] t1_r0_c9_rr1;
  wire [15:0] t1_r0_c9_rr2;
  wire [15:0] t1_r0_c9_rr3;
  wire [15:0] t1_r0_c9_rr4;
  wire [15:0] t1_r0_c9_rr5;
  wire [15:0] t1_r0_c9_rr6;
  wire [15:0] t1_r0_c9_rr7;
  wire [15:0] t2_r0_c9_rr0;
  wire [15:0] t2_r0_c9_rr1;
  wire [15:0] t2_r0_c9_rr2;
  wire [15:0] t2_r0_c9_rr3;
  wire [15:0] t3_r0_c9_rr0;
  wire [15:0] t3_r0_c9_rr1;
  wire [15:0] t4_r0_c9_rr0;
  wire [15:0] t0_r0_c10_rr0;
  wire [15:0] t0_r0_c10_rr1;
  wire [15:0] t0_r0_c10_rr2;
  wire [15:0] t0_r0_c10_rr3;
  wire [15:0] t0_r0_c10_rr4;
  wire [15:0] t0_r0_c10_rr5;
  wire [15:0] t0_r0_c10_rr6;
  wire [15:0] t0_r0_c10_rr7;
  wire [15:0] t0_r0_c10_rr8;
  wire [15:0] t0_r0_c10_rr9;
  wire [15:0] t0_r0_c10_rr10;
  wire [15:0] t0_r0_c10_rr11;
  wire [15:0] t0_r0_c10_rr12;
  wire [15:0] t0_r0_c10_rr13;
  wire [15:0] t0_r0_c10_rr14;
  wire [15:0] t1_r0_c10_rr0;
  wire [15:0] t1_r0_c10_rr1;
  wire [15:0] t1_r0_c10_rr2;
  wire [15:0] t1_r0_c10_rr3;
  wire [15:0] t1_r0_c10_rr4;
  wire [15:0] t1_r0_c10_rr5;
  wire [15:0] t1_r0_c10_rr6;
  wire [15:0] t1_r0_c10_rr7;
  wire [15:0] t2_r0_c10_rr0;
  wire [15:0] t2_r0_c10_rr1;
  wire [15:0] t2_r0_c10_rr2;
  wire [15:0] t2_r0_c10_rr3;
  wire [15:0] t3_r0_c10_rr0;
  wire [15:0] t3_r0_c10_rr1;
  wire [15:0] t4_r0_c10_rr0;
  wire [15:0] t0_r0_c11_rr0;
  wire [15:0] t0_r0_c11_rr1;
  wire [15:0] t0_r0_c11_rr2;
  wire [15:0] t0_r0_c11_rr3;
  wire [15:0] t0_r0_c11_rr4;
  wire [15:0] t0_r0_c11_rr5;
  wire [15:0] t0_r0_c11_rr6;
  wire [15:0] t0_r0_c11_rr7;
  wire [15:0] t0_r0_c11_rr8;
  wire [15:0] t0_r0_c11_rr9;
  wire [15:0] t0_r0_c11_rr10;
  wire [15:0] t0_r0_c11_rr11;
  wire [15:0] t0_r0_c11_rr12;
  wire [15:0] t0_r0_c11_rr13;
  wire [15:0] t0_r0_c11_rr14;
  wire [15:0] t1_r0_c11_rr0;
  wire [15:0] t1_r0_c11_rr1;
  wire [15:0] t1_r0_c11_rr2;
  wire [15:0] t1_r0_c11_rr3;
  wire [15:0] t1_r0_c11_rr4;
  wire [15:0] t1_r0_c11_rr5;
  wire [15:0] t1_r0_c11_rr6;
  wire [15:0] t1_r0_c11_rr7;
  wire [15:0] t2_r0_c11_rr0;
  wire [15:0] t2_r0_c11_rr1;
  wire [15:0] t2_r0_c11_rr2;
  wire [15:0] t2_r0_c11_rr3;
  wire [15:0] t3_r0_c11_rr0;
  wire [15:0] t3_r0_c11_rr1;
  wire [15:0] t4_r0_c11_rr0;
  wire [15:0] t0_r0_c12_rr0;
  wire [15:0] t0_r0_c12_rr1;
  wire [15:0] t0_r0_c12_rr2;
  wire [15:0] t0_r0_c12_rr3;
  wire [15:0] t0_r0_c12_rr4;
  wire [15:0] t0_r0_c12_rr5;
  wire [15:0] t0_r0_c12_rr6;
  wire [15:0] t0_r0_c12_rr7;
  wire [15:0] t0_r0_c12_rr8;
  wire [15:0] t0_r0_c12_rr9;
  wire [15:0] t0_r0_c12_rr10;
  wire [15:0] t0_r0_c12_rr11;
  wire [15:0] t0_r0_c12_rr12;
  wire [15:0] t0_r0_c12_rr13;
  wire [15:0] t0_r0_c12_rr14;
  wire [15:0] t1_r0_c12_rr0;
  wire [15:0] t1_r0_c12_rr1;
  wire [15:0] t1_r0_c12_rr2;
  wire [15:0] t1_r0_c12_rr3;
  wire [15:0] t1_r0_c12_rr4;
  wire [15:0] t1_r0_c12_rr5;
  wire [15:0] t1_r0_c12_rr6;
  wire [15:0] t1_r0_c12_rr7;
  wire [15:0] t2_r0_c12_rr0;
  wire [15:0] t2_r0_c12_rr1;
  wire [15:0] t2_r0_c12_rr2;
  wire [15:0] t2_r0_c12_rr3;
  wire [15:0] t3_r0_c12_rr0;
  wire [15:0] t3_r0_c12_rr1;
  wire [15:0] t4_r0_c12_rr0;
  wire [15:0] t0_r0_c13_rr0;
  wire [15:0] t0_r0_c13_rr1;
  wire [15:0] t0_r0_c13_rr2;
  wire [15:0] t0_r0_c13_rr3;
  wire [15:0] t0_r0_c13_rr4;
  wire [15:0] t0_r0_c13_rr5;
  wire [15:0] t0_r0_c13_rr6;
  wire [15:0] t0_r0_c13_rr7;
  wire [15:0] t0_r0_c13_rr8;
  wire [15:0] t0_r0_c13_rr9;
  wire [15:0] t0_r0_c13_rr10;
  wire [15:0] t0_r0_c13_rr11;
  wire [15:0] t0_r0_c13_rr12;
  wire [15:0] t0_r0_c13_rr13;
  wire [15:0] t0_r0_c13_rr14;
  wire [15:0] t1_r0_c13_rr0;
  wire [15:0] t1_r0_c13_rr1;
  wire [15:0] t1_r0_c13_rr2;
  wire [15:0] t1_r0_c13_rr3;
  wire [15:0] t1_r0_c13_rr4;
  wire [15:0] t1_r0_c13_rr5;
  wire [15:0] t1_r0_c13_rr6;
  wire [15:0] t1_r0_c13_rr7;
  wire [15:0] t2_r0_c13_rr0;
  wire [15:0] t2_r0_c13_rr1;
  wire [15:0] t2_r0_c13_rr2;
  wire [15:0] t2_r0_c13_rr3;
  wire [15:0] t3_r0_c13_rr0;
  wire [15:0] t3_r0_c13_rr1;
  wire [15:0] t4_r0_c13_rr0;
  wire [15:0] t0_r0_c14_rr0;
  wire [15:0] t0_r0_c14_rr1;
  wire [15:0] t0_r0_c14_rr2;
  wire [15:0] t0_r0_c14_rr3;
  wire [15:0] t0_r0_c14_rr4;
  wire [15:0] t0_r0_c14_rr5;
  wire [15:0] t0_r0_c14_rr6;
  wire [15:0] t0_r0_c14_rr7;
  wire [15:0] t0_r0_c14_rr8;
  wire [15:0] t0_r0_c14_rr9;
  wire [15:0] t0_r0_c14_rr10;
  wire [15:0] t0_r0_c14_rr11;
  wire [15:0] t0_r0_c14_rr12;
  wire [15:0] t0_r0_c14_rr13;
  wire [15:0] t0_r0_c14_rr14;
  wire [15:0] t1_r0_c14_rr0;
  wire [15:0] t1_r0_c14_rr1;
  wire [15:0] t1_r0_c14_rr2;
  wire [15:0] t1_r0_c14_rr3;
  wire [15:0] t1_r0_c14_rr4;
  wire [15:0] t1_r0_c14_rr5;
  wire [15:0] t1_r0_c14_rr6;
  wire [15:0] t1_r0_c14_rr7;
  wire [15:0] t2_r0_c14_rr0;
  wire [15:0] t2_r0_c14_rr1;
  wire [15:0] t2_r0_c14_rr2;
  wire [15:0] t2_r0_c14_rr3;
  wire [15:0] t3_r0_c14_rr0;
  wire [15:0] t3_r0_c14_rr1;
  wire [15:0] t4_r0_c14_rr0;
  wire [15:0] t0_r1_c0_rr0;
  wire [15:0] t0_r1_c0_rr1;
  wire [15:0] t0_r1_c0_rr2;
  wire [15:0] t0_r1_c0_rr3;
  wire [15:0] t0_r1_c0_rr4;
  wire [15:0] t0_r1_c0_rr5;
  wire [15:0] t0_r1_c0_rr6;
  wire [15:0] t0_r1_c0_rr7;
  wire [15:0] t0_r1_c0_rr8;
  wire [15:0] t0_r1_c0_rr9;
  wire [15:0] t0_r1_c0_rr10;
  wire [15:0] t0_r1_c0_rr11;
  wire [15:0] t0_r1_c0_rr12;
  wire [15:0] t0_r1_c0_rr13;
  wire [15:0] t0_r1_c0_rr14;
  wire [15:0] t1_r1_c0_rr0;
  wire [15:0] t1_r1_c0_rr1;
  wire [15:0] t1_r1_c0_rr2;
  wire [15:0] t1_r1_c0_rr3;
  wire [15:0] t1_r1_c0_rr4;
  wire [15:0] t1_r1_c0_rr5;
  wire [15:0] t1_r1_c0_rr6;
  wire [15:0] t1_r1_c0_rr7;
  wire [15:0] t2_r1_c0_rr0;
  wire [15:0] t2_r1_c0_rr1;
  wire [15:0] t2_r1_c0_rr2;
  wire [15:0] t2_r1_c0_rr3;
  wire [15:0] t3_r1_c0_rr0;
  wire [15:0] t3_r1_c0_rr1;
  wire [15:0] t4_r1_c0_rr0;
  wire [15:0] t0_r1_c1_rr0;
  wire [15:0] t0_r1_c1_rr1;
  wire [15:0] t0_r1_c1_rr2;
  wire [15:0] t0_r1_c1_rr3;
  wire [15:0] t0_r1_c1_rr4;
  wire [15:0] t0_r1_c1_rr5;
  wire [15:0] t0_r1_c1_rr6;
  wire [15:0] t0_r1_c1_rr7;
  wire [15:0] t0_r1_c1_rr8;
  wire [15:0] t0_r1_c1_rr9;
  wire [15:0] t0_r1_c1_rr10;
  wire [15:0] t0_r1_c1_rr11;
  wire [15:0] t0_r1_c1_rr12;
  wire [15:0] t0_r1_c1_rr13;
  wire [15:0] t0_r1_c1_rr14;
  wire [15:0] t1_r1_c1_rr0;
  wire [15:0] t1_r1_c1_rr1;
  wire [15:0] t1_r1_c1_rr2;
  wire [15:0] t1_r1_c1_rr3;
  wire [15:0] t1_r1_c1_rr4;
  wire [15:0] t1_r1_c1_rr5;
  wire [15:0] t1_r1_c1_rr6;
  wire [15:0] t1_r1_c1_rr7;
  wire [15:0] t2_r1_c1_rr0;
  wire [15:0] t2_r1_c1_rr1;
  wire [15:0] t2_r1_c1_rr2;
  wire [15:0] t2_r1_c1_rr3;
  wire [15:0] t3_r1_c1_rr0;
  wire [15:0] t3_r1_c1_rr1;
  wire [15:0] t4_r1_c1_rr0;
  wire [15:0] t0_r1_c2_rr0;
  wire [15:0] t0_r1_c2_rr1;
  wire [15:0] t0_r1_c2_rr2;
  wire [15:0] t0_r1_c2_rr3;
  wire [15:0] t0_r1_c2_rr4;
  wire [15:0] t0_r1_c2_rr5;
  wire [15:0] t0_r1_c2_rr6;
  wire [15:0] t0_r1_c2_rr7;
  wire [15:0] t0_r1_c2_rr8;
  wire [15:0] t0_r1_c2_rr9;
  wire [15:0] t0_r1_c2_rr10;
  wire [15:0] t0_r1_c2_rr11;
  wire [15:0] t0_r1_c2_rr12;
  wire [15:0] t0_r1_c2_rr13;
  wire [15:0] t0_r1_c2_rr14;
  wire [15:0] t1_r1_c2_rr0;
  wire [15:0] t1_r1_c2_rr1;
  wire [15:0] t1_r1_c2_rr2;
  wire [15:0] t1_r1_c2_rr3;
  wire [15:0] t1_r1_c2_rr4;
  wire [15:0] t1_r1_c2_rr5;
  wire [15:0] t1_r1_c2_rr6;
  wire [15:0] t1_r1_c2_rr7;
  wire [15:0] t2_r1_c2_rr0;
  wire [15:0] t2_r1_c2_rr1;
  wire [15:0] t2_r1_c2_rr2;
  wire [15:0] t2_r1_c2_rr3;
  wire [15:0] t3_r1_c2_rr0;
  wire [15:0] t3_r1_c2_rr1;
  wire [15:0] t4_r1_c2_rr0;
  wire [15:0] t0_r1_c3_rr0;
  wire [15:0] t0_r1_c3_rr1;
  wire [15:0] t0_r1_c3_rr2;
  wire [15:0] t0_r1_c3_rr3;
  wire [15:0] t0_r1_c3_rr4;
  wire [15:0] t0_r1_c3_rr5;
  wire [15:0] t0_r1_c3_rr6;
  wire [15:0] t0_r1_c3_rr7;
  wire [15:0] t0_r1_c3_rr8;
  wire [15:0] t0_r1_c3_rr9;
  wire [15:0] t0_r1_c3_rr10;
  wire [15:0] t0_r1_c3_rr11;
  wire [15:0] t0_r1_c3_rr12;
  wire [15:0] t0_r1_c3_rr13;
  wire [15:0] t0_r1_c3_rr14;
  wire [15:0] t1_r1_c3_rr0;
  wire [15:0] t1_r1_c3_rr1;
  wire [15:0] t1_r1_c3_rr2;
  wire [15:0] t1_r1_c3_rr3;
  wire [15:0] t1_r1_c3_rr4;
  wire [15:0] t1_r1_c3_rr5;
  wire [15:0] t1_r1_c3_rr6;
  wire [15:0] t1_r1_c3_rr7;
  wire [15:0] t2_r1_c3_rr0;
  wire [15:0] t2_r1_c3_rr1;
  wire [15:0] t2_r1_c3_rr2;
  wire [15:0] t2_r1_c3_rr3;
  wire [15:0] t3_r1_c3_rr0;
  wire [15:0] t3_r1_c3_rr1;
  wire [15:0] t4_r1_c3_rr0;
  wire [15:0] t0_r1_c4_rr0;
  wire [15:0] t0_r1_c4_rr1;
  wire [15:0] t0_r1_c4_rr2;
  wire [15:0] t0_r1_c4_rr3;
  wire [15:0] t0_r1_c4_rr4;
  wire [15:0] t0_r1_c4_rr5;
  wire [15:0] t0_r1_c4_rr6;
  wire [15:0] t0_r1_c4_rr7;
  wire [15:0] t0_r1_c4_rr8;
  wire [15:0] t0_r1_c4_rr9;
  wire [15:0] t0_r1_c4_rr10;
  wire [15:0] t0_r1_c4_rr11;
  wire [15:0] t0_r1_c4_rr12;
  wire [15:0] t0_r1_c4_rr13;
  wire [15:0] t0_r1_c4_rr14;
  wire [15:0] t1_r1_c4_rr0;
  wire [15:0] t1_r1_c4_rr1;
  wire [15:0] t1_r1_c4_rr2;
  wire [15:0] t1_r1_c4_rr3;
  wire [15:0] t1_r1_c4_rr4;
  wire [15:0] t1_r1_c4_rr5;
  wire [15:0] t1_r1_c4_rr6;
  wire [15:0] t1_r1_c4_rr7;
  wire [15:0] t2_r1_c4_rr0;
  wire [15:0] t2_r1_c4_rr1;
  wire [15:0] t2_r1_c4_rr2;
  wire [15:0] t2_r1_c4_rr3;
  wire [15:0] t3_r1_c4_rr0;
  wire [15:0] t3_r1_c4_rr1;
  wire [15:0] t4_r1_c4_rr0;
  wire [15:0] t0_r1_c5_rr0;
  wire [15:0] t0_r1_c5_rr1;
  wire [15:0] t0_r1_c5_rr2;
  wire [15:0] t0_r1_c5_rr3;
  wire [15:0] t0_r1_c5_rr4;
  wire [15:0] t0_r1_c5_rr5;
  wire [15:0] t0_r1_c5_rr6;
  wire [15:0] t0_r1_c5_rr7;
  wire [15:0] t0_r1_c5_rr8;
  wire [15:0] t0_r1_c5_rr9;
  wire [15:0] t0_r1_c5_rr10;
  wire [15:0] t0_r1_c5_rr11;
  wire [15:0] t0_r1_c5_rr12;
  wire [15:0] t0_r1_c5_rr13;
  wire [15:0] t0_r1_c5_rr14;
  wire [15:0] t1_r1_c5_rr0;
  wire [15:0] t1_r1_c5_rr1;
  wire [15:0] t1_r1_c5_rr2;
  wire [15:0] t1_r1_c5_rr3;
  wire [15:0] t1_r1_c5_rr4;
  wire [15:0] t1_r1_c5_rr5;
  wire [15:0] t1_r1_c5_rr6;
  wire [15:0] t1_r1_c5_rr7;
  wire [15:0] t2_r1_c5_rr0;
  wire [15:0] t2_r1_c5_rr1;
  wire [15:0] t2_r1_c5_rr2;
  wire [15:0] t2_r1_c5_rr3;
  wire [15:0] t3_r1_c5_rr0;
  wire [15:0] t3_r1_c5_rr1;
  wire [15:0] t4_r1_c5_rr0;
  wire [15:0] t0_r1_c6_rr0;
  wire [15:0] t0_r1_c6_rr1;
  wire [15:0] t0_r1_c6_rr2;
  wire [15:0] t0_r1_c6_rr3;
  wire [15:0] t0_r1_c6_rr4;
  wire [15:0] t0_r1_c6_rr5;
  wire [15:0] t0_r1_c6_rr6;
  wire [15:0] t0_r1_c6_rr7;
  wire [15:0] t0_r1_c6_rr8;
  wire [15:0] t0_r1_c6_rr9;
  wire [15:0] t0_r1_c6_rr10;
  wire [15:0] t0_r1_c6_rr11;
  wire [15:0] t0_r1_c6_rr12;
  wire [15:0] t0_r1_c6_rr13;
  wire [15:0] t0_r1_c6_rr14;
  wire [15:0] t1_r1_c6_rr0;
  wire [15:0] t1_r1_c6_rr1;
  wire [15:0] t1_r1_c6_rr2;
  wire [15:0] t1_r1_c6_rr3;
  wire [15:0] t1_r1_c6_rr4;
  wire [15:0] t1_r1_c6_rr5;
  wire [15:0] t1_r1_c6_rr6;
  wire [15:0] t1_r1_c6_rr7;
  wire [15:0] t2_r1_c6_rr0;
  wire [15:0] t2_r1_c6_rr1;
  wire [15:0] t2_r1_c6_rr2;
  wire [15:0] t2_r1_c6_rr3;
  wire [15:0] t3_r1_c6_rr0;
  wire [15:0] t3_r1_c6_rr1;
  wire [15:0] t4_r1_c6_rr0;
  wire [15:0] t0_r1_c7_rr0;
  wire [15:0] t0_r1_c7_rr1;
  wire [15:0] t0_r1_c7_rr2;
  wire [15:0] t0_r1_c7_rr3;
  wire [15:0] t0_r1_c7_rr4;
  wire [15:0] t0_r1_c7_rr5;
  wire [15:0] t0_r1_c7_rr6;
  wire [15:0] t0_r1_c7_rr7;
  wire [15:0] t0_r1_c7_rr8;
  wire [15:0] t0_r1_c7_rr9;
  wire [15:0] t0_r1_c7_rr10;
  wire [15:0] t0_r1_c7_rr11;
  wire [15:0] t0_r1_c7_rr12;
  wire [15:0] t0_r1_c7_rr13;
  wire [15:0] t0_r1_c7_rr14;
  wire [15:0] t1_r1_c7_rr0;
  wire [15:0] t1_r1_c7_rr1;
  wire [15:0] t1_r1_c7_rr2;
  wire [15:0] t1_r1_c7_rr3;
  wire [15:0] t1_r1_c7_rr4;
  wire [15:0] t1_r1_c7_rr5;
  wire [15:0] t1_r1_c7_rr6;
  wire [15:0] t1_r1_c7_rr7;
  wire [15:0] t2_r1_c7_rr0;
  wire [15:0] t2_r1_c7_rr1;
  wire [15:0] t2_r1_c7_rr2;
  wire [15:0] t2_r1_c7_rr3;
  wire [15:0] t3_r1_c7_rr0;
  wire [15:0] t3_r1_c7_rr1;
  wire [15:0] t4_r1_c7_rr0;
  wire [15:0] t0_r1_c8_rr0;
  wire [15:0] t0_r1_c8_rr1;
  wire [15:0] t0_r1_c8_rr2;
  wire [15:0] t0_r1_c8_rr3;
  wire [15:0] t0_r1_c8_rr4;
  wire [15:0] t0_r1_c8_rr5;
  wire [15:0] t0_r1_c8_rr6;
  wire [15:0] t0_r1_c8_rr7;
  wire [15:0] t0_r1_c8_rr8;
  wire [15:0] t0_r1_c8_rr9;
  wire [15:0] t0_r1_c8_rr10;
  wire [15:0] t0_r1_c8_rr11;
  wire [15:0] t0_r1_c8_rr12;
  wire [15:0] t0_r1_c8_rr13;
  wire [15:0] t0_r1_c8_rr14;
  wire [15:0] t1_r1_c8_rr0;
  wire [15:0] t1_r1_c8_rr1;
  wire [15:0] t1_r1_c8_rr2;
  wire [15:0] t1_r1_c8_rr3;
  wire [15:0] t1_r1_c8_rr4;
  wire [15:0] t1_r1_c8_rr5;
  wire [15:0] t1_r1_c8_rr6;
  wire [15:0] t1_r1_c8_rr7;
  wire [15:0] t2_r1_c8_rr0;
  wire [15:0] t2_r1_c8_rr1;
  wire [15:0] t2_r1_c8_rr2;
  wire [15:0] t2_r1_c8_rr3;
  wire [15:0] t3_r1_c8_rr0;
  wire [15:0] t3_r1_c8_rr1;
  wire [15:0] t4_r1_c8_rr0;
  wire [15:0] t0_r1_c9_rr0;
  wire [15:0] t0_r1_c9_rr1;
  wire [15:0] t0_r1_c9_rr2;
  wire [15:0] t0_r1_c9_rr3;
  wire [15:0] t0_r1_c9_rr4;
  wire [15:0] t0_r1_c9_rr5;
  wire [15:0] t0_r1_c9_rr6;
  wire [15:0] t0_r1_c9_rr7;
  wire [15:0] t0_r1_c9_rr8;
  wire [15:0] t0_r1_c9_rr9;
  wire [15:0] t0_r1_c9_rr10;
  wire [15:0] t0_r1_c9_rr11;
  wire [15:0] t0_r1_c9_rr12;
  wire [15:0] t0_r1_c9_rr13;
  wire [15:0] t0_r1_c9_rr14;
  wire [15:0] t1_r1_c9_rr0;
  wire [15:0] t1_r1_c9_rr1;
  wire [15:0] t1_r1_c9_rr2;
  wire [15:0] t1_r1_c9_rr3;
  wire [15:0] t1_r1_c9_rr4;
  wire [15:0] t1_r1_c9_rr5;
  wire [15:0] t1_r1_c9_rr6;
  wire [15:0] t1_r1_c9_rr7;
  wire [15:0] t2_r1_c9_rr0;
  wire [15:0] t2_r1_c9_rr1;
  wire [15:0] t2_r1_c9_rr2;
  wire [15:0] t2_r1_c9_rr3;
  wire [15:0] t3_r1_c9_rr0;
  wire [15:0] t3_r1_c9_rr1;
  wire [15:0] t4_r1_c9_rr0;
  wire [15:0] t0_r1_c10_rr0;
  wire [15:0] t0_r1_c10_rr1;
  wire [15:0] t0_r1_c10_rr2;
  wire [15:0] t0_r1_c10_rr3;
  wire [15:0] t0_r1_c10_rr4;
  wire [15:0] t0_r1_c10_rr5;
  wire [15:0] t0_r1_c10_rr6;
  wire [15:0] t0_r1_c10_rr7;
  wire [15:0] t0_r1_c10_rr8;
  wire [15:0] t0_r1_c10_rr9;
  wire [15:0] t0_r1_c10_rr10;
  wire [15:0] t0_r1_c10_rr11;
  wire [15:0] t0_r1_c10_rr12;
  wire [15:0] t0_r1_c10_rr13;
  wire [15:0] t0_r1_c10_rr14;
  wire [15:0] t1_r1_c10_rr0;
  wire [15:0] t1_r1_c10_rr1;
  wire [15:0] t1_r1_c10_rr2;
  wire [15:0] t1_r1_c10_rr3;
  wire [15:0] t1_r1_c10_rr4;
  wire [15:0] t1_r1_c10_rr5;
  wire [15:0] t1_r1_c10_rr6;
  wire [15:0] t1_r1_c10_rr7;
  wire [15:0] t2_r1_c10_rr0;
  wire [15:0] t2_r1_c10_rr1;
  wire [15:0] t2_r1_c10_rr2;
  wire [15:0] t2_r1_c10_rr3;
  wire [15:0] t3_r1_c10_rr0;
  wire [15:0] t3_r1_c10_rr1;
  wire [15:0] t4_r1_c10_rr0;
  wire [15:0] t0_r1_c11_rr0;
  wire [15:0] t0_r1_c11_rr1;
  wire [15:0] t0_r1_c11_rr2;
  wire [15:0] t0_r1_c11_rr3;
  wire [15:0] t0_r1_c11_rr4;
  wire [15:0] t0_r1_c11_rr5;
  wire [15:0] t0_r1_c11_rr6;
  wire [15:0] t0_r1_c11_rr7;
  wire [15:0] t0_r1_c11_rr8;
  wire [15:0] t0_r1_c11_rr9;
  wire [15:0] t0_r1_c11_rr10;
  wire [15:0] t0_r1_c11_rr11;
  wire [15:0] t0_r1_c11_rr12;
  wire [15:0] t0_r1_c11_rr13;
  wire [15:0] t0_r1_c11_rr14;
  wire [15:0] t1_r1_c11_rr0;
  wire [15:0] t1_r1_c11_rr1;
  wire [15:0] t1_r1_c11_rr2;
  wire [15:0] t1_r1_c11_rr3;
  wire [15:0] t1_r1_c11_rr4;
  wire [15:0] t1_r1_c11_rr5;
  wire [15:0] t1_r1_c11_rr6;
  wire [15:0] t1_r1_c11_rr7;
  wire [15:0] t2_r1_c11_rr0;
  wire [15:0] t2_r1_c11_rr1;
  wire [15:0] t2_r1_c11_rr2;
  wire [15:0] t2_r1_c11_rr3;
  wire [15:0] t3_r1_c11_rr0;
  wire [15:0] t3_r1_c11_rr1;
  wire [15:0] t4_r1_c11_rr0;
  wire [15:0] t0_r1_c12_rr0;
  wire [15:0] t0_r1_c12_rr1;
  wire [15:0] t0_r1_c12_rr2;
  wire [15:0] t0_r1_c12_rr3;
  wire [15:0] t0_r1_c12_rr4;
  wire [15:0] t0_r1_c12_rr5;
  wire [15:0] t0_r1_c12_rr6;
  wire [15:0] t0_r1_c12_rr7;
  wire [15:0] t0_r1_c12_rr8;
  wire [15:0] t0_r1_c12_rr9;
  wire [15:0] t0_r1_c12_rr10;
  wire [15:0] t0_r1_c12_rr11;
  wire [15:0] t0_r1_c12_rr12;
  wire [15:0] t0_r1_c12_rr13;
  wire [15:0] t0_r1_c12_rr14;
  wire [15:0] t1_r1_c12_rr0;
  wire [15:0] t1_r1_c12_rr1;
  wire [15:0] t1_r1_c12_rr2;
  wire [15:0] t1_r1_c12_rr3;
  wire [15:0] t1_r1_c12_rr4;
  wire [15:0] t1_r1_c12_rr5;
  wire [15:0] t1_r1_c12_rr6;
  wire [15:0] t1_r1_c12_rr7;
  wire [15:0] t2_r1_c12_rr0;
  wire [15:0] t2_r1_c12_rr1;
  wire [15:0] t2_r1_c12_rr2;
  wire [15:0] t2_r1_c12_rr3;
  wire [15:0] t3_r1_c12_rr0;
  wire [15:0] t3_r1_c12_rr1;
  wire [15:0] t4_r1_c12_rr0;
  wire [15:0] t0_r1_c13_rr0;
  wire [15:0] t0_r1_c13_rr1;
  wire [15:0] t0_r1_c13_rr2;
  wire [15:0] t0_r1_c13_rr3;
  wire [15:0] t0_r1_c13_rr4;
  wire [15:0] t0_r1_c13_rr5;
  wire [15:0] t0_r1_c13_rr6;
  wire [15:0] t0_r1_c13_rr7;
  wire [15:0] t0_r1_c13_rr8;
  wire [15:0] t0_r1_c13_rr9;
  wire [15:0] t0_r1_c13_rr10;
  wire [15:0] t0_r1_c13_rr11;
  wire [15:0] t0_r1_c13_rr12;
  wire [15:0] t0_r1_c13_rr13;
  wire [15:0] t0_r1_c13_rr14;
  wire [15:0] t1_r1_c13_rr0;
  wire [15:0] t1_r1_c13_rr1;
  wire [15:0] t1_r1_c13_rr2;
  wire [15:0] t1_r1_c13_rr3;
  wire [15:0] t1_r1_c13_rr4;
  wire [15:0] t1_r1_c13_rr5;
  wire [15:0] t1_r1_c13_rr6;
  wire [15:0] t1_r1_c13_rr7;
  wire [15:0] t2_r1_c13_rr0;
  wire [15:0] t2_r1_c13_rr1;
  wire [15:0] t2_r1_c13_rr2;
  wire [15:0] t2_r1_c13_rr3;
  wire [15:0] t3_r1_c13_rr0;
  wire [15:0] t3_r1_c13_rr1;
  wire [15:0] t4_r1_c13_rr0;
  wire [15:0] t0_r1_c14_rr0;
  wire [15:0] t0_r1_c14_rr1;
  wire [15:0] t0_r1_c14_rr2;
  wire [15:0] t0_r1_c14_rr3;
  wire [15:0] t0_r1_c14_rr4;
  wire [15:0] t0_r1_c14_rr5;
  wire [15:0] t0_r1_c14_rr6;
  wire [15:0] t0_r1_c14_rr7;
  wire [15:0] t0_r1_c14_rr8;
  wire [15:0] t0_r1_c14_rr9;
  wire [15:0] t0_r1_c14_rr10;
  wire [15:0] t0_r1_c14_rr11;
  wire [15:0] t0_r1_c14_rr12;
  wire [15:0] t0_r1_c14_rr13;
  wire [15:0] t0_r1_c14_rr14;
  wire [15:0] t1_r1_c14_rr0;
  wire [15:0] t1_r1_c14_rr1;
  wire [15:0] t1_r1_c14_rr2;
  wire [15:0] t1_r1_c14_rr3;
  wire [15:0] t1_r1_c14_rr4;
  wire [15:0] t1_r1_c14_rr5;
  wire [15:0] t1_r1_c14_rr6;
  wire [15:0] t1_r1_c14_rr7;
  wire [15:0] t2_r1_c14_rr0;
  wire [15:0] t2_r1_c14_rr1;
  wire [15:0] t2_r1_c14_rr2;
  wire [15:0] t2_r1_c14_rr3;
  wire [15:0] t3_r1_c14_rr0;
  wire [15:0] t3_r1_c14_rr1;
  wire [15:0] t4_r1_c14_rr0;
  wire [15:0] t0_r2_c0_rr0;
  wire [15:0] t0_r2_c0_rr1;
  wire [15:0] t0_r2_c0_rr2;
  wire [15:0] t0_r2_c0_rr3;
  wire [15:0] t0_r2_c0_rr4;
  wire [15:0] t0_r2_c0_rr5;
  wire [15:0] t0_r2_c0_rr6;
  wire [15:0] t0_r2_c0_rr7;
  wire [15:0] t0_r2_c0_rr8;
  wire [15:0] t0_r2_c0_rr9;
  wire [15:0] t0_r2_c0_rr10;
  wire [15:0] t0_r2_c0_rr11;
  wire [15:0] t0_r2_c0_rr12;
  wire [15:0] t0_r2_c0_rr13;
  wire [15:0] t0_r2_c0_rr14;
  wire [15:0] t1_r2_c0_rr0;
  wire [15:0] t1_r2_c0_rr1;
  wire [15:0] t1_r2_c0_rr2;
  wire [15:0] t1_r2_c0_rr3;
  wire [15:0] t1_r2_c0_rr4;
  wire [15:0] t1_r2_c0_rr5;
  wire [15:0] t1_r2_c0_rr6;
  wire [15:0] t1_r2_c0_rr7;
  wire [15:0] t2_r2_c0_rr0;
  wire [15:0] t2_r2_c0_rr1;
  wire [15:0] t2_r2_c0_rr2;
  wire [15:0] t2_r2_c0_rr3;
  wire [15:0] t3_r2_c0_rr0;
  wire [15:0] t3_r2_c0_rr1;
  wire [15:0] t4_r2_c0_rr0;
  wire [15:0] t0_r2_c1_rr0;
  wire [15:0] t0_r2_c1_rr1;
  wire [15:0] t0_r2_c1_rr2;
  wire [15:0] t0_r2_c1_rr3;
  wire [15:0] t0_r2_c1_rr4;
  wire [15:0] t0_r2_c1_rr5;
  wire [15:0] t0_r2_c1_rr6;
  wire [15:0] t0_r2_c1_rr7;
  wire [15:0] t0_r2_c1_rr8;
  wire [15:0] t0_r2_c1_rr9;
  wire [15:0] t0_r2_c1_rr10;
  wire [15:0] t0_r2_c1_rr11;
  wire [15:0] t0_r2_c1_rr12;
  wire [15:0] t0_r2_c1_rr13;
  wire [15:0] t0_r2_c1_rr14;
  wire [15:0] t1_r2_c1_rr0;
  wire [15:0] t1_r2_c1_rr1;
  wire [15:0] t1_r2_c1_rr2;
  wire [15:0] t1_r2_c1_rr3;
  wire [15:0] t1_r2_c1_rr4;
  wire [15:0] t1_r2_c1_rr5;
  wire [15:0] t1_r2_c1_rr6;
  wire [15:0] t1_r2_c1_rr7;
  wire [15:0] t2_r2_c1_rr0;
  wire [15:0] t2_r2_c1_rr1;
  wire [15:0] t2_r2_c1_rr2;
  wire [15:0] t2_r2_c1_rr3;
  wire [15:0] t3_r2_c1_rr0;
  wire [15:0] t3_r2_c1_rr1;
  wire [15:0] t4_r2_c1_rr0;
  wire [15:0] t0_r2_c2_rr0;
  wire [15:0] t0_r2_c2_rr1;
  wire [15:0] t0_r2_c2_rr2;
  wire [15:0] t0_r2_c2_rr3;
  wire [15:0] t0_r2_c2_rr4;
  wire [15:0] t0_r2_c2_rr5;
  wire [15:0] t0_r2_c2_rr6;
  wire [15:0] t0_r2_c2_rr7;
  wire [15:0] t0_r2_c2_rr8;
  wire [15:0] t0_r2_c2_rr9;
  wire [15:0] t0_r2_c2_rr10;
  wire [15:0] t0_r2_c2_rr11;
  wire [15:0] t0_r2_c2_rr12;
  wire [15:0] t0_r2_c2_rr13;
  wire [15:0] t0_r2_c2_rr14;
  wire [15:0] t1_r2_c2_rr0;
  wire [15:0] t1_r2_c2_rr1;
  wire [15:0] t1_r2_c2_rr2;
  wire [15:0] t1_r2_c2_rr3;
  wire [15:0] t1_r2_c2_rr4;
  wire [15:0] t1_r2_c2_rr5;
  wire [15:0] t1_r2_c2_rr6;
  wire [15:0] t1_r2_c2_rr7;
  wire [15:0] t2_r2_c2_rr0;
  wire [15:0] t2_r2_c2_rr1;
  wire [15:0] t2_r2_c2_rr2;
  wire [15:0] t2_r2_c2_rr3;
  wire [15:0] t3_r2_c2_rr0;
  wire [15:0] t3_r2_c2_rr1;
  wire [15:0] t4_r2_c2_rr0;
  wire [15:0] t0_r2_c3_rr0;
  wire [15:0] t0_r2_c3_rr1;
  wire [15:0] t0_r2_c3_rr2;
  wire [15:0] t0_r2_c3_rr3;
  wire [15:0] t0_r2_c3_rr4;
  wire [15:0] t0_r2_c3_rr5;
  wire [15:0] t0_r2_c3_rr6;
  wire [15:0] t0_r2_c3_rr7;
  wire [15:0] t0_r2_c3_rr8;
  wire [15:0] t0_r2_c3_rr9;
  wire [15:0] t0_r2_c3_rr10;
  wire [15:0] t0_r2_c3_rr11;
  wire [15:0] t0_r2_c3_rr12;
  wire [15:0] t0_r2_c3_rr13;
  wire [15:0] t0_r2_c3_rr14;
  wire [15:0] t1_r2_c3_rr0;
  wire [15:0] t1_r2_c3_rr1;
  wire [15:0] t1_r2_c3_rr2;
  wire [15:0] t1_r2_c3_rr3;
  wire [15:0] t1_r2_c3_rr4;
  wire [15:0] t1_r2_c3_rr5;
  wire [15:0] t1_r2_c3_rr6;
  wire [15:0] t1_r2_c3_rr7;
  wire [15:0] t2_r2_c3_rr0;
  wire [15:0] t2_r2_c3_rr1;
  wire [15:0] t2_r2_c3_rr2;
  wire [15:0] t2_r2_c3_rr3;
  wire [15:0] t3_r2_c3_rr0;
  wire [15:0] t3_r2_c3_rr1;
  wire [15:0] t4_r2_c3_rr0;
  wire [15:0] t0_r2_c4_rr0;
  wire [15:0] t0_r2_c4_rr1;
  wire [15:0] t0_r2_c4_rr2;
  wire [15:0] t0_r2_c4_rr3;
  wire [15:0] t0_r2_c4_rr4;
  wire [15:0] t0_r2_c4_rr5;
  wire [15:0] t0_r2_c4_rr6;
  wire [15:0] t0_r2_c4_rr7;
  wire [15:0] t0_r2_c4_rr8;
  wire [15:0] t0_r2_c4_rr9;
  wire [15:0] t0_r2_c4_rr10;
  wire [15:0] t0_r2_c4_rr11;
  wire [15:0] t0_r2_c4_rr12;
  wire [15:0] t0_r2_c4_rr13;
  wire [15:0] t0_r2_c4_rr14;
  wire [15:0] t1_r2_c4_rr0;
  wire [15:0] t1_r2_c4_rr1;
  wire [15:0] t1_r2_c4_rr2;
  wire [15:0] t1_r2_c4_rr3;
  wire [15:0] t1_r2_c4_rr4;
  wire [15:0] t1_r2_c4_rr5;
  wire [15:0] t1_r2_c4_rr6;
  wire [15:0] t1_r2_c4_rr7;
  wire [15:0] t2_r2_c4_rr0;
  wire [15:0] t2_r2_c4_rr1;
  wire [15:0] t2_r2_c4_rr2;
  wire [15:0] t2_r2_c4_rr3;
  wire [15:0] t3_r2_c4_rr0;
  wire [15:0] t3_r2_c4_rr1;
  wire [15:0] t4_r2_c4_rr0;
  wire [15:0] t0_r2_c5_rr0;
  wire [15:0] t0_r2_c5_rr1;
  wire [15:0] t0_r2_c5_rr2;
  wire [15:0] t0_r2_c5_rr3;
  wire [15:0] t0_r2_c5_rr4;
  wire [15:0] t0_r2_c5_rr5;
  wire [15:0] t0_r2_c5_rr6;
  wire [15:0] t0_r2_c5_rr7;
  wire [15:0] t0_r2_c5_rr8;
  wire [15:0] t0_r2_c5_rr9;
  wire [15:0] t0_r2_c5_rr10;
  wire [15:0] t0_r2_c5_rr11;
  wire [15:0] t0_r2_c5_rr12;
  wire [15:0] t0_r2_c5_rr13;
  wire [15:0] t0_r2_c5_rr14;
  wire [15:0] t1_r2_c5_rr0;
  wire [15:0] t1_r2_c5_rr1;
  wire [15:0] t1_r2_c5_rr2;
  wire [15:0] t1_r2_c5_rr3;
  wire [15:0] t1_r2_c5_rr4;
  wire [15:0] t1_r2_c5_rr5;
  wire [15:0] t1_r2_c5_rr6;
  wire [15:0] t1_r2_c5_rr7;
  wire [15:0] t2_r2_c5_rr0;
  wire [15:0] t2_r2_c5_rr1;
  wire [15:0] t2_r2_c5_rr2;
  wire [15:0] t2_r2_c5_rr3;
  wire [15:0] t3_r2_c5_rr0;
  wire [15:0] t3_r2_c5_rr1;
  wire [15:0] t4_r2_c5_rr0;
  wire [15:0] t0_r2_c6_rr0;
  wire [15:0] t0_r2_c6_rr1;
  wire [15:0] t0_r2_c6_rr2;
  wire [15:0] t0_r2_c6_rr3;
  wire [15:0] t0_r2_c6_rr4;
  wire [15:0] t0_r2_c6_rr5;
  wire [15:0] t0_r2_c6_rr6;
  wire [15:0] t0_r2_c6_rr7;
  wire [15:0] t0_r2_c6_rr8;
  wire [15:0] t0_r2_c6_rr9;
  wire [15:0] t0_r2_c6_rr10;
  wire [15:0] t0_r2_c6_rr11;
  wire [15:0] t0_r2_c6_rr12;
  wire [15:0] t0_r2_c6_rr13;
  wire [15:0] t0_r2_c6_rr14;
  wire [15:0] t1_r2_c6_rr0;
  wire [15:0] t1_r2_c6_rr1;
  wire [15:0] t1_r2_c6_rr2;
  wire [15:0] t1_r2_c6_rr3;
  wire [15:0] t1_r2_c6_rr4;
  wire [15:0] t1_r2_c6_rr5;
  wire [15:0] t1_r2_c6_rr6;
  wire [15:0] t1_r2_c6_rr7;
  wire [15:0] t2_r2_c6_rr0;
  wire [15:0] t2_r2_c6_rr1;
  wire [15:0] t2_r2_c6_rr2;
  wire [15:0] t2_r2_c6_rr3;
  wire [15:0] t3_r2_c6_rr0;
  wire [15:0] t3_r2_c6_rr1;
  wire [15:0] t4_r2_c6_rr0;
  wire [15:0] t0_r2_c7_rr0;
  wire [15:0] t0_r2_c7_rr1;
  wire [15:0] t0_r2_c7_rr2;
  wire [15:0] t0_r2_c7_rr3;
  wire [15:0] t0_r2_c7_rr4;
  wire [15:0] t0_r2_c7_rr5;
  wire [15:0] t0_r2_c7_rr6;
  wire [15:0] t0_r2_c7_rr7;
  wire [15:0] t0_r2_c7_rr8;
  wire [15:0] t0_r2_c7_rr9;
  wire [15:0] t0_r2_c7_rr10;
  wire [15:0] t0_r2_c7_rr11;
  wire [15:0] t0_r2_c7_rr12;
  wire [15:0] t0_r2_c7_rr13;
  wire [15:0] t0_r2_c7_rr14;
  wire [15:0] t1_r2_c7_rr0;
  wire [15:0] t1_r2_c7_rr1;
  wire [15:0] t1_r2_c7_rr2;
  wire [15:0] t1_r2_c7_rr3;
  wire [15:0] t1_r2_c7_rr4;
  wire [15:0] t1_r2_c7_rr5;
  wire [15:0] t1_r2_c7_rr6;
  wire [15:0] t1_r2_c7_rr7;
  wire [15:0] t2_r2_c7_rr0;
  wire [15:0] t2_r2_c7_rr1;
  wire [15:0] t2_r2_c7_rr2;
  wire [15:0] t2_r2_c7_rr3;
  wire [15:0] t3_r2_c7_rr0;
  wire [15:0] t3_r2_c7_rr1;
  wire [15:0] t4_r2_c7_rr0;
  wire [15:0] t0_r2_c8_rr0;
  wire [15:0] t0_r2_c8_rr1;
  wire [15:0] t0_r2_c8_rr2;
  wire [15:0] t0_r2_c8_rr3;
  wire [15:0] t0_r2_c8_rr4;
  wire [15:0] t0_r2_c8_rr5;
  wire [15:0] t0_r2_c8_rr6;
  wire [15:0] t0_r2_c8_rr7;
  wire [15:0] t0_r2_c8_rr8;
  wire [15:0] t0_r2_c8_rr9;
  wire [15:0] t0_r2_c8_rr10;
  wire [15:0] t0_r2_c8_rr11;
  wire [15:0] t0_r2_c8_rr12;
  wire [15:0] t0_r2_c8_rr13;
  wire [15:0] t0_r2_c8_rr14;
  wire [15:0] t1_r2_c8_rr0;
  wire [15:0] t1_r2_c8_rr1;
  wire [15:0] t1_r2_c8_rr2;
  wire [15:0] t1_r2_c8_rr3;
  wire [15:0] t1_r2_c8_rr4;
  wire [15:0] t1_r2_c8_rr5;
  wire [15:0] t1_r2_c8_rr6;
  wire [15:0] t1_r2_c8_rr7;
  wire [15:0] t2_r2_c8_rr0;
  wire [15:0] t2_r2_c8_rr1;
  wire [15:0] t2_r2_c8_rr2;
  wire [15:0] t2_r2_c8_rr3;
  wire [15:0] t3_r2_c8_rr0;
  wire [15:0] t3_r2_c8_rr1;
  wire [15:0] t4_r2_c8_rr0;
  wire [15:0] t0_r2_c9_rr0;
  wire [15:0] t0_r2_c9_rr1;
  wire [15:0] t0_r2_c9_rr2;
  wire [15:0] t0_r2_c9_rr3;
  wire [15:0] t0_r2_c9_rr4;
  wire [15:0] t0_r2_c9_rr5;
  wire [15:0] t0_r2_c9_rr6;
  wire [15:0] t0_r2_c9_rr7;
  wire [15:0] t0_r2_c9_rr8;
  wire [15:0] t0_r2_c9_rr9;
  wire [15:0] t0_r2_c9_rr10;
  wire [15:0] t0_r2_c9_rr11;
  wire [15:0] t0_r2_c9_rr12;
  wire [15:0] t0_r2_c9_rr13;
  wire [15:0] t0_r2_c9_rr14;
  wire [15:0] t1_r2_c9_rr0;
  wire [15:0] t1_r2_c9_rr1;
  wire [15:0] t1_r2_c9_rr2;
  wire [15:0] t1_r2_c9_rr3;
  wire [15:0] t1_r2_c9_rr4;
  wire [15:0] t1_r2_c9_rr5;
  wire [15:0] t1_r2_c9_rr6;
  wire [15:0] t1_r2_c9_rr7;
  wire [15:0] t2_r2_c9_rr0;
  wire [15:0] t2_r2_c9_rr1;
  wire [15:0] t2_r2_c9_rr2;
  wire [15:0] t2_r2_c9_rr3;
  wire [15:0] t3_r2_c9_rr0;
  wire [15:0] t3_r2_c9_rr1;
  wire [15:0] t4_r2_c9_rr0;
  wire [15:0] t0_r2_c10_rr0;
  wire [15:0] t0_r2_c10_rr1;
  wire [15:0] t0_r2_c10_rr2;
  wire [15:0] t0_r2_c10_rr3;
  wire [15:0] t0_r2_c10_rr4;
  wire [15:0] t0_r2_c10_rr5;
  wire [15:0] t0_r2_c10_rr6;
  wire [15:0] t0_r2_c10_rr7;
  wire [15:0] t0_r2_c10_rr8;
  wire [15:0] t0_r2_c10_rr9;
  wire [15:0] t0_r2_c10_rr10;
  wire [15:0] t0_r2_c10_rr11;
  wire [15:0] t0_r2_c10_rr12;
  wire [15:0] t0_r2_c10_rr13;
  wire [15:0] t0_r2_c10_rr14;
  wire [15:0] t1_r2_c10_rr0;
  wire [15:0] t1_r2_c10_rr1;
  wire [15:0] t1_r2_c10_rr2;
  wire [15:0] t1_r2_c10_rr3;
  wire [15:0] t1_r2_c10_rr4;
  wire [15:0] t1_r2_c10_rr5;
  wire [15:0] t1_r2_c10_rr6;
  wire [15:0] t1_r2_c10_rr7;
  wire [15:0] t2_r2_c10_rr0;
  wire [15:0] t2_r2_c10_rr1;
  wire [15:0] t2_r2_c10_rr2;
  wire [15:0] t2_r2_c10_rr3;
  wire [15:0] t3_r2_c10_rr0;
  wire [15:0] t3_r2_c10_rr1;
  wire [15:0] t4_r2_c10_rr0;
  wire [15:0] t0_r2_c11_rr0;
  wire [15:0] t0_r2_c11_rr1;
  wire [15:0] t0_r2_c11_rr2;
  wire [15:0] t0_r2_c11_rr3;
  wire [15:0] t0_r2_c11_rr4;
  wire [15:0] t0_r2_c11_rr5;
  wire [15:0] t0_r2_c11_rr6;
  wire [15:0] t0_r2_c11_rr7;
  wire [15:0] t0_r2_c11_rr8;
  wire [15:0] t0_r2_c11_rr9;
  wire [15:0] t0_r2_c11_rr10;
  wire [15:0] t0_r2_c11_rr11;
  wire [15:0] t0_r2_c11_rr12;
  wire [15:0] t0_r2_c11_rr13;
  wire [15:0] t0_r2_c11_rr14;
  wire [15:0] t1_r2_c11_rr0;
  wire [15:0] t1_r2_c11_rr1;
  wire [15:0] t1_r2_c11_rr2;
  wire [15:0] t1_r2_c11_rr3;
  wire [15:0] t1_r2_c11_rr4;
  wire [15:0] t1_r2_c11_rr5;
  wire [15:0] t1_r2_c11_rr6;
  wire [15:0] t1_r2_c11_rr7;
  wire [15:0] t2_r2_c11_rr0;
  wire [15:0] t2_r2_c11_rr1;
  wire [15:0] t2_r2_c11_rr2;
  wire [15:0] t2_r2_c11_rr3;
  wire [15:0] t3_r2_c11_rr0;
  wire [15:0] t3_r2_c11_rr1;
  wire [15:0] t4_r2_c11_rr0;
  wire [15:0] t0_r2_c12_rr0;
  wire [15:0] t0_r2_c12_rr1;
  wire [15:0] t0_r2_c12_rr2;
  wire [15:0] t0_r2_c12_rr3;
  wire [15:0] t0_r2_c12_rr4;
  wire [15:0] t0_r2_c12_rr5;
  wire [15:0] t0_r2_c12_rr6;
  wire [15:0] t0_r2_c12_rr7;
  wire [15:0] t0_r2_c12_rr8;
  wire [15:0] t0_r2_c12_rr9;
  wire [15:0] t0_r2_c12_rr10;
  wire [15:0] t0_r2_c12_rr11;
  wire [15:0] t0_r2_c12_rr12;
  wire [15:0] t0_r2_c12_rr13;
  wire [15:0] t0_r2_c12_rr14;
  wire [15:0] t1_r2_c12_rr0;
  wire [15:0] t1_r2_c12_rr1;
  wire [15:0] t1_r2_c12_rr2;
  wire [15:0] t1_r2_c12_rr3;
  wire [15:0] t1_r2_c12_rr4;
  wire [15:0] t1_r2_c12_rr5;
  wire [15:0] t1_r2_c12_rr6;
  wire [15:0] t1_r2_c12_rr7;
  wire [15:0] t2_r2_c12_rr0;
  wire [15:0] t2_r2_c12_rr1;
  wire [15:0] t2_r2_c12_rr2;
  wire [15:0] t2_r2_c12_rr3;
  wire [15:0] t3_r2_c12_rr0;
  wire [15:0] t3_r2_c12_rr1;
  wire [15:0] t4_r2_c12_rr0;
  wire [15:0] t0_r2_c13_rr0;
  wire [15:0] t0_r2_c13_rr1;
  wire [15:0] t0_r2_c13_rr2;
  wire [15:0] t0_r2_c13_rr3;
  wire [15:0] t0_r2_c13_rr4;
  wire [15:0] t0_r2_c13_rr5;
  wire [15:0] t0_r2_c13_rr6;
  wire [15:0] t0_r2_c13_rr7;
  wire [15:0] t0_r2_c13_rr8;
  wire [15:0] t0_r2_c13_rr9;
  wire [15:0] t0_r2_c13_rr10;
  wire [15:0] t0_r2_c13_rr11;
  wire [15:0] t0_r2_c13_rr12;
  wire [15:0] t0_r2_c13_rr13;
  wire [15:0] t0_r2_c13_rr14;
  wire [15:0] t1_r2_c13_rr0;
  wire [15:0] t1_r2_c13_rr1;
  wire [15:0] t1_r2_c13_rr2;
  wire [15:0] t1_r2_c13_rr3;
  wire [15:0] t1_r2_c13_rr4;
  wire [15:0] t1_r2_c13_rr5;
  wire [15:0] t1_r2_c13_rr6;
  wire [15:0] t1_r2_c13_rr7;
  wire [15:0] t2_r2_c13_rr0;
  wire [15:0] t2_r2_c13_rr1;
  wire [15:0] t2_r2_c13_rr2;
  wire [15:0] t2_r2_c13_rr3;
  wire [15:0] t3_r2_c13_rr0;
  wire [15:0] t3_r2_c13_rr1;
  wire [15:0] t4_r2_c13_rr0;
  wire [15:0] t0_r2_c14_rr0;
  wire [15:0] t0_r2_c14_rr1;
  wire [15:0] t0_r2_c14_rr2;
  wire [15:0] t0_r2_c14_rr3;
  wire [15:0] t0_r2_c14_rr4;
  wire [15:0] t0_r2_c14_rr5;
  wire [15:0] t0_r2_c14_rr6;
  wire [15:0] t0_r2_c14_rr7;
  wire [15:0] t0_r2_c14_rr8;
  wire [15:0] t0_r2_c14_rr9;
  wire [15:0] t0_r2_c14_rr10;
  wire [15:0] t0_r2_c14_rr11;
  wire [15:0] t0_r2_c14_rr12;
  wire [15:0] t0_r2_c14_rr13;
  wire [15:0] t0_r2_c14_rr14;
  wire [15:0] t1_r2_c14_rr0;
  wire [15:0] t1_r2_c14_rr1;
  wire [15:0] t1_r2_c14_rr2;
  wire [15:0] t1_r2_c14_rr3;
  wire [15:0] t1_r2_c14_rr4;
  wire [15:0] t1_r2_c14_rr5;
  wire [15:0] t1_r2_c14_rr6;
  wire [15:0] t1_r2_c14_rr7;
  wire [15:0] t2_r2_c14_rr0;
  wire [15:0] t2_r2_c14_rr1;
  wire [15:0] t2_r2_c14_rr2;
  wire [15:0] t2_r2_c14_rr3;
  wire [15:0] t3_r2_c14_rr0;
  wire [15:0] t3_r2_c14_rr1;
  wire [15:0] t4_r2_c14_rr0;
  wire [15:0] t0_r3_c0_rr0;
  wire [15:0] t0_r3_c0_rr1;
  wire [15:0] t0_r3_c0_rr2;
  wire [15:0] t0_r3_c0_rr3;
  wire [15:0] t0_r3_c0_rr4;
  wire [15:0] t0_r3_c0_rr5;
  wire [15:0] t0_r3_c0_rr6;
  wire [15:0] t0_r3_c0_rr7;
  wire [15:0] t0_r3_c0_rr8;
  wire [15:0] t0_r3_c0_rr9;
  wire [15:0] t0_r3_c0_rr10;
  wire [15:0] t0_r3_c0_rr11;
  wire [15:0] t0_r3_c0_rr12;
  wire [15:0] t0_r3_c0_rr13;
  wire [15:0] t0_r3_c0_rr14;
  wire [15:0] t1_r3_c0_rr0;
  wire [15:0] t1_r3_c0_rr1;
  wire [15:0] t1_r3_c0_rr2;
  wire [15:0] t1_r3_c0_rr3;
  wire [15:0] t1_r3_c0_rr4;
  wire [15:0] t1_r3_c0_rr5;
  wire [15:0] t1_r3_c0_rr6;
  wire [15:0] t1_r3_c0_rr7;
  wire [15:0] t2_r3_c0_rr0;
  wire [15:0] t2_r3_c0_rr1;
  wire [15:0] t2_r3_c0_rr2;
  wire [15:0] t2_r3_c0_rr3;
  wire [15:0] t3_r3_c0_rr0;
  wire [15:0] t3_r3_c0_rr1;
  wire [15:0] t4_r3_c0_rr0;
  wire [15:0] t0_r3_c1_rr0;
  wire [15:0] t0_r3_c1_rr1;
  wire [15:0] t0_r3_c1_rr2;
  wire [15:0] t0_r3_c1_rr3;
  wire [15:0] t0_r3_c1_rr4;
  wire [15:0] t0_r3_c1_rr5;
  wire [15:0] t0_r3_c1_rr6;
  wire [15:0] t0_r3_c1_rr7;
  wire [15:0] t0_r3_c1_rr8;
  wire [15:0] t0_r3_c1_rr9;
  wire [15:0] t0_r3_c1_rr10;
  wire [15:0] t0_r3_c1_rr11;
  wire [15:0] t0_r3_c1_rr12;
  wire [15:0] t0_r3_c1_rr13;
  wire [15:0] t0_r3_c1_rr14;
  wire [15:0] t1_r3_c1_rr0;
  wire [15:0] t1_r3_c1_rr1;
  wire [15:0] t1_r3_c1_rr2;
  wire [15:0] t1_r3_c1_rr3;
  wire [15:0] t1_r3_c1_rr4;
  wire [15:0] t1_r3_c1_rr5;
  wire [15:0] t1_r3_c1_rr6;
  wire [15:0] t1_r3_c1_rr7;
  wire [15:0] t2_r3_c1_rr0;
  wire [15:0] t2_r3_c1_rr1;
  wire [15:0] t2_r3_c1_rr2;
  wire [15:0] t2_r3_c1_rr3;
  wire [15:0] t3_r3_c1_rr0;
  wire [15:0] t3_r3_c1_rr1;
  wire [15:0] t4_r3_c1_rr0;
  wire [15:0] t0_r3_c2_rr0;
  wire [15:0] t0_r3_c2_rr1;
  wire [15:0] t0_r3_c2_rr2;
  wire [15:0] t0_r3_c2_rr3;
  wire [15:0] t0_r3_c2_rr4;
  wire [15:0] t0_r3_c2_rr5;
  wire [15:0] t0_r3_c2_rr6;
  wire [15:0] t0_r3_c2_rr7;
  wire [15:0] t0_r3_c2_rr8;
  wire [15:0] t0_r3_c2_rr9;
  wire [15:0] t0_r3_c2_rr10;
  wire [15:0] t0_r3_c2_rr11;
  wire [15:0] t0_r3_c2_rr12;
  wire [15:0] t0_r3_c2_rr13;
  wire [15:0] t0_r3_c2_rr14;
  wire [15:0] t1_r3_c2_rr0;
  wire [15:0] t1_r3_c2_rr1;
  wire [15:0] t1_r3_c2_rr2;
  wire [15:0] t1_r3_c2_rr3;
  wire [15:0] t1_r3_c2_rr4;
  wire [15:0] t1_r3_c2_rr5;
  wire [15:0] t1_r3_c2_rr6;
  wire [15:0] t1_r3_c2_rr7;
  wire [15:0] t2_r3_c2_rr0;
  wire [15:0] t2_r3_c2_rr1;
  wire [15:0] t2_r3_c2_rr2;
  wire [15:0] t2_r3_c2_rr3;
  wire [15:0] t3_r3_c2_rr0;
  wire [15:0] t3_r3_c2_rr1;
  wire [15:0] t4_r3_c2_rr0;
  wire [15:0] t0_r3_c3_rr0;
  wire [15:0] t0_r3_c3_rr1;
  wire [15:0] t0_r3_c3_rr2;
  wire [15:0] t0_r3_c3_rr3;
  wire [15:0] t0_r3_c3_rr4;
  wire [15:0] t0_r3_c3_rr5;
  wire [15:0] t0_r3_c3_rr6;
  wire [15:0] t0_r3_c3_rr7;
  wire [15:0] t0_r3_c3_rr8;
  wire [15:0] t0_r3_c3_rr9;
  wire [15:0] t0_r3_c3_rr10;
  wire [15:0] t0_r3_c3_rr11;
  wire [15:0] t0_r3_c3_rr12;
  wire [15:0] t0_r3_c3_rr13;
  wire [15:0] t0_r3_c3_rr14;
  wire [15:0] t1_r3_c3_rr0;
  wire [15:0] t1_r3_c3_rr1;
  wire [15:0] t1_r3_c3_rr2;
  wire [15:0] t1_r3_c3_rr3;
  wire [15:0] t1_r3_c3_rr4;
  wire [15:0] t1_r3_c3_rr5;
  wire [15:0] t1_r3_c3_rr6;
  wire [15:0] t1_r3_c3_rr7;
  wire [15:0] t2_r3_c3_rr0;
  wire [15:0] t2_r3_c3_rr1;
  wire [15:0] t2_r3_c3_rr2;
  wire [15:0] t2_r3_c3_rr3;
  wire [15:0] t3_r3_c3_rr0;
  wire [15:0] t3_r3_c3_rr1;
  wire [15:0] t4_r3_c3_rr0;
  wire [15:0] t0_r3_c4_rr0;
  wire [15:0] t0_r3_c4_rr1;
  wire [15:0] t0_r3_c4_rr2;
  wire [15:0] t0_r3_c4_rr3;
  wire [15:0] t0_r3_c4_rr4;
  wire [15:0] t0_r3_c4_rr5;
  wire [15:0] t0_r3_c4_rr6;
  wire [15:0] t0_r3_c4_rr7;
  wire [15:0] t0_r3_c4_rr8;
  wire [15:0] t0_r3_c4_rr9;
  wire [15:0] t0_r3_c4_rr10;
  wire [15:0] t0_r3_c4_rr11;
  wire [15:0] t0_r3_c4_rr12;
  wire [15:0] t0_r3_c4_rr13;
  wire [15:0] t0_r3_c4_rr14;
  wire [15:0] t1_r3_c4_rr0;
  wire [15:0] t1_r3_c4_rr1;
  wire [15:0] t1_r3_c4_rr2;
  wire [15:0] t1_r3_c4_rr3;
  wire [15:0] t1_r3_c4_rr4;
  wire [15:0] t1_r3_c4_rr5;
  wire [15:0] t1_r3_c4_rr6;
  wire [15:0] t1_r3_c4_rr7;
  wire [15:0] t2_r3_c4_rr0;
  wire [15:0] t2_r3_c4_rr1;
  wire [15:0] t2_r3_c4_rr2;
  wire [15:0] t2_r3_c4_rr3;
  wire [15:0] t3_r3_c4_rr0;
  wire [15:0] t3_r3_c4_rr1;
  wire [15:0] t4_r3_c4_rr0;
  wire [15:0] t0_r3_c5_rr0;
  wire [15:0] t0_r3_c5_rr1;
  wire [15:0] t0_r3_c5_rr2;
  wire [15:0] t0_r3_c5_rr3;
  wire [15:0] t0_r3_c5_rr4;
  wire [15:0] t0_r3_c5_rr5;
  wire [15:0] t0_r3_c5_rr6;
  wire [15:0] t0_r3_c5_rr7;
  wire [15:0] t0_r3_c5_rr8;
  wire [15:0] t0_r3_c5_rr9;
  wire [15:0] t0_r3_c5_rr10;
  wire [15:0] t0_r3_c5_rr11;
  wire [15:0] t0_r3_c5_rr12;
  wire [15:0] t0_r3_c5_rr13;
  wire [15:0] t0_r3_c5_rr14;
  wire [15:0] t1_r3_c5_rr0;
  wire [15:0] t1_r3_c5_rr1;
  wire [15:0] t1_r3_c5_rr2;
  wire [15:0] t1_r3_c5_rr3;
  wire [15:0] t1_r3_c5_rr4;
  wire [15:0] t1_r3_c5_rr5;
  wire [15:0] t1_r3_c5_rr6;
  wire [15:0] t1_r3_c5_rr7;
  wire [15:0] t2_r3_c5_rr0;
  wire [15:0] t2_r3_c5_rr1;
  wire [15:0] t2_r3_c5_rr2;
  wire [15:0] t2_r3_c5_rr3;
  wire [15:0] t3_r3_c5_rr0;
  wire [15:0] t3_r3_c5_rr1;
  wire [15:0] t4_r3_c5_rr0;
  wire [15:0] t0_r3_c6_rr0;
  wire [15:0] t0_r3_c6_rr1;
  wire [15:0] t0_r3_c6_rr2;
  wire [15:0] t0_r3_c6_rr3;
  wire [15:0] t0_r3_c6_rr4;
  wire [15:0] t0_r3_c6_rr5;
  wire [15:0] t0_r3_c6_rr6;
  wire [15:0] t0_r3_c6_rr7;
  wire [15:0] t0_r3_c6_rr8;
  wire [15:0] t0_r3_c6_rr9;
  wire [15:0] t0_r3_c6_rr10;
  wire [15:0] t0_r3_c6_rr11;
  wire [15:0] t0_r3_c6_rr12;
  wire [15:0] t0_r3_c6_rr13;
  wire [15:0] t0_r3_c6_rr14;
  wire [15:0] t1_r3_c6_rr0;
  wire [15:0] t1_r3_c6_rr1;
  wire [15:0] t1_r3_c6_rr2;
  wire [15:0] t1_r3_c6_rr3;
  wire [15:0] t1_r3_c6_rr4;
  wire [15:0] t1_r3_c6_rr5;
  wire [15:0] t1_r3_c6_rr6;
  wire [15:0] t1_r3_c6_rr7;
  wire [15:0] t2_r3_c6_rr0;
  wire [15:0] t2_r3_c6_rr1;
  wire [15:0] t2_r3_c6_rr2;
  wire [15:0] t2_r3_c6_rr3;
  wire [15:0] t3_r3_c6_rr0;
  wire [15:0] t3_r3_c6_rr1;
  wire [15:0] t4_r3_c6_rr0;
  wire [15:0] t0_r3_c7_rr0;
  wire [15:0] t0_r3_c7_rr1;
  wire [15:0] t0_r3_c7_rr2;
  wire [15:0] t0_r3_c7_rr3;
  wire [15:0] t0_r3_c7_rr4;
  wire [15:0] t0_r3_c7_rr5;
  wire [15:0] t0_r3_c7_rr6;
  wire [15:0] t0_r3_c7_rr7;
  wire [15:0] t0_r3_c7_rr8;
  wire [15:0] t0_r3_c7_rr9;
  wire [15:0] t0_r3_c7_rr10;
  wire [15:0] t0_r3_c7_rr11;
  wire [15:0] t0_r3_c7_rr12;
  wire [15:0] t0_r3_c7_rr13;
  wire [15:0] t0_r3_c7_rr14;
  wire [15:0] t1_r3_c7_rr0;
  wire [15:0] t1_r3_c7_rr1;
  wire [15:0] t1_r3_c7_rr2;
  wire [15:0] t1_r3_c7_rr3;
  wire [15:0] t1_r3_c7_rr4;
  wire [15:0] t1_r3_c7_rr5;
  wire [15:0] t1_r3_c7_rr6;
  wire [15:0] t1_r3_c7_rr7;
  wire [15:0] t2_r3_c7_rr0;
  wire [15:0] t2_r3_c7_rr1;
  wire [15:0] t2_r3_c7_rr2;
  wire [15:0] t2_r3_c7_rr3;
  wire [15:0] t3_r3_c7_rr0;
  wire [15:0] t3_r3_c7_rr1;
  wire [15:0] t4_r3_c7_rr0;
  wire [15:0] t0_r3_c8_rr0;
  wire [15:0] t0_r3_c8_rr1;
  wire [15:0] t0_r3_c8_rr2;
  wire [15:0] t0_r3_c8_rr3;
  wire [15:0] t0_r3_c8_rr4;
  wire [15:0] t0_r3_c8_rr5;
  wire [15:0] t0_r3_c8_rr6;
  wire [15:0] t0_r3_c8_rr7;
  wire [15:0] t0_r3_c8_rr8;
  wire [15:0] t0_r3_c8_rr9;
  wire [15:0] t0_r3_c8_rr10;
  wire [15:0] t0_r3_c8_rr11;
  wire [15:0] t0_r3_c8_rr12;
  wire [15:0] t0_r3_c8_rr13;
  wire [15:0] t0_r3_c8_rr14;
  wire [15:0] t1_r3_c8_rr0;
  wire [15:0] t1_r3_c8_rr1;
  wire [15:0] t1_r3_c8_rr2;
  wire [15:0] t1_r3_c8_rr3;
  wire [15:0] t1_r3_c8_rr4;
  wire [15:0] t1_r3_c8_rr5;
  wire [15:0] t1_r3_c8_rr6;
  wire [15:0] t1_r3_c8_rr7;
  wire [15:0] t2_r3_c8_rr0;
  wire [15:0] t2_r3_c8_rr1;
  wire [15:0] t2_r3_c8_rr2;
  wire [15:0] t2_r3_c8_rr3;
  wire [15:0] t3_r3_c8_rr0;
  wire [15:0] t3_r3_c8_rr1;
  wire [15:0] t4_r3_c8_rr0;
  wire [15:0] t0_r3_c9_rr0;
  wire [15:0] t0_r3_c9_rr1;
  wire [15:0] t0_r3_c9_rr2;
  wire [15:0] t0_r3_c9_rr3;
  wire [15:0] t0_r3_c9_rr4;
  wire [15:0] t0_r3_c9_rr5;
  wire [15:0] t0_r3_c9_rr6;
  wire [15:0] t0_r3_c9_rr7;
  wire [15:0] t0_r3_c9_rr8;
  wire [15:0] t0_r3_c9_rr9;
  wire [15:0] t0_r3_c9_rr10;
  wire [15:0] t0_r3_c9_rr11;
  wire [15:0] t0_r3_c9_rr12;
  wire [15:0] t0_r3_c9_rr13;
  wire [15:0] t0_r3_c9_rr14;
  wire [15:0] t1_r3_c9_rr0;
  wire [15:0] t1_r3_c9_rr1;
  wire [15:0] t1_r3_c9_rr2;
  wire [15:0] t1_r3_c9_rr3;
  wire [15:0] t1_r3_c9_rr4;
  wire [15:0] t1_r3_c9_rr5;
  wire [15:0] t1_r3_c9_rr6;
  wire [15:0] t1_r3_c9_rr7;
  wire [15:0] t2_r3_c9_rr0;
  wire [15:0] t2_r3_c9_rr1;
  wire [15:0] t2_r3_c9_rr2;
  wire [15:0] t2_r3_c9_rr3;
  wire [15:0] t3_r3_c9_rr0;
  wire [15:0] t3_r3_c9_rr1;
  wire [15:0] t4_r3_c9_rr0;
  wire [15:0] t0_r3_c10_rr0;
  wire [15:0] t0_r3_c10_rr1;
  wire [15:0] t0_r3_c10_rr2;
  wire [15:0] t0_r3_c10_rr3;
  wire [15:0] t0_r3_c10_rr4;
  wire [15:0] t0_r3_c10_rr5;
  wire [15:0] t0_r3_c10_rr6;
  wire [15:0] t0_r3_c10_rr7;
  wire [15:0] t0_r3_c10_rr8;
  wire [15:0] t0_r3_c10_rr9;
  wire [15:0] t0_r3_c10_rr10;
  wire [15:0] t0_r3_c10_rr11;
  wire [15:0] t0_r3_c10_rr12;
  wire [15:0] t0_r3_c10_rr13;
  wire [15:0] t0_r3_c10_rr14;
  wire [15:0] t1_r3_c10_rr0;
  wire [15:0] t1_r3_c10_rr1;
  wire [15:0] t1_r3_c10_rr2;
  wire [15:0] t1_r3_c10_rr3;
  wire [15:0] t1_r3_c10_rr4;
  wire [15:0] t1_r3_c10_rr5;
  wire [15:0] t1_r3_c10_rr6;
  wire [15:0] t1_r3_c10_rr7;
  wire [15:0] t2_r3_c10_rr0;
  wire [15:0] t2_r3_c10_rr1;
  wire [15:0] t2_r3_c10_rr2;
  wire [15:0] t2_r3_c10_rr3;
  wire [15:0] t3_r3_c10_rr0;
  wire [15:0] t3_r3_c10_rr1;
  wire [15:0] t4_r3_c10_rr0;
  wire [15:0] t0_r3_c11_rr0;
  wire [15:0] t0_r3_c11_rr1;
  wire [15:0] t0_r3_c11_rr2;
  wire [15:0] t0_r3_c11_rr3;
  wire [15:0] t0_r3_c11_rr4;
  wire [15:0] t0_r3_c11_rr5;
  wire [15:0] t0_r3_c11_rr6;
  wire [15:0] t0_r3_c11_rr7;
  wire [15:0] t0_r3_c11_rr8;
  wire [15:0] t0_r3_c11_rr9;
  wire [15:0] t0_r3_c11_rr10;
  wire [15:0] t0_r3_c11_rr11;
  wire [15:0] t0_r3_c11_rr12;
  wire [15:0] t0_r3_c11_rr13;
  wire [15:0] t0_r3_c11_rr14;
  wire [15:0] t1_r3_c11_rr0;
  wire [15:0] t1_r3_c11_rr1;
  wire [15:0] t1_r3_c11_rr2;
  wire [15:0] t1_r3_c11_rr3;
  wire [15:0] t1_r3_c11_rr4;
  wire [15:0] t1_r3_c11_rr5;
  wire [15:0] t1_r3_c11_rr6;
  wire [15:0] t1_r3_c11_rr7;
  wire [15:0] t2_r3_c11_rr0;
  wire [15:0] t2_r3_c11_rr1;
  wire [15:0] t2_r3_c11_rr2;
  wire [15:0] t2_r3_c11_rr3;
  wire [15:0] t3_r3_c11_rr0;
  wire [15:0] t3_r3_c11_rr1;
  wire [15:0] t4_r3_c11_rr0;
  wire [15:0] t0_r3_c12_rr0;
  wire [15:0] t0_r3_c12_rr1;
  wire [15:0] t0_r3_c12_rr2;
  wire [15:0] t0_r3_c12_rr3;
  wire [15:0] t0_r3_c12_rr4;
  wire [15:0] t0_r3_c12_rr5;
  wire [15:0] t0_r3_c12_rr6;
  wire [15:0] t0_r3_c12_rr7;
  wire [15:0] t0_r3_c12_rr8;
  wire [15:0] t0_r3_c12_rr9;
  wire [15:0] t0_r3_c12_rr10;
  wire [15:0] t0_r3_c12_rr11;
  wire [15:0] t0_r3_c12_rr12;
  wire [15:0] t0_r3_c12_rr13;
  wire [15:0] t0_r3_c12_rr14;
  wire [15:0] t1_r3_c12_rr0;
  wire [15:0] t1_r3_c12_rr1;
  wire [15:0] t1_r3_c12_rr2;
  wire [15:0] t1_r3_c12_rr3;
  wire [15:0] t1_r3_c12_rr4;
  wire [15:0] t1_r3_c12_rr5;
  wire [15:0] t1_r3_c12_rr6;
  wire [15:0] t1_r3_c12_rr7;
  wire [15:0] t2_r3_c12_rr0;
  wire [15:0] t2_r3_c12_rr1;
  wire [15:0] t2_r3_c12_rr2;
  wire [15:0] t2_r3_c12_rr3;
  wire [15:0] t3_r3_c12_rr0;
  wire [15:0] t3_r3_c12_rr1;
  wire [15:0] t4_r3_c12_rr0;
  wire [15:0] t0_r3_c13_rr0;
  wire [15:0] t0_r3_c13_rr1;
  wire [15:0] t0_r3_c13_rr2;
  wire [15:0] t0_r3_c13_rr3;
  wire [15:0] t0_r3_c13_rr4;
  wire [15:0] t0_r3_c13_rr5;
  wire [15:0] t0_r3_c13_rr6;
  wire [15:0] t0_r3_c13_rr7;
  wire [15:0] t0_r3_c13_rr8;
  wire [15:0] t0_r3_c13_rr9;
  wire [15:0] t0_r3_c13_rr10;
  wire [15:0] t0_r3_c13_rr11;
  wire [15:0] t0_r3_c13_rr12;
  wire [15:0] t0_r3_c13_rr13;
  wire [15:0] t0_r3_c13_rr14;
  wire [15:0] t1_r3_c13_rr0;
  wire [15:0] t1_r3_c13_rr1;
  wire [15:0] t1_r3_c13_rr2;
  wire [15:0] t1_r3_c13_rr3;
  wire [15:0] t1_r3_c13_rr4;
  wire [15:0] t1_r3_c13_rr5;
  wire [15:0] t1_r3_c13_rr6;
  wire [15:0] t1_r3_c13_rr7;
  wire [15:0] t2_r3_c13_rr0;
  wire [15:0] t2_r3_c13_rr1;
  wire [15:0] t2_r3_c13_rr2;
  wire [15:0] t2_r3_c13_rr3;
  wire [15:0] t3_r3_c13_rr0;
  wire [15:0] t3_r3_c13_rr1;
  wire [15:0] t4_r3_c13_rr0;
  wire [15:0] t0_r3_c14_rr0;
  wire [15:0] t0_r3_c14_rr1;
  wire [15:0] t0_r3_c14_rr2;
  wire [15:0] t0_r3_c14_rr3;
  wire [15:0] t0_r3_c14_rr4;
  wire [15:0] t0_r3_c14_rr5;
  wire [15:0] t0_r3_c14_rr6;
  wire [15:0] t0_r3_c14_rr7;
  wire [15:0] t0_r3_c14_rr8;
  wire [15:0] t0_r3_c14_rr9;
  wire [15:0] t0_r3_c14_rr10;
  wire [15:0] t0_r3_c14_rr11;
  wire [15:0] t0_r3_c14_rr12;
  wire [15:0] t0_r3_c14_rr13;
  wire [15:0] t0_r3_c14_rr14;
  wire [15:0] t1_r3_c14_rr0;
  wire [15:0] t1_r3_c14_rr1;
  wire [15:0] t1_r3_c14_rr2;
  wire [15:0] t1_r3_c14_rr3;
  wire [15:0] t1_r3_c14_rr4;
  wire [15:0] t1_r3_c14_rr5;
  wire [15:0] t1_r3_c14_rr6;
  wire [15:0] t1_r3_c14_rr7;
  wire [15:0] t2_r3_c14_rr0;
  wire [15:0] t2_r3_c14_rr1;
  wire [15:0] t2_r3_c14_rr2;
  wire [15:0] t2_r3_c14_rr3;
  wire [15:0] t3_r3_c14_rr0;
  wire [15:0] t3_r3_c14_rr1;
  wire [15:0] t4_r3_c14_rr0;
  wire [15:0] t0_r4_c0_rr0;
  wire [15:0] t0_r4_c0_rr1;
  wire [15:0] t0_r4_c0_rr2;
  wire [15:0] t0_r4_c0_rr3;
  wire [15:0] t0_r4_c0_rr4;
  wire [15:0] t0_r4_c0_rr5;
  wire [15:0] t0_r4_c0_rr6;
  wire [15:0] t0_r4_c0_rr7;
  wire [15:0] t0_r4_c0_rr8;
  wire [15:0] t0_r4_c0_rr9;
  wire [15:0] t0_r4_c0_rr10;
  wire [15:0] t0_r4_c0_rr11;
  wire [15:0] t0_r4_c0_rr12;
  wire [15:0] t0_r4_c0_rr13;
  wire [15:0] t0_r4_c0_rr14;
  wire [15:0] t1_r4_c0_rr0;
  wire [15:0] t1_r4_c0_rr1;
  wire [15:0] t1_r4_c0_rr2;
  wire [15:0] t1_r4_c0_rr3;
  wire [15:0] t1_r4_c0_rr4;
  wire [15:0] t1_r4_c0_rr5;
  wire [15:0] t1_r4_c0_rr6;
  wire [15:0] t1_r4_c0_rr7;
  wire [15:0] t2_r4_c0_rr0;
  wire [15:0] t2_r4_c0_rr1;
  wire [15:0] t2_r4_c0_rr2;
  wire [15:0] t2_r4_c0_rr3;
  wire [15:0] t3_r4_c0_rr0;
  wire [15:0] t3_r4_c0_rr1;
  wire [15:0] t4_r4_c0_rr0;
  wire [15:0] t0_r4_c1_rr0;
  wire [15:0] t0_r4_c1_rr1;
  wire [15:0] t0_r4_c1_rr2;
  wire [15:0] t0_r4_c1_rr3;
  wire [15:0] t0_r4_c1_rr4;
  wire [15:0] t0_r4_c1_rr5;
  wire [15:0] t0_r4_c1_rr6;
  wire [15:0] t0_r4_c1_rr7;
  wire [15:0] t0_r4_c1_rr8;
  wire [15:0] t0_r4_c1_rr9;
  wire [15:0] t0_r4_c1_rr10;
  wire [15:0] t0_r4_c1_rr11;
  wire [15:0] t0_r4_c1_rr12;
  wire [15:0] t0_r4_c1_rr13;
  wire [15:0] t0_r4_c1_rr14;
  wire [15:0] t1_r4_c1_rr0;
  wire [15:0] t1_r4_c1_rr1;
  wire [15:0] t1_r4_c1_rr2;
  wire [15:0] t1_r4_c1_rr3;
  wire [15:0] t1_r4_c1_rr4;
  wire [15:0] t1_r4_c1_rr5;
  wire [15:0] t1_r4_c1_rr6;
  wire [15:0] t1_r4_c1_rr7;
  wire [15:0] t2_r4_c1_rr0;
  wire [15:0] t2_r4_c1_rr1;
  wire [15:0] t2_r4_c1_rr2;
  wire [15:0] t2_r4_c1_rr3;
  wire [15:0] t3_r4_c1_rr0;
  wire [15:0] t3_r4_c1_rr1;
  wire [15:0] t4_r4_c1_rr0;
  wire [15:0] t0_r4_c2_rr0;
  wire [15:0] t0_r4_c2_rr1;
  wire [15:0] t0_r4_c2_rr2;
  wire [15:0] t0_r4_c2_rr3;
  wire [15:0] t0_r4_c2_rr4;
  wire [15:0] t0_r4_c2_rr5;
  wire [15:0] t0_r4_c2_rr6;
  wire [15:0] t0_r4_c2_rr7;
  wire [15:0] t0_r4_c2_rr8;
  wire [15:0] t0_r4_c2_rr9;
  wire [15:0] t0_r4_c2_rr10;
  wire [15:0] t0_r4_c2_rr11;
  wire [15:0] t0_r4_c2_rr12;
  wire [15:0] t0_r4_c2_rr13;
  wire [15:0] t0_r4_c2_rr14;
  wire [15:0] t1_r4_c2_rr0;
  wire [15:0] t1_r4_c2_rr1;
  wire [15:0] t1_r4_c2_rr2;
  wire [15:0] t1_r4_c2_rr3;
  wire [15:0] t1_r4_c2_rr4;
  wire [15:0] t1_r4_c2_rr5;
  wire [15:0] t1_r4_c2_rr6;
  wire [15:0] t1_r4_c2_rr7;
  wire [15:0] t2_r4_c2_rr0;
  wire [15:0] t2_r4_c2_rr1;
  wire [15:0] t2_r4_c2_rr2;
  wire [15:0] t2_r4_c2_rr3;
  wire [15:0] t3_r4_c2_rr0;
  wire [15:0] t3_r4_c2_rr1;
  wire [15:0] t4_r4_c2_rr0;
  wire [15:0] t0_r4_c3_rr0;
  wire [15:0] t0_r4_c3_rr1;
  wire [15:0] t0_r4_c3_rr2;
  wire [15:0] t0_r4_c3_rr3;
  wire [15:0] t0_r4_c3_rr4;
  wire [15:0] t0_r4_c3_rr5;
  wire [15:0] t0_r4_c3_rr6;
  wire [15:0] t0_r4_c3_rr7;
  wire [15:0] t0_r4_c3_rr8;
  wire [15:0] t0_r4_c3_rr9;
  wire [15:0] t0_r4_c3_rr10;
  wire [15:0] t0_r4_c3_rr11;
  wire [15:0] t0_r4_c3_rr12;
  wire [15:0] t0_r4_c3_rr13;
  wire [15:0] t0_r4_c3_rr14;
  wire [15:0] t1_r4_c3_rr0;
  wire [15:0] t1_r4_c3_rr1;
  wire [15:0] t1_r4_c3_rr2;
  wire [15:0] t1_r4_c3_rr3;
  wire [15:0] t1_r4_c3_rr4;
  wire [15:0] t1_r4_c3_rr5;
  wire [15:0] t1_r4_c3_rr6;
  wire [15:0] t1_r4_c3_rr7;
  wire [15:0] t2_r4_c3_rr0;
  wire [15:0] t2_r4_c3_rr1;
  wire [15:0] t2_r4_c3_rr2;
  wire [15:0] t2_r4_c3_rr3;
  wire [15:0] t3_r4_c3_rr0;
  wire [15:0] t3_r4_c3_rr1;
  wire [15:0] t4_r4_c3_rr0;
  wire [15:0] t0_r4_c4_rr0;
  wire [15:0] t0_r4_c4_rr1;
  wire [15:0] t0_r4_c4_rr2;
  wire [15:0] t0_r4_c4_rr3;
  wire [15:0] t0_r4_c4_rr4;
  wire [15:0] t0_r4_c4_rr5;
  wire [15:0] t0_r4_c4_rr6;
  wire [15:0] t0_r4_c4_rr7;
  wire [15:0] t0_r4_c4_rr8;
  wire [15:0] t0_r4_c4_rr9;
  wire [15:0] t0_r4_c4_rr10;
  wire [15:0] t0_r4_c4_rr11;
  wire [15:0] t0_r4_c4_rr12;
  wire [15:0] t0_r4_c4_rr13;
  wire [15:0] t0_r4_c4_rr14;
  wire [15:0] t1_r4_c4_rr0;
  wire [15:0] t1_r4_c4_rr1;
  wire [15:0] t1_r4_c4_rr2;
  wire [15:0] t1_r4_c4_rr3;
  wire [15:0] t1_r4_c4_rr4;
  wire [15:0] t1_r4_c4_rr5;
  wire [15:0] t1_r4_c4_rr6;
  wire [15:0] t1_r4_c4_rr7;
  wire [15:0] t2_r4_c4_rr0;
  wire [15:0] t2_r4_c4_rr1;
  wire [15:0] t2_r4_c4_rr2;
  wire [15:0] t2_r4_c4_rr3;
  wire [15:0] t3_r4_c4_rr0;
  wire [15:0] t3_r4_c4_rr1;
  wire [15:0] t4_r4_c4_rr0;
  wire [15:0] t0_r4_c5_rr0;
  wire [15:0] t0_r4_c5_rr1;
  wire [15:0] t0_r4_c5_rr2;
  wire [15:0] t0_r4_c5_rr3;
  wire [15:0] t0_r4_c5_rr4;
  wire [15:0] t0_r4_c5_rr5;
  wire [15:0] t0_r4_c5_rr6;
  wire [15:0] t0_r4_c5_rr7;
  wire [15:0] t0_r4_c5_rr8;
  wire [15:0] t0_r4_c5_rr9;
  wire [15:0] t0_r4_c5_rr10;
  wire [15:0] t0_r4_c5_rr11;
  wire [15:0] t0_r4_c5_rr12;
  wire [15:0] t0_r4_c5_rr13;
  wire [15:0] t0_r4_c5_rr14;
  wire [15:0] t1_r4_c5_rr0;
  wire [15:0] t1_r4_c5_rr1;
  wire [15:0] t1_r4_c5_rr2;
  wire [15:0] t1_r4_c5_rr3;
  wire [15:0] t1_r4_c5_rr4;
  wire [15:0] t1_r4_c5_rr5;
  wire [15:0] t1_r4_c5_rr6;
  wire [15:0] t1_r4_c5_rr7;
  wire [15:0] t2_r4_c5_rr0;
  wire [15:0] t2_r4_c5_rr1;
  wire [15:0] t2_r4_c5_rr2;
  wire [15:0] t2_r4_c5_rr3;
  wire [15:0] t3_r4_c5_rr0;
  wire [15:0] t3_r4_c5_rr1;
  wire [15:0] t4_r4_c5_rr0;
  wire [15:0] t0_r4_c6_rr0;
  wire [15:0] t0_r4_c6_rr1;
  wire [15:0] t0_r4_c6_rr2;
  wire [15:0] t0_r4_c6_rr3;
  wire [15:0] t0_r4_c6_rr4;
  wire [15:0] t0_r4_c6_rr5;
  wire [15:0] t0_r4_c6_rr6;
  wire [15:0] t0_r4_c6_rr7;
  wire [15:0] t0_r4_c6_rr8;
  wire [15:0] t0_r4_c6_rr9;
  wire [15:0] t0_r4_c6_rr10;
  wire [15:0] t0_r4_c6_rr11;
  wire [15:0] t0_r4_c6_rr12;
  wire [15:0] t0_r4_c6_rr13;
  wire [15:0] t0_r4_c6_rr14;
  wire [15:0] t1_r4_c6_rr0;
  wire [15:0] t1_r4_c6_rr1;
  wire [15:0] t1_r4_c6_rr2;
  wire [15:0] t1_r4_c6_rr3;
  wire [15:0] t1_r4_c6_rr4;
  wire [15:0] t1_r4_c6_rr5;
  wire [15:0] t1_r4_c6_rr6;
  wire [15:0] t1_r4_c6_rr7;
  wire [15:0] t2_r4_c6_rr0;
  wire [15:0] t2_r4_c6_rr1;
  wire [15:0] t2_r4_c6_rr2;
  wire [15:0] t2_r4_c6_rr3;
  wire [15:0] t3_r4_c6_rr0;
  wire [15:0] t3_r4_c6_rr1;
  wire [15:0] t4_r4_c6_rr0;
  wire [15:0] t0_r4_c7_rr0;
  wire [15:0] t0_r4_c7_rr1;
  wire [15:0] t0_r4_c7_rr2;
  wire [15:0] t0_r4_c7_rr3;
  wire [15:0] t0_r4_c7_rr4;
  wire [15:0] t0_r4_c7_rr5;
  wire [15:0] t0_r4_c7_rr6;
  wire [15:0] t0_r4_c7_rr7;
  wire [15:0] t0_r4_c7_rr8;
  wire [15:0] t0_r4_c7_rr9;
  wire [15:0] t0_r4_c7_rr10;
  wire [15:0] t0_r4_c7_rr11;
  wire [15:0] t0_r4_c7_rr12;
  wire [15:0] t0_r4_c7_rr13;
  wire [15:0] t0_r4_c7_rr14;
  wire [15:0] t1_r4_c7_rr0;
  wire [15:0] t1_r4_c7_rr1;
  wire [15:0] t1_r4_c7_rr2;
  wire [15:0] t1_r4_c7_rr3;
  wire [15:0] t1_r4_c7_rr4;
  wire [15:0] t1_r4_c7_rr5;
  wire [15:0] t1_r4_c7_rr6;
  wire [15:0] t1_r4_c7_rr7;
  wire [15:0] t2_r4_c7_rr0;
  wire [15:0] t2_r4_c7_rr1;
  wire [15:0] t2_r4_c7_rr2;
  wire [15:0] t2_r4_c7_rr3;
  wire [15:0] t3_r4_c7_rr0;
  wire [15:0] t3_r4_c7_rr1;
  wire [15:0] t4_r4_c7_rr0;
  wire [15:0] t0_r4_c8_rr0;
  wire [15:0] t0_r4_c8_rr1;
  wire [15:0] t0_r4_c8_rr2;
  wire [15:0] t0_r4_c8_rr3;
  wire [15:0] t0_r4_c8_rr4;
  wire [15:0] t0_r4_c8_rr5;
  wire [15:0] t0_r4_c8_rr6;
  wire [15:0] t0_r4_c8_rr7;
  wire [15:0] t0_r4_c8_rr8;
  wire [15:0] t0_r4_c8_rr9;
  wire [15:0] t0_r4_c8_rr10;
  wire [15:0] t0_r4_c8_rr11;
  wire [15:0] t0_r4_c8_rr12;
  wire [15:0] t0_r4_c8_rr13;
  wire [15:0] t0_r4_c8_rr14;
  wire [15:0] t1_r4_c8_rr0;
  wire [15:0] t1_r4_c8_rr1;
  wire [15:0] t1_r4_c8_rr2;
  wire [15:0] t1_r4_c8_rr3;
  wire [15:0] t1_r4_c8_rr4;
  wire [15:0] t1_r4_c8_rr5;
  wire [15:0] t1_r4_c8_rr6;
  wire [15:0] t1_r4_c8_rr7;
  wire [15:0] t2_r4_c8_rr0;
  wire [15:0] t2_r4_c8_rr1;
  wire [15:0] t2_r4_c8_rr2;
  wire [15:0] t2_r4_c8_rr3;
  wire [15:0] t3_r4_c8_rr0;
  wire [15:0] t3_r4_c8_rr1;
  wire [15:0] t4_r4_c8_rr0;
  wire [15:0] t0_r4_c9_rr0;
  wire [15:0] t0_r4_c9_rr1;
  wire [15:0] t0_r4_c9_rr2;
  wire [15:0] t0_r4_c9_rr3;
  wire [15:0] t0_r4_c9_rr4;
  wire [15:0] t0_r4_c9_rr5;
  wire [15:0] t0_r4_c9_rr6;
  wire [15:0] t0_r4_c9_rr7;
  wire [15:0] t0_r4_c9_rr8;
  wire [15:0] t0_r4_c9_rr9;
  wire [15:0] t0_r4_c9_rr10;
  wire [15:0] t0_r4_c9_rr11;
  wire [15:0] t0_r4_c9_rr12;
  wire [15:0] t0_r4_c9_rr13;
  wire [15:0] t0_r4_c9_rr14;
  wire [15:0] t1_r4_c9_rr0;
  wire [15:0] t1_r4_c9_rr1;
  wire [15:0] t1_r4_c9_rr2;
  wire [15:0] t1_r4_c9_rr3;
  wire [15:0] t1_r4_c9_rr4;
  wire [15:0] t1_r4_c9_rr5;
  wire [15:0] t1_r4_c9_rr6;
  wire [15:0] t1_r4_c9_rr7;
  wire [15:0] t2_r4_c9_rr0;
  wire [15:0] t2_r4_c9_rr1;
  wire [15:0] t2_r4_c9_rr2;
  wire [15:0] t2_r4_c9_rr3;
  wire [15:0] t3_r4_c9_rr0;
  wire [15:0] t3_r4_c9_rr1;
  wire [15:0] t4_r4_c9_rr0;
  wire [15:0] t0_r4_c10_rr0;
  wire [15:0] t0_r4_c10_rr1;
  wire [15:0] t0_r4_c10_rr2;
  wire [15:0] t0_r4_c10_rr3;
  wire [15:0] t0_r4_c10_rr4;
  wire [15:0] t0_r4_c10_rr5;
  wire [15:0] t0_r4_c10_rr6;
  wire [15:0] t0_r4_c10_rr7;
  wire [15:0] t0_r4_c10_rr8;
  wire [15:0] t0_r4_c10_rr9;
  wire [15:0] t0_r4_c10_rr10;
  wire [15:0] t0_r4_c10_rr11;
  wire [15:0] t0_r4_c10_rr12;
  wire [15:0] t0_r4_c10_rr13;
  wire [15:0] t0_r4_c10_rr14;
  wire [15:0] t1_r4_c10_rr0;
  wire [15:0] t1_r4_c10_rr1;
  wire [15:0] t1_r4_c10_rr2;
  wire [15:0] t1_r4_c10_rr3;
  wire [15:0] t1_r4_c10_rr4;
  wire [15:0] t1_r4_c10_rr5;
  wire [15:0] t1_r4_c10_rr6;
  wire [15:0] t1_r4_c10_rr7;
  wire [15:0] t2_r4_c10_rr0;
  wire [15:0] t2_r4_c10_rr1;
  wire [15:0] t2_r4_c10_rr2;
  wire [15:0] t2_r4_c10_rr3;
  wire [15:0] t3_r4_c10_rr0;
  wire [15:0] t3_r4_c10_rr1;
  wire [15:0] t4_r4_c10_rr0;
  wire [15:0] t0_r4_c11_rr0;
  wire [15:0] t0_r4_c11_rr1;
  wire [15:0] t0_r4_c11_rr2;
  wire [15:0] t0_r4_c11_rr3;
  wire [15:0] t0_r4_c11_rr4;
  wire [15:0] t0_r4_c11_rr5;
  wire [15:0] t0_r4_c11_rr6;
  wire [15:0] t0_r4_c11_rr7;
  wire [15:0] t0_r4_c11_rr8;
  wire [15:0] t0_r4_c11_rr9;
  wire [15:0] t0_r4_c11_rr10;
  wire [15:0] t0_r4_c11_rr11;
  wire [15:0] t0_r4_c11_rr12;
  wire [15:0] t0_r4_c11_rr13;
  wire [15:0] t0_r4_c11_rr14;
  wire [15:0] t1_r4_c11_rr0;
  wire [15:0] t1_r4_c11_rr1;
  wire [15:0] t1_r4_c11_rr2;
  wire [15:0] t1_r4_c11_rr3;
  wire [15:0] t1_r4_c11_rr4;
  wire [15:0] t1_r4_c11_rr5;
  wire [15:0] t1_r4_c11_rr6;
  wire [15:0] t1_r4_c11_rr7;
  wire [15:0] t2_r4_c11_rr0;
  wire [15:0] t2_r4_c11_rr1;
  wire [15:0] t2_r4_c11_rr2;
  wire [15:0] t2_r4_c11_rr3;
  wire [15:0] t3_r4_c11_rr0;
  wire [15:0] t3_r4_c11_rr1;
  wire [15:0] t4_r4_c11_rr0;
  wire [15:0] t0_r4_c12_rr0;
  wire [15:0] t0_r4_c12_rr1;
  wire [15:0] t0_r4_c12_rr2;
  wire [15:0] t0_r4_c12_rr3;
  wire [15:0] t0_r4_c12_rr4;
  wire [15:0] t0_r4_c12_rr5;
  wire [15:0] t0_r4_c12_rr6;
  wire [15:0] t0_r4_c12_rr7;
  wire [15:0] t0_r4_c12_rr8;
  wire [15:0] t0_r4_c12_rr9;
  wire [15:0] t0_r4_c12_rr10;
  wire [15:0] t0_r4_c12_rr11;
  wire [15:0] t0_r4_c12_rr12;
  wire [15:0] t0_r4_c12_rr13;
  wire [15:0] t0_r4_c12_rr14;
  wire [15:0] t1_r4_c12_rr0;
  wire [15:0] t1_r4_c12_rr1;
  wire [15:0] t1_r4_c12_rr2;
  wire [15:0] t1_r4_c12_rr3;
  wire [15:0] t1_r4_c12_rr4;
  wire [15:0] t1_r4_c12_rr5;
  wire [15:0] t1_r4_c12_rr6;
  wire [15:0] t1_r4_c12_rr7;
  wire [15:0] t2_r4_c12_rr0;
  wire [15:0] t2_r4_c12_rr1;
  wire [15:0] t2_r4_c12_rr2;
  wire [15:0] t2_r4_c12_rr3;
  wire [15:0] t3_r4_c12_rr0;
  wire [15:0] t3_r4_c12_rr1;
  wire [15:0] t4_r4_c12_rr0;
  wire [15:0] t0_r4_c13_rr0;
  wire [15:0] t0_r4_c13_rr1;
  wire [15:0] t0_r4_c13_rr2;
  wire [15:0] t0_r4_c13_rr3;
  wire [15:0] t0_r4_c13_rr4;
  wire [15:0] t0_r4_c13_rr5;
  wire [15:0] t0_r4_c13_rr6;
  wire [15:0] t0_r4_c13_rr7;
  wire [15:0] t0_r4_c13_rr8;
  wire [15:0] t0_r4_c13_rr9;
  wire [15:0] t0_r4_c13_rr10;
  wire [15:0] t0_r4_c13_rr11;
  wire [15:0] t0_r4_c13_rr12;
  wire [15:0] t0_r4_c13_rr13;
  wire [15:0] t0_r4_c13_rr14;
  wire [15:0] t1_r4_c13_rr0;
  wire [15:0] t1_r4_c13_rr1;
  wire [15:0] t1_r4_c13_rr2;
  wire [15:0] t1_r4_c13_rr3;
  wire [15:0] t1_r4_c13_rr4;
  wire [15:0] t1_r4_c13_rr5;
  wire [15:0] t1_r4_c13_rr6;
  wire [15:0] t1_r4_c13_rr7;
  wire [15:0] t2_r4_c13_rr0;
  wire [15:0] t2_r4_c13_rr1;
  wire [15:0] t2_r4_c13_rr2;
  wire [15:0] t2_r4_c13_rr3;
  wire [15:0] t3_r4_c13_rr0;
  wire [15:0] t3_r4_c13_rr1;
  wire [15:0] t4_r4_c13_rr0;
  wire [15:0] t0_r4_c14_rr0;
  wire [15:0] t0_r4_c14_rr1;
  wire [15:0] t0_r4_c14_rr2;
  wire [15:0] t0_r4_c14_rr3;
  wire [15:0] t0_r4_c14_rr4;
  wire [15:0] t0_r4_c14_rr5;
  wire [15:0] t0_r4_c14_rr6;
  wire [15:0] t0_r4_c14_rr7;
  wire [15:0] t0_r4_c14_rr8;
  wire [15:0] t0_r4_c14_rr9;
  wire [15:0] t0_r4_c14_rr10;
  wire [15:0] t0_r4_c14_rr11;
  wire [15:0] t0_r4_c14_rr12;
  wire [15:0] t0_r4_c14_rr13;
  wire [15:0] t0_r4_c14_rr14;
  wire [15:0] t1_r4_c14_rr0;
  wire [15:0] t1_r4_c14_rr1;
  wire [15:0] t1_r4_c14_rr2;
  wire [15:0] t1_r4_c14_rr3;
  wire [15:0] t1_r4_c14_rr4;
  wire [15:0] t1_r4_c14_rr5;
  wire [15:0] t1_r4_c14_rr6;
  wire [15:0] t1_r4_c14_rr7;
  wire [15:0] t2_r4_c14_rr0;
  wire [15:0] t2_r4_c14_rr1;
  wire [15:0] t2_r4_c14_rr2;
  wire [15:0] t2_r4_c14_rr3;
  wire [15:0] t3_r4_c14_rr0;
  wire [15:0] t3_r4_c14_rr1;
  wire [15:0] t4_r4_c14_rr0;
  wire [15:0] t0_r5_c0_rr0;
  wire [15:0] t0_r5_c0_rr1;
  wire [15:0] t0_r5_c0_rr2;
  wire [15:0] t0_r5_c0_rr3;
  wire [15:0] t0_r5_c0_rr4;
  wire [15:0] t0_r5_c0_rr5;
  wire [15:0] t0_r5_c0_rr6;
  wire [15:0] t0_r5_c0_rr7;
  wire [15:0] t0_r5_c0_rr8;
  wire [15:0] t0_r5_c0_rr9;
  wire [15:0] t0_r5_c0_rr10;
  wire [15:0] t0_r5_c0_rr11;
  wire [15:0] t0_r5_c0_rr12;
  wire [15:0] t0_r5_c0_rr13;
  wire [15:0] t0_r5_c0_rr14;
  wire [15:0] t1_r5_c0_rr0;
  wire [15:0] t1_r5_c0_rr1;
  wire [15:0] t1_r5_c0_rr2;
  wire [15:0] t1_r5_c0_rr3;
  wire [15:0] t1_r5_c0_rr4;
  wire [15:0] t1_r5_c0_rr5;
  wire [15:0] t1_r5_c0_rr6;
  wire [15:0] t1_r5_c0_rr7;
  wire [15:0] t2_r5_c0_rr0;
  wire [15:0] t2_r5_c0_rr1;
  wire [15:0] t2_r5_c0_rr2;
  wire [15:0] t2_r5_c0_rr3;
  wire [15:0] t3_r5_c0_rr0;
  wire [15:0] t3_r5_c0_rr1;
  wire [15:0] t4_r5_c0_rr0;
  wire [15:0] t0_r5_c1_rr0;
  wire [15:0] t0_r5_c1_rr1;
  wire [15:0] t0_r5_c1_rr2;
  wire [15:0] t0_r5_c1_rr3;
  wire [15:0] t0_r5_c1_rr4;
  wire [15:0] t0_r5_c1_rr5;
  wire [15:0] t0_r5_c1_rr6;
  wire [15:0] t0_r5_c1_rr7;
  wire [15:0] t0_r5_c1_rr8;
  wire [15:0] t0_r5_c1_rr9;
  wire [15:0] t0_r5_c1_rr10;
  wire [15:0] t0_r5_c1_rr11;
  wire [15:0] t0_r5_c1_rr12;
  wire [15:0] t0_r5_c1_rr13;
  wire [15:0] t0_r5_c1_rr14;
  wire [15:0] t1_r5_c1_rr0;
  wire [15:0] t1_r5_c1_rr1;
  wire [15:0] t1_r5_c1_rr2;
  wire [15:0] t1_r5_c1_rr3;
  wire [15:0] t1_r5_c1_rr4;
  wire [15:0] t1_r5_c1_rr5;
  wire [15:0] t1_r5_c1_rr6;
  wire [15:0] t1_r5_c1_rr7;
  wire [15:0] t2_r5_c1_rr0;
  wire [15:0] t2_r5_c1_rr1;
  wire [15:0] t2_r5_c1_rr2;
  wire [15:0] t2_r5_c1_rr3;
  wire [15:0] t3_r5_c1_rr0;
  wire [15:0] t3_r5_c1_rr1;
  wire [15:0] t4_r5_c1_rr0;
  wire [15:0] t0_r5_c2_rr0;
  wire [15:0] t0_r5_c2_rr1;
  wire [15:0] t0_r5_c2_rr2;
  wire [15:0] t0_r5_c2_rr3;
  wire [15:0] t0_r5_c2_rr4;
  wire [15:0] t0_r5_c2_rr5;
  wire [15:0] t0_r5_c2_rr6;
  wire [15:0] t0_r5_c2_rr7;
  wire [15:0] t0_r5_c2_rr8;
  wire [15:0] t0_r5_c2_rr9;
  wire [15:0] t0_r5_c2_rr10;
  wire [15:0] t0_r5_c2_rr11;
  wire [15:0] t0_r5_c2_rr12;
  wire [15:0] t0_r5_c2_rr13;
  wire [15:0] t0_r5_c2_rr14;
  wire [15:0] t1_r5_c2_rr0;
  wire [15:0] t1_r5_c2_rr1;
  wire [15:0] t1_r5_c2_rr2;
  wire [15:0] t1_r5_c2_rr3;
  wire [15:0] t1_r5_c2_rr4;
  wire [15:0] t1_r5_c2_rr5;
  wire [15:0] t1_r5_c2_rr6;
  wire [15:0] t1_r5_c2_rr7;
  wire [15:0] t2_r5_c2_rr0;
  wire [15:0] t2_r5_c2_rr1;
  wire [15:0] t2_r5_c2_rr2;
  wire [15:0] t2_r5_c2_rr3;
  wire [15:0] t3_r5_c2_rr0;
  wire [15:0] t3_r5_c2_rr1;
  wire [15:0] t4_r5_c2_rr0;
  wire [15:0] t0_r5_c3_rr0;
  wire [15:0] t0_r5_c3_rr1;
  wire [15:0] t0_r5_c3_rr2;
  wire [15:0] t0_r5_c3_rr3;
  wire [15:0] t0_r5_c3_rr4;
  wire [15:0] t0_r5_c3_rr5;
  wire [15:0] t0_r5_c3_rr6;
  wire [15:0] t0_r5_c3_rr7;
  wire [15:0] t0_r5_c3_rr8;
  wire [15:0] t0_r5_c3_rr9;
  wire [15:0] t0_r5_c3_rr10;
  wire [15:0] t0_r5_c3_rr11;
  wire [15:0] t0_r5_c3_rr12;
  wire [15:0] t0_r5_c3_rr13;
  wire [15:0] t0_r5_c3_rr14;
  wire [15:0] t1_r5_c3_rr0;
  wire [15:0] t1_r5_c3_rr1;
  wire [15:0] t1_r5_c3_rr2;
  wire [15:0] t1_r5_c3_rr3;
  wire [15:0] t1_r5_c3_rr4;
  wire [15:0] t1_r5_c3_rr5;
  wire [15:0] t1_r5_c3_rr6;
  wire [15:0] t1_r5_c3_rr7;
  wire [15:0] t2_r5_c3_rr0;
  wire [15:0] t2_r5_c3_rr1;
  wire [15:0] t2_r5_c3_rr2;
  wire [15:0] t2_r5_c3_rr3;
  wire [15:0] t3_r5_c3_rr0;
  wire [15:0] t3_r5_c3_rr1;
  wire [15:0] t4_r5_c3_rr0;
  wire [15:0] t0_r5_c4_rr0;
  wire [15:0] t0_r5_c4_rr1;
  wire [15:0] t0_r5_c4_rr2;
  wire [15:0] t0_r5_c4_rr3;
  wire [15:0] t0_r5_c4_rr4;
  wire [15:0] t0_r5_c4_rr5;
  wire [15:0] t0_r5_c4_rr6;
  wire [15:0] t0_r5_c4_rr7;
  wire [15:0] t0_r5_c4_rr8;
  wire [15:0] t0_r5_c4_rr9;
  wire [15:0] t0_r5_c4_rr10;
  wire [15:0] t0_r5_c4_rr11;
  wire [15:0] t0_r5_c4_rr12;
  wire [15:0] t0_r5_c4_rr13;
  wire [15:0] t0_r5_c4_rr14;
  wire [15:0] t1_r5_c4_rr0;
  wire [15:0] t1_r5_c4_rr1;
  wire [15:0] t1_r5_c4_rr2;
  wire [15:0] t1_r5_c4_rr3;
  wire [15:0] t1_r5_c4_rr4;
  wire [15:0] t1_r5_c4_rr5;
  wire [15:0] t1_r5_c4_rr6;
  wire [15:0] t1_r5_c4_rr7;
  wire [15:0] t2_r5_c4_rr0;
  wire [15:0] t2_r5_c4_rr1;
  wire [15:0] t2_r5_c4_rr2;
  wire [15:0] t2_r5_c4_rr3;
  wire [15:0] t3_r5_c4_rr0;
  wire [15:0] t3_r5_c4_rr1;
  wire [15:0] t4_r5_c4_rr0;
  wire [15:0] t0_r5_c5_rr0;
  wire [15:0] t0_r5_c5_rr1;
  wire [15:0] t0_r5_c5_rr2;
  wire [15:0] t0_r5_c5_rr3;
  wire [15:0] t0_r5_c5_rr4;
  wire [15:0] t0_r5_c5_rr5;
  wire [15:0] t0_r5_c5_rr6;
  wire [15:0] t0_r5_c5_rr7;
  wire [15:0] t0_r5_c5_rr8;
  wire [15:0] t0_r5_c5_rr9;
  wire [15:0] t0_r5_c5_rr10;
  wire [15:0] t0_r5_c5_rr11;
  wire [15:0] t0_r5_c5_rr12;
  wire [15:0] t0_r5_c5_rr13;
  wire [15:0] t0_r5_c5_rr14;
  wire [15:0] t1_r5_c5_rr0;
  wire [15:0] t1_r5_c5_rr1;
  wire [15:0] t1_r5_c5_rr2;
  wire [15:0] t1_r5_c5_rr3;
  wire [15:0] t1_r5_c5_rr4;
  wire [15:0] t1_r5_c5_rr5;
  wire [15:0] t1_r5_c5_rr6;
  wire [15:0] t1_r5_c5_rr7;
  wire [15:0] t2_r5_c5_rr0;
  wire [15:0] t2_r5_c5_rr1;
  wire [15:0] t2_r5_c5_rr2;
  wire [15:0] t2_r5_c5_rr3;
  wire [15:0] t3_r5_c5_rr0;
  wire [15:0] t3_r5_c5_rr1;
  wire [15:0] t4_r5_c5_rr0;
  wire [15:0] t0_r5_c6_rr0;
  wire [15:0] t0_r5_c6_rr1;
  wire [15:0] t0_r5_c6_rr2;
  wire [15:0] t0_r5_c6_rr3;
  wire [15:0] t0_r5_c6_rr4;
  wire [15:0] t0_r5_c6_rr5;
  wire [15:0] t0_r5_c6_rr6;
  wire [15:0] t0_r5_c6_rr7;
  wire [15:0] t0_r5_c6_rr8;
  wire [15:0] t0_r5_c6_rr9;
  wire [15:0] t0_r5_c6_rr10;
  wire [15:0] t0_r5_c6_rr11;
  wire [15:0] t0_r5_c6_rr12;
  wire [15:0] t0_r5_c6_rr13;
  wire [15:0] t0_r5_c6_rr14;
  wire [15:0] t1_r5_c6_rr0;
  wire [15:0] t1_r5_c6_rr1;
  wire [15:0] t1_r5_c6_rr2;
  wire [15:0] t1_r5_c6_rr3;
  wire [15:0] t1_r5_c6_rr4;
  wire [15:0] t1_r5_c6_rr5;
  wire [15:0] t1_r5_c6_rr6;
  wire [15:0] t1_r5_c6_rr7;
  wire [15:0] t2_r5_c6_rr0;
  wire [15:0] t2_r5_c6_rr1;
  wire [15:0] t2_r5_c6_rr2;
  wire [15:0] t2_r5_c6_rr3;
  wire [15:0] t3_r5_c6_rr0;
  wire [15:0] t3_r5_c6_rr1;
  wire [15:0] t4_r5_c6_rr0;
  wire [15:0] t0_r5_c7_rr0;
  wire [15:0] t0_r5_c7_rr1;
  wire [15:0] t0_r5_c7_rr2;
  wire [15:0] t0_r5_c7_rr3;
  wire [15:0] t0_r5_c7_rr4;
  wire [15:0] t0_r5_c7_rr5;
  wire [15:0] t0_r5_c7_rr6;
  wire [15:0] t0_r5_c7_rr7;
  wire [15:0] t0_r5_c7_rr8;
  wire [15:0] t0_r5_c7_rr9;
  wire [15:0] t0_r5_c7_rr10;
  wire [15:0] t0_r5_c7_rr11;
  wire [15:0] t0_r5_c7_rr12;
  wire [15:0] t0_r5_c7_rr13;
  wire [15:0] t0_r5_c7_rr14;
  wire [15:0] t1_r5_c7_rr0;
  wire [15:0] t1_r5_c7_rr1;
  wire [15:0] t1_r5_c7_rr2;
  wire [15:0] t1_r5_c7_rr3;
  wire [15:0] t1_r5_c7_rr4;
  wire [15:0] t1_r5_c7_rr5;
  wire [15:0] t1_r5_c7_rr6;
  wire [15:0] t1_r5_c7_rr7;
  wire [15:0] t2_r5_c7_rr0;
  wire [15:0] t2_r5_c7_rr1;
  wire [15:0] t2_r5_c7_rr2;
  wire [15:0] t2_r5_c7_rr3;
  wire [15:0] t3_r5_c7_rr0;
  wire [15:0] t3_r5_c7_rr1;
  wire [15:0] t4_r5_c7_rr0;
  wire [15:0] t0_r5_c8_rr0;
  wire [15:0] t0_r5_c8_rr1;
  wire [15:0] t0_r5_c8_rr2;
  wire [15:0] t0_r5_c8_rr3;
  wire [15:0] t0_r5_c8_rr4;
  wire [15:0] t0_r5_c8_rr5;
  wire [15:0] t0_r5_c8_rr6;
  wire [15:0] t0_r5_c8_rr7;
  wire [15:0] t0_r5_c8_rr8;
  wire [15:0] t0_r5_c8_rr9;
  wire [15:0] t0_r5_c8_rr10;
  wire [15:0] t0_r5_c8_rr11;
  wire [15:0] t0_r5_c8_rr12;
  wire [15:0] t0_r5_c8_rr13;
  wire [15:0] t0_r5_c8_rr14;
  wire [15:0] t1_r5_c8_rr0;
  wire [15:0] t1_r5_c8_rr1;
  wire [15:0] t1_r5_c8_rr2;
  wire [15:0] t1_r5_c8_rr3;
  wire [15:0] t1_r5_c8_rr4;
  wire [15:0] t1_r5_c8_rr5;
  wire [15:0] t1_r5_c8_rr6;
  wire [15:0] t1_r5_c8_rr7;
  wire [15:0] t2_r5_c8_rr0;
  wire [15:0] t2_r5_c8_rr1;
  wire [15:0] t2_r5_c8_rr2;
  wire [15:0] t2_r5_c8_rr3;
  wire [15:0] t3_r5_c8_rr0;
  wire [15:0] t3_r5_c8_rr1;
  wire [15:0] t4_r5_c8_rr0;
  wire [15:0] t0_r5_c9_rr0;
  wire [15:0] t0_r5_c9_rr1;
  wire [15:0] t0_r5_c9_rr2;
  wire [15:0] t0_r5_c9_rr3;
  wire [15:0] t0_r5_c9_rr4;
  wire [15:0] t0_r5_c9_rr5;
  wire [15:0] t0_r5_c9_rr6;
  wire [15:0] t0_r5_c9_rr7;
  wire [15:0] t0_r5_c9_rr8;
  wire [15:0] t0_r5_c9_rr9;
  wire [15:0] t0_r5_c9_rr10;
  wire [15:0] t0_r5_c9_rr11;
  wire [15:0] t0_r5_c9_rr12;
  wire [15:0] t0_r5_c9_rr13;
  wire [15:0] t0_r5_c9_rr14;
  wire [15:0] t1_r5_c9_rr0;
  wire [15:0] t1_r5_c9_rr1;
  wire [15:0] t1_r5_c9_rr2;
  wire [15:0] t1_r5_c9_rr3;
  wire [15:0] t1_r5_c9_rr4;
  wire [15:0] t1_r5_c9_rr5;
  wire [15:0] t1_r5_c9_rr6;
  wire [15:0] t1_r5_c9_rr7;
  wire [15:0] t2_r5_c9_rr0;
  wire [15:0] t2_r5_c9_rr1;
  wire [15:0] t2_r5_c9_rr2;
  wire [15:0] t2_r5_c9_rr3;
  wire [15:0] t3_r5_c9_rr0;
  wire [15:0] t3_r5_c9_rr1;
  wire [15:0] t4_r5_c9_rr0;
  wire [15:0] t0_r5_c10_rr0;
  wire [15:0] t0_r5_c10_rr1;
  wire [15:0] t0_r5_c10_rr2;
  wire [15:0] t0_r5_c10_rr3;
  wire [15:0] t0_r5_c10_rr4;
  wire [15:0] t0_r5_c10_rr5;
  wire [15:0] t0_r5_c10_rr6;
  wire [15:0] t0_r5_c10_rr7;
  wire [15:0] t0_r5_c10_rr8;
  wire [15:0] t0_r5_c10_rr9;
  wire [15:0] t0_r5_c10_rr10;
  wire [15:0] t0_r5_c10_rr11;
  wire [15:0] t0_r5_c10_rr12;
  wire [15:0] t0_r5_c10_rr13;
  wire [15:0] t0_r5_c10_rr14;
  wire [15:0] t1_r5_c10_rr0;
  wire [15:0] t1_r5_c10_rr1;
  wire [15:0] t1_r5_c10_rr2;
  wire [15:0] t1_r5_c10_rr3;
  wire [15:0] t1_r5_c10_rr4;
  wire [15:0] t1_r5_c10_rr5;
  wire [15:0] t1_r5_c10_rr6;
  wire [15:0] t1_r5_c10_rr7;
  wire [15:0] t2_r5_c10_rr0;
  wire [15:0] t2_r5_c10_rr1;
  wire [15:0] t2_r5_c10_rr2;
  wire [15:0] t2_r5_c10_rr3;
  wire [15:0] t3_r5_c10_rr0;
  wire [15:0] t3_r5_c10_rr1;
  wire [15:0] t4_r5_c10_rr0;
  wire [15:0] t0_r5_c11_rr0;
  wire [15:0] t0_r5_c11_rr1;
  wire [15:0] t0_r5_c11_rr2;
  wire [15:0] t0_r5_c11_rr3;
  wire [15:0] t0_r5_c11_rr4;
  wire [15:0] t0_r5_c11_rr5;
  wire [15:0] t0_r5_c11_rr6;
  wire [15:0] t0_r5_c11_rr7;
  wire [15:0] t0_r5_c11_rr8;
  wire [15:0] t0_r5_c11_rr9;
  wire [15:0] t0_r5_c11_rr10;
  wire [15:0] t0_r5_c11_rr11;
  wire [15:0] t0_r5_c11_rr12;
  wire [15:0] t0_r5_c11_rr13;
  wire [15:0] t0_r5_c11_rr14;
  wire [15:0] t1_r5_c11_rr0;
  wire [15:0] t1_r5_c11_rr1;
  wire [15:0] t1_r5_c11_rr2;
  wire [15:0] t1_r5_c11_rr3;
  wire [15:0] t1_r5_c11_rr4;
  wire [15:0] t1_r5_c11_rr5;
  wire [15:0] t1_r5_c11_rr6;
  wire [15:0] t1_r5_c11_rr7;
  wire [15:0] t2_r5_c11_rr0;
  wire [15:0] t2_r5_c11_rr1;
  wire [15:0] t2_r5_c11_rr2;
  wire [15:0] t2_r5_c11_rr3;
  wire [15:0] t3_r5_c11_rr0;
  wire [15:0] t3_r5_c11_rr1;
  wire [15:0] t4_r5_c11_rr0;
  wire [15:0] t0_r5_c12_rr0;
  wire [15:0] t0_r5_c12_rr1;
  wire [15:0] t0_r5_c12_rr2;
  wire [15:0] t0_r5_c12_rr3;
  wire [15:0] t0_r5_c12_rr4;
  wire [15:0] t0_r5_c12_rr5;
  wire [15:0] t0_r5_c12_rr6;
  wire [15:0] t0_r5_c12_rr7;
  wire [15:0] t0_r5_c12_rr8;
  wire [15:0] t0_r5_c12_rr9;
  wire [15:0] t0_r5_c12_rr10;
  wire [15:0] t0_r5_c12_rr11;
  wire [15:0] t0_r5_c12_rr12;
  wire [15:0] t0_r5_c12_rr13;
  wire [15:0] t0_r5_c12_rr14;
  wire [15:0] t1_r5_c12_rr0;
  wire [15:0] t1_r5_c12_rr1;
  wire [15:0] t1_r5_c12_rr2;
  wire [15:0] t1_r5_c12_rr3;
  wire [15:0] t1_r5_c12_rr4;
  wire [15:0] t1_r5_c12_rr5;
  wire [15:0] t1_r5_c12_rr6;
  wire [15:0] t1_r5_c12_rr7;
  wire [15:0] t2_r5_c12_rr0;
  wire [15:0] t2_r5_c12_rr1;
  wire [15:0] t2_r5_c12_rr2;
  wire [15:0] t2_r5_c12_rr3;
  wire [15:0] t3_r5_c12_rr0;
  wire [15:0] t3_r5_c12_rr1;
  wire [15:0] t4_r5_c12_rr0;
  wire [15:0] t0_r5_c13_rr0;
  wire [15:0] t0_r5_c13_rr1;
  wire [15:0] t0_r5_c13_rr2;
  wire [15:0] t0_r5_c13_rr3;
  wire [15:0] t0_r5_c13_rr4;
  wire [15:0] t0_r5_c13_rr5;
  wire [15:0] t0_r5_c13_rr6;
  wire [15:0] t0_r5_c13_rr7;
  wire [15:0] t0_r5_c13_rr8;
  wire [15:0] t0_r5_c13_rr9;
  wire [15:0] t0_r5_c13_rr10;
  wire [15:0] t0_r5_c13_rr11;
  wire [15:0] t0_r5_c13_rr12;
  wire [15:0] t0_r5_c13_rr13;
  wire [15:0] t0_r5_c13_rr14;
  wire [15:0] t1_r5_c13_rr0;
  wire [15:0] t1_r5_c13_rr1;
  wire [15:0] t1_r5_c13_rr2;
  wire [15:0] t1_r5_c13_rr3;
  wire [15:0] t1_r5_c13_rr4;
  wire [15:0] t1_r5_c13_rr5;
  wire [15:0] t1_r5_c13_rr6;
  wire [15:0] t1_r5_c13_rr7;
  wire [15:0] t2_r5_c13_rr0;
  wire [15:0] t2_r5_c13_rr1;
  wire [15:0] t2_r5_c13_rr2;
  wire [15:0] t2_r5_c13_rr3;
  wire [15:0] t3_r5_c13_rr0;
  wire [15:0] t3_r5_c13_rr1;
  wire [15:0] t4_r5_c13_rr0;
  wire [15:0] t0_r5_c14_rr0;
  wire [15:0] t0_r5_c14_rr1;
  wire [15:0] t0_r5_c14_rr2;
  wire [15:0] t0_r5_c14_rr3;
  wire [15:0] t0_r5_c14_rr4;
  wire [15:0] t0_r5_c14_rr5;
  wire [15:0] t0_r5_c14_rr6;
  wire [15:0] t0_r5_c14_rr7;
  wire [15:0] t0_r5_c14_rr8;
  wire [15:0] t0_r5_c14_rr9;
  wire [15:0] t0_r5_c14_rr10;
  wire [15:0] t0_r5_c14_rr11;
  wire [15:0] t0_r5_c14_rr12;
  wire [15:0] t0_r5_c14_rr13;
  wire [15:0] t0_r5_c14_rr14;
  wire [15:0] t1_r5_c14_rr0;
  wire [15:0] t1_r5_c14_rr1;
  wire [15:0] t1_r5_c14_rr2;
  wire [15:0] t1_r5_c14_rr3;
  wire [15:0] t1_r5_c14_rr4;
  wire [15:0] t1_r5_c14_rr5;
  wire [15:0] t1_r5_c14_rr6;
  wire [15:0] t1_r5_c14_rr7;
  wire [15:0] t2_r5_c14_rr0;
  wire [15:0] t2_r5_c14_rr1;
  wire [15:0] t2_r5_c14_rr2;
  wire [15:0] t2_r5_c14_rr3;
  wire [15:0] t3_r5_c14_rr0;
  wire [15:0] t3_r5_c14_rr1;
  wire [15:0] t4_r5_c14_rr0;
  wire [15:0] t0_r6_c0_rr0;
  wire [15:0] t0_r6_c0_rr1;
  wire [15:0] t0_r6_c0_rr2;
  wire [15:0] t0_r6_c0_rr3;
  wire [15:0] t0_r6_c0_rr4;
  wire [15:0] t0_r6_c0_rr5;
  wire [15:0] t0_r6_c0_rr6;
  wire [15:0] t0_r6_c0_rr7;
  wire [15:0] t0_r6_c0_rr8;
  wire [15:0] t0_r6_c0_rr9;
  wire [15:0] t0_r6_c0_rr10;
  wire [15:0] t0_r6_c0_rr11;
  wire [15:0] t0_r6_c0_rr12;
  wire [15:0] t0_r6_c0_rr13;
  wire [15:0] t0_r6_c0_rr14;
  wire [15:0] t1_r6_c0_rr0;
  wire [15:0] t1_r6_c0_rr1;
  wire [15:0] t1_r6_c0_rr2;
  wire [15:0] t1_r6_c0_rr3;
  wire [15:0] t1_r6_c0_rr4;
  wire [15:0] t1_r6_c0_rr5;
  wire [15:0] t1_r6_c0_rr6;
  wire [15:0] t1_r6_c0_rr7;
  wire [15:0] t2_r6_c0_rr0;
  wire [15:0] t2_r6_c0_rr1;
  wire [15:0] t2_r6_c0_rr2;
  wire [15:0] t2_r6_c0_rr3;
  wire [15:0] t3_r6_c0_rr0;
  wire [15:0] t3_r6_c0_rr1;
  wire [15:0] t4_r6_c0_rr0;
  wire [15:0] t0_r6_c1_rr0;
  wire [15:0] t0_r6_c1_rr1;
  wire [15:0] t0_r6_c1_rr2;
  wire [15:0] t0_r6_c1_rr3;
  wire [15:0] t0_r6_c1_rr4;
  wire [15:0] t0_r6_c1_rr5;
  wire [15:0] t0_r6_c1_rr6;
  wire [15:0] t0_r6_c1_rr7;
  wire [15:0] t0_r6_c1_rr8;
  wire [15:0] t0_r6_c1_rr9;
  wire [15:0] t0_r6_c1_rr10;
  wire [15:0] t0_r6_c1_rr11;
  wire [15:0] t0_r6_c1_rr12;
  wire [15:0] t0_r6_c1_rr13;
  wire [15:0] t0_r6_c1_rr14;
  wire [15:0] t1_r6_c1_rr0;
  wire [15:0] t1_r6_c1_rr1;
  wire [15:0] t1_r6_c1_rr2;
  wire [15:0] t1_r6_c1_rr3;
  wire [15:0] t1_r6_c1_rr4;
  wire [15:0] t1_r6_c1_rr5;
  wire [15:0] t1_r6_c1_rr6;
  wire [15:0] t1_r6_c1_rr7;
  wire [15:0] t2_r6_c1_rr0;
  wire [15:0] t2_r6_c1_rr1;
  wire [15:0] t2_r6_c1_rr2;
  wire [15:0] t2_r6_c1_rr3;
  wire [15:0] t3_r6_c1_rr0;
  wire [15:0] t3_r6_c1_rr1;
  wire [15:0] t4_r6_c1_rr0;
  wire [15:0] t0_r6_c2_rr0;
  wire [15:0] t0_r6_c2_rr1;
  wire [15:0] t0_r6_c2_rr2;
  wire [15:0] t0_r6_c2_rr3;
  wire [15:0] t0_r6_c2_rr4;
  wire [15:0] t0_r6_c2_rr5;
  wire [15:0] t0_r6_c2_rr6;
  wire [15:0] t0_r6_c2_rr7;
  wire [15:0] t0_r6_c2_rr8;
  wire [15:0] t0_r6_c2_rr9;
  wire [15:0] t0_r6_c2_rr10;
  wire [15:0] t0_r6_c2_rr11;
  wire [15:0] t0_r6_c2_rr12;
  wire [15:0] t0_r6_c2_rr13;
  wire [15:0] t0_r6_c2_rr14;
  wire [15:0] t1_r6_c2_rr0;
  wire [15:0] t1_r6_c2_rr1;
  wire [15:0] t1_r6_c2_rr2;
  wire [15:0] t1_r6_c2_rr3;
  wire [15:0] t1_r6_c2_rr4;
  wire [15:0] t1_r6_c2_rr5;
  wire [15:0] t1_r6_c2_rr6;
  wire [15:0] t1_r6_c2_rr7;
  wire [15:0] t2_r6_c2_rr0;
  wire [15:0] t2_r6_c2_rr1;
  wire [15:0] t2_r6_c2_rr2;
  wire [15:0] t2_r6_c2_rr3;
  wire [15:0] t3_r6_c2_rr0;
  wire [15:0] t3_r6_c2_rr1;
  wire [15:0] t4_r6_c2_rr0;
  wire [15:0] t0_r6_c3_rr0;
  wire [15:0] t0_r6_c3_rr1;
  wire [15:0] t0_r6_c3_rr2;
  wire [15:0] t0_r6_c3_rr3;
  wire [15:0] t0_r6_c3_rr4;
  wire [15:0] t0_r6_c3_rr5;
  wire [15:0] t0_r6_c3_rr6;
  wire [15:0] t0_r6_c3_rr7;
  wire [15:0] t0_r6_c3_rr8;
  wire [15:0] t0_r6_c3_rr9;
  wire [15:0] t0_r6_c3_rr10;
  wire [15:0] t0_r6_c3_rr11;
  wire [15:0] t0_r6_c3_rr12;
  wire [15:0] t0_r6_c3_rr13;
  wire [15:0] t0_r6_c3_rr14;
  wire [15:0] t1_r6_c3_rr0;
  wire [15:0] t1_r6_c3_rr1;
  wire [15:0] t1_r6_c3_rr2;
  wire [15:0] t1_r6_c3_rr3;
  wire [15:0] t1_r6_c3_rr4;
  wire [15:0] t1_r6_c3_rr5;
  wire [15:0] t1_r6_c3_rr6;
  wire [15:0] t1_r6_c3_rr7;
  wire [15:0] t2_r6_c3_rr0;
  wire [15:0] t2_r6_c3_rr1;
  wire [15:0] t2_r6_c3_rr2;
  wire [15:0] t2_r6_c3_rr3;
  wire [15:0] t3_r6_c3_rr0;
  wire [15:0] t3_r6_c3_rr1;
  wire [15:0] t4_r6_c3_rr0;
  wire [15:0] t0_r6_c4_rr0;
  wire [15:0] t0_r6_c4_rr1;
  wire [15:0] t0_r6_c4_rr2;
  wire [15:0] t0_r6_c4_rr3;
  wire [15:0] t0_r6_c4_rr4;
  wire [15:0] t0_r6_c4_rr5;
  wire [15:0] t0_r6_c4_rr6;
  wire [15:0] t0_r6_c4_rr7;
  wire [15:0] t0_r6_c4_rr8;
  wire [15:0] t0_r6_c4_rr9;
  wire [15:0] t0_r6_c4_rr10;
  wire [15:0] t0_r6_c4_rr11;
  wire [15:0] t0_r6_c4_rr12;
  wire [15:0] t0_r6_c4_rr13;
  wire [15:0] t0_r6_c4_rr14;
  wire [15:0] t1_r6_c4_rr0;
  wire [15:0] t1_r6_c4_rr1;
  wire [15:0] t1_r6_c4_rr2;
  wire [15:0] t1_r6_c4_rr3;
  wire [15:0] t1_r6_c4_rr4;
  wire [15:0] t1_r6_c4_rr5;
  wire [15:0] t1_r6_c4_rr6;
  wire [15:0] t1_r6_c4_rr7;
  wire [15:0] t2_r6_c4_rr0;
  wire [15:0] t2_r6_c4_rr1;
  wire [15:0] t2_r6_c4_rr2;
  wire [15:0] t2_r6_c4_rr3;
  wire [15:0] t3_r6_c4_rr0;
  wire [15:0] t3_r6_c4_rr1;
  wire [15:0] t4_r6_c4_rr0;
  wire [15:0] t0_r6_c5_rr0;
  wire [15:0] t0_r6_c5_rr1;
  wire [15:0] t0_r6_c5_rr2;
  wire [15:0] t0_r6_c5_rr3;
  wire [15:0] t0_r6_c5_rr4;
  wire [15:0] t0_r6_c5_rr5;
  wire [15:0] t0_r6_c5_rr6;
  wire [15:0] t0_r6_c5_rr7;
  wire [15:0] t0_r6_c5_rr8;
  wire [15:0] t0_r6_c5_rr9;
  wire [15:0] t0_r6_c5_rr10;
  wire [15:0] t0_r6_c5_rr11;
  wire [15:0] t0_r6_c5_rr12;
  wire [15:0] t0_r6_c5_rr13;
  wire [15:0] t0_r6_c5_rr14;
  wire [15:0] t1_r6_c5_rr0;
  wire [15:0] t1_r6_c5_rr1;
  wire [15:0] t1_r6_c5_rr2;
  wire [15:0] t1_r6_c5_rr3;
  wire [15:0] t1_r6_c5_rr4;
  wire [15:0] t1_r6_c5_rr5;
  wire [15:0] t1_r6_c5_rr6;
  wire [15:0] t1_r6_c5_rr7;
  wire [15:0] t2_r6_c5_rr0;
  wire [15:0] t2_r6_c5_rr1;
  wire [15:0] t2_r6_c5_rr2;
  wire [15:0] t2_r6_c5_rr3;
  wire [15:0] t3_r6_c5_rr0;
  wire [15:0] t3_r6_c5_rr1;
  wire [15:0] t4_r6_c5_rr0;
  wire [15:0] t0_r6_c6_rr0;
  wire [15:0] t0_r6_c6_rr1;
  wire [15:0] t0_r6_c6_rr2;
  wire [15:0] t0_r6_c6_rr3;
  wire [15:0] t0_r6_c6_rr4;
  wire [15:0] t0_r6_c6_rr5;
  wire [15:0] t0_r6_c6_rr6;
  wire [15:0] t0_r6_c6_rr7;
  wire [15:0] t0_r6_c6_rr8;
  wire [15:0] t0_r6_c6_rr9;
  wire [15:0] t0_r6_c6_rr10;
  wire [15:0] t0_r6_c6_rr11;
  wire [15:0] t0_r6_c6_rr12;
  wire [15:0] t0_r6_c6_rr13;
  wire [15:0] t0_r6_c6_rr14;
  wire [15:0] t1_r6_c6_rr0;
  wire [15:0] t1_r6_c6_rr1;
  wire [15:0] t1_r6_c6_rr2;
  wire [15:0] t1_r6_c6_rr3;
  wire [15:0] t1_r6_c6_rr4;
  wire [15:0] t1_r6_c6_rr5;
  wire [15:0] t1_r6_c6_rr6;
  wire [15:0] t1_r6_c6_rr7;
  wire [15:0] t2_r6_c6_rr0;
  wire [15:0] t2_r6_c6_rr1;
  wire [15:0] t2_r6_c6_rr2;
  wire [15:0] t2_r6_c6_rr3;
  wire [15:0] t3_r6_c6_rr0;
  wire [15:0] t3_r6_c6_rr1;
  wire [15:0] t4_r6_c6_rr0;
  wire [15:0] t0_r6_c7_rr0;
  wire [15:0] t0_r6_c7_rr1;
  wire [15:0] t0_r6_c7_rr2;
  wire [15:0] t0_r6_c7_rr3;
  wire [15:0] t0_r6_c7_rr4;
  wire [15:0] t0_r6_c7_rr5;
  wire [15:0] t0_r6_c7_rr6;
  wire [15:0] t0_r6_c7_rr7;
  wire [15:0] t0_r6_c7_rr8;
  wire [15:0] t0_r6_c7_rr9;
  wire [15:0] t0_r6_c7_rr10;
  wire [15:0] t0_r6_c7_rr11;
  wire [15:0] t0_r6_c7_rr12;
  wire [15:0] t0_r6_c7_rr13;
  wire [15:0] t0_r6_c7_rr14;
  wire [15:0] t1_r6_c7_rr0;
  wire [15:0] t1_r6_c7_rr1;
  wire [15:0] t1_r6_c7_rr2;
  wire [15:0] t1_r6_c7_rr3;
  wire [15:0] t1_r6_c7_rr4;
  wire [15:0] t1_r6_c7_rr5;
  wire [15:0] t1_r6_c7_rr6;
  wire [15:0] t1_r6_c7_rr7;
  wire [15:0] t2_r6_c7_rr0;
  wire [15:0] t2_r6_c7_rr1;
  wire [15:0] t2_r6_c7_rr2;
  wire [15:0] t2_r6_c7_rr3;
  wire [15:0] t3_r6_c7_rr0;
  wire [15:0] t3_r6_c7_rr1;
  wire [15:0] t4_r6_c7_rr0;
  wire [15:0] t0_r6_c8_rr0;
  wire [15:0] t0_r6_c8_rr1;
  wire [15:0] t0_r6_c8_rr2;
  wire [15:0] t0_r6_c8_rr3;
  wire [15:0] t0_r6_c8_rr4;
  wire [15:0] t0_r6_c8_rr5;
  wire [15:0] t0_r6_c8_rr6;
  wire [15:0] t0_r6_c8_rr7;
  wire [15:0] t0_r6_c8_rr8;
  wire [15:0] t0_r6_c8_rr9;
  wire [15:0] t0_r6_c8_rr10;
  wire [15:0] t0_r6_c8_rr11;
  wire [15:0] t0_r6_c8_rr12;
  wire [15:0] t0_r6_c8_rr13;
  wire [15:0] t0_r6_c8_rr14;
  wire [15:0] t1_r6_c8_rr0;
  wire [15:0] t1_r6_c8_rr1;
  wire [15:0] t1_r6_c8_rr2;
  wire [15:0] t1_r6_c8_rr3;
  wire [15:0] t1_r6_c8_rr4;
  wire [15:0] t1_r6_c8_rr5;
  wire [15:0] t1_r6_c8_rr6;
  wire [15:0] t1_r6_c8_rr7;
  wire [15:0] t2_r6_c8_rr0;
  wire [15:0] t2_r6_c8_rr1;
  wire [15:0] t2_r6_c8_rr2;
  wire [15:0] t2_r6_c8_rr3;
  wire [15:0] t3_r6_c8_rr0;
  wire [15:0] t3_r6_c8_rr1;
  wire [15:0] t4_r6_c8_rr0;
  wire [15:0] t0_r6_c9_rr0;
  wire [15:0] t0_r6_c9_rr1;
  wire [15:0] t0_r6_c9_rr2;
  wire [15:0] t0_r6_c9_rr3;
  wire [15:0] t0_r6_c9_rr4;
  wire [15:0] t0_r6_c9_rr5;
  wire [15:0] t0_r6_c9_rr6;
  wire [15:0] t0_r6_c9_rr7;
  wire [15:0] t0_r6_c9_rr8;
  wire [15:0] t0_r6_c9_rr9;
  wire [15:0] t0_r6_c9_rr10;
  wire [15:0] t0_r6_c9_rr11;
  wire [15:0] t0_r6_c9_rr12;
  wire [15:0] t0_r6_c9_rr13;
  wire [15:0] t0_r6_c9_rr14;
  wire [15:0] t1_r6_c9_rr0;
  wire [15:0] t1_r6_c9_rr1;
  wire [15:0] t1_r6_c9_rr2;
  wire [15:0] t1_r6_c9_rr3;
  wire [15:0] t1_r6_c9_rr4;
  wire [15:0] t1_r6_c9_rr5;
  wire [15:0] t1_r6_c9_rr6;
  wire [15:0] t1_r6_c9_rr7;
  wire [15:0] t2_r6_c9_rr0;
  wire [15:0] t2_r6_c9_rr1;
  wire [15:0] t2_r6_c9_rr2;
  wire [15:0] t2_r6_c9_rr3;
  wire [15:0] t3_r6_c9_rr0;
  wire [15:0] t3_r6_c9_rr1;
  wire [15:0] t4_r6_c9_rr0;
  wire [15:0] t0_r6_c10_rr0;
  wire [15:0] t0_r6_c10_rr1;
  wire [15:0] t0_r6_c10_rr2;
  wire [15:0] t0_r6_c10_rr3;
  wire [15:0] t0_r6_c10_rr4;
  wire [15:0] t0_r6_c10_rr5;
  wire [15:0] t0_r6_c10_rr6;
  wire [15:0] t0_r6_c10_rr7;
  wire [15:0] t0_r6_c10_rr8;
  wire [15:0] t0_r6_c10_rr9;
  wire [15:0] t0_r6_c10_rr10;
  wire [15:0] t0_r6_c10_rr11;
  wire [15:0] t0_r6_c10_rr12;
  wire [15:0] t0_r6_c10_rr13;
  wire [15:0] t0_r6_c10_rr14;
  wire [15:0] t1_r6_c10_rr0;
  wire [15:0] t1_r6_c10_rr1;
  wire [15:0] t1_r6_c10_rr2;
  wire [15:0] t1_r6_c10_rr3;
  wire [15:0] t1_r6_c10_rr4;
  wire [15:0] t1_r6_c10_rr5;
  wire [15:0] t1_r6_c10_rr6;
  wire [15:0] t1_r6_c10_rr7;
  wire [15:0] t2_r6_c10_rr0;
  wire [15:0] t2_r6_c10_rr1;
  wire [15:0] t2_r6_c10_rr2;
  wire [15:0] t2_r6_c10_rr3;
  wire [15:0] t3_r6_c10_rr0;
  wire [15:0] t3_r6_c10_rr1;
  wire [15:0] t4_r6_c10_rr0;
  wire [15:0] t0_r6_c11_rr0;
  wire [15:0] t0_r6_c11_rr1;
  wire [15:0] t0_r6_c11_rr2;
  wire [15:0] t0_r6_c11_rr3;
  wire [15:0] t0_r6_c11_rr4;
  wire [15:0] t0_r6_c11_rr5;
  wire [15:0] t0_r6_c11_rr6;
  wire [15:0] t0_r6_c11_rr7;
  wire [15:0] t0_r6_c11_rr8;
  wire [15:0] t0_r6_c11_rr9;
  wire [15:0] t0_r6_c11_rr10;
  wire [15:0] t0_r6_c11_rr11;
  wire [15:0] t0_r6_c11_rr12;
  wire [15:0] t0_r6_c11_rr13;
  wire [15:0] t0_r6_c11_rr14;
  wire [15:0] t1_r6_c11_rr0;
  wire [15:0] t1_r6_c11_rr1;
  wire [15:0] t1_r6_c11_rr2;
  wire [15:0] t1_r6_c11_rr3;
  wire [15:0] t1_r6_c11_rr4;
  wire [15:0] t1_r6_c11_rr5;
  wire [15:0] t1_r6_c11_rr6;
  wire [15:0] t1_r6_c11_rr7;
  wire [15:0] t2_r6_c11_rr0;
  wire [15:0] t2_r6_c11_rr1;
  wire [15:0] t2_r6_c11_rr2;
  wire [15:0] t2_r6_c11_rr3;
  wire [15:0] t3_r6_c11_rr0;
  wire [15:0] t3_r6_c11_rr1;
  wire [15:0] t4_r6_c11_rr0;
  wire [15:0] t0_r6_c12_rr0;
  wire [15:0] t0_r6_c12_rr1;
  wire [15:0] t0_r6_c12_rr2;
  wire [15:0] t0_r6_c12_rr3;
  wire [15:0] t0_r6_c12_rr4;
  wire [15:0] t0_r6_c12_rr5;
  wire [15:0] t0_r6_c12_rr6;
  wire [15:0] t0_r6_c12_rr7;
  wire [15:0] t0_r6_c12_rr8;
  wire [15:0] t0_r6_c12_rr9;
  wire [15:0] t0_r6_c12_rr10;
  wire [15:0] t0_r6_c12_rr11;
  wire [15:0] t0_r6_c12_rr12;
  wire [15:0] t0_r6_c12_rr13;
  wire [15:0] t0_r6_c12_rr14;
  wire [15:0] t1_r6_c12_rr0;
  wire [15:0] t1_r6_c12_rr1;
  wire [15:0] t1_r6_c12_rr2;
  wire [15:0] t1_r6_c12_rr3;
  wire [15:0] t1_r6_c12_rr4;
  wire [15:0] t1_r6_c12_rr5;
  wire [15:0] t1_r6_c12_rr6;
  wire [15:0] t1_r6_c12_rr7;
  wire [15:0] t2_r6_c12_rr0;
  wire [15:0] t2_r6_c12_rr1;
  wire [15:0] t2_r6_c12_rr2;
  wire [15:0] t2_r6_c12_rr3;
  wire [15:0] t3_r6_c12_rr0;
  wire [15:0] t3_r6_c12_rr1;
  wire [15:0] t4_r6_c12_rr0;
  wire [15:0] t0_r6_c13_rr0;
  wire [15:0] t0_r6_c13_rr1;
  wire [15:0] t0_r6_c13_rr2;
  wire [15:0] t0_r6_c13_rr3;
  wire [15:0] t0_r6_c13_rr4;
  wire [15:0] t0_r6_c13_rr5;
  wire [15:0] t0_r6_c13_rr6;
  wire [15:0] t0_r6_c13_rr7;
  wire [15:0] t0_r6_c13_rr8;
  wire [15:0] t0_r6_c13_rr9;
  wire [15:0] t0_r6_c13_rr10;
  wire [15:0] t0_r6_c13_rr11;
  wire [15:0] t0_r6_c13_rr12;
  wire [15:0] t0_r6_c13_rr13;
  wire [15:0] t0_r6_c13_rr14;
  wire [15:0] t1_r6_c13_rr0;
  wire [15:0] t1_r6_c13_rr1;
  wire [15:0] t1_r6_c13_rr2;
  wire [15:0] t1_r6_c13_rr3;
  wire [15:0] t1_r6_c13_rr4;
  wire [15:0] t1_r6_c13_rr5;
  wire [15:0] t1_r6_c13_rr6;
  wire [15:0] t1_r6_c13_rr7;
  wire [15:0] t2_r6_c13_rr0;
  wire [15:0] t2_r6_c13_rr1;
  wire [15:0] t2_r6_c13_rr2;
  wire [15:0] t2_r6_c13_rr3;
  wire [15:0] t3_r6_c13_rr0;
  wire [15:0] t3_r6_c13_rr1;
  wire [15:0] t4_r6_c13_rr0;
  wire [15:0] t0_r6_c14_rr0;
  wire [15:0] t0_r6_c14_rr1;
  wire [15:0] t0_r6_c14_rr2;
  wire [15:0] t0_r6_c14_rr3;
  wire [15:0] t0_r6_c14_rr4;
  wire [15:0] t0_r6_c14_rr5;
  wire [15:0] t0_r6_c14_rr6;
  wire [15:0] t0_r6_c14_rr7;
  wire [15:0] t0_r6_c14_rr8;
  wire [15:0] t0_r6_c14_rr9;
  wire [15:0] t0_r6_c14_rr10;
  wire [15:0] t0_r6_c14_rr11;
  wire [15:0] t0_r6_c14_rr12;
  wire [15:0] t0_r6_c14_rr13;
  wire [15:0] t0_r6_c14_rr14;
  wire [15:0] t1_r6_c14_rr0;
  wire [15:0] t1_r6_c14_rr1;
  wire [15:0] t1_r6_c14_rr2;
  wire [15:0] t1_r6_c14_rr3;
  wire [15:0] t1_r6_c14_rr4;
  wire [15:0] t1_r6_c14_rr5;
  wire [15:0] t1_r6_c14_rr6;
  wire [15:0] t1_r6_c14_rr7;
  wire [15:0] t2_r6_c14_rr0;
  wire [15:0] t2_r6_c14_rr1;
  wire [15:0] t2_r6_c14_rr2;
  wire [15:0] t2_r6_c14_rr3;
  wire [15:0] t3_r6_c14_rr0;
  wire [15:0] t3_r6_c14_rr1;
  wire [15:0] t4_r6_c14_rr0;
  wire [15:0] t0_r7_c0_rr0;
  wire [15:0] t0_r7_c0_rr1;
  wire [15:0] t0_r7_c0_rr2;
  wire [15:0] t0_r7_c0_rr3;
  wire [15:0] t0_r7_c0_rr4;
  wire [15:0] t0_r7_c0_rr5;
  wire [15:0] t0_r7_c0_rr6;
  wire [15:0] t0_r7_c0_rr7;
  wire [15:0] t0_r7_c0_rr8;
  wire [15:0] t0_r7_c0_rr9;
  wire [15:0] t0_r7_c0_rr10;
  wire [15:0] t0_r7_c0_rr11;
  wire [15:0] t0_r7_c0_rr12;
  wire [15:0] t0_r7_c0_rr13;
  wire [15:0] t0_r7_c0_rr14;
  wire [15:0] t1_r7_c0_rr0;
  wire [15:0] t1_r7_c0_rr1;
  wire [15:0] t1_r7_c0_rr2;
  wire [15:0] t1_r7_c0_rr3;
  wire [15:0] t1_r7_c0_rr4;
  wire [15:0] t1_r7_c0_rr5;
  wire [15:0] t1_r7_c0_rr6;
  wire [15:0] t1_r7_c0_rr7;
  wire [15:0] t2_r7_c0_rr0;
  wire [15:0] t2_r7_c0_rr1;
  wire [15:0] t2_r7_c0_rr2;
  wire [15:0] t2_r7_c0_rr3;
  wire [15:0] t3_r7_c0_rr0;
  wire [15:0] t3_r7_c0_rr1;
  wire [15:0] t4_r7_c0_rr0;
  wire [15:0] t0_r7_c1_rr0;
  wire [15:0] t0_r7_c1_rr1;
  wire [15:0] t0_r7_c1_rr2;
  wire [15:0] t0_r7_c1_rr3;
  wire [15:0] t0_r7_c1_rr4;
  wire [15:0] t0_r7_c1_rr5;
  wire [15:0] t0_r7_c1_rr6;
  wire [15:0] t0_r7_c1_rr7;
  wire [15:0] t0_r7_c1_rr8;
  wire [15:0] t0_r7_c1_rr9;
  wire [15:0] t0_r7_c1_rr10;
  wire [15:0] t0_r7_c1_rr11;
  wire [15:0] t0_r7_c1_rr12;
  wire [15:0] t0_r7_c1_rr13;
  wire [15:0] t0_r7_c1_rr14;
  wire [15:0] t1_r7_c1_rr0;
  wire [15:0] t1_r7_c1_rr1;
  wire [15:0] t1_r7_c1_rr2;
  wire [15:0] t1_r7_c1_rr3;
  wire [15:0] t1_r7_c1_rr4;
  wire [15:0] t1_r7_c1_rr5;
  wire [15:0] t1_r7_c1_rr6;
  wire [15:0] t1_r7_c1_rr7;
  wire [15:0] t2_r7_c1_rr0;
  wire [15:0] t2_r7_c1_rr1;
  wire [15:0] t2_r7_c1_rr2;
  wire [15:0] t2_r7_c1_rr3;
  wire [15:0] t3_r7_c1_rr0;
  wire [15:0] t3_r7_c1_rr1;
  wire [15:0] t4_r7_c1_rr0;
  wire [15:0] t0_r7_c2_rr0;
  wire [15:0] t0_r7_c2_rr1;
  wire [15:0] t0_r7_c2_rr2;
  wire [15:0] t0_r7_c2_rr3;
  wire [15:0] t0_r7_c2_rr4;
  wire [15:0] t0_r7_c2_rr5;
  wire [15:0] t0_r7_c2_rr6;
  wire [15:0] t0_r7_c2_rr7;
  wire [15:0] t0_r7_c2_rr8;
  wire [15:0] t0_r7_c2_rr9;
  wire [15:0] t0_r7_c2_rr10;
  wire [15:0] t0_r7_c2_rr11;
  wire [15:0] t0_r7_c2_rr12;
  wire [15:0] t0_r7_c2_rr13;
  wire [15:0] t0_r7_c2_rr14;
  wire [15:0] t1_r7_c2_rr0;
  wire [15:0] t1_r7_c2_rr1;
  wire [15:0] t1_r7_c2_rr2;
  wire [15:0] t1_r7_c2_rr3;
  wire [15:0] t1_r7_c2_rr4;
  wire [15:0] t1_r7_c2_rr5;
  wire [15:0] t1_r7_c2_rr6;
  wire [15:0] t1_r7_c2_rr7;
  wire [15:0] t2_r7_c2_rr0;
  wire [15:0] t2_r7_c2_rr1;
  wire [15:0] t2_r7_c2_rr2;
  wire [15:0] t2_r7_c2_rr3;
  wire [15:0] t3_r7_c2_rr0;
  wire [15:0] t3_r7_c2_rr1;
  wire [15:0] t4_r7_c2_rr0;
  wire [15:0] t0_r7_c3_rr0;
  wire [15:0] t0_r7_c3_rr1;
  wire [15:0] t0_r7_c3_rr2;
  wire [15:0] t0_r7_c3_rr3;
  wire [15:0] t0_r7_c3_rr4;
  wire [15:0] t0_r7_c3_rr5;
  wire [15:0] t0_r7_c3_rr6;
  wire [15:0] t0_r7_c3_rr7;
  wire [15:0] t0_r7_c3_rr8;
  wire [15:0] t0_r7_c3_rr9;
  wire [15:0] t0_r7_c3_rr10;
  wire [15:0] t0_r7_c3_rr11;
  wire [15:0] t0_r7_c3_rr12;
  wire [15:0] t0_r7_c3_rr13;
  wire [15:0] t0_r7_c3_rr14;
  wire [15:0] t1_r7_c3_rr0;
  wire [15:0] t1_r7_c3_rr1;
  wire [15:0] t1_r7_c3_rr2;
  wire [15:0] t1_r7_c3_rr3;
  wire [15:0] t1_r7_c3_rr4;
  wire [15:0] t1_r7_c3_rr5;
  wire [15:0] t1_r7_c3_rr6;
  wire [15:0] t1_r7_c3_rr7;
  wire [15:0] t2_r7_c3_rr0;
  wire [15:0] t2_r7_c3_rr1;
  wire [15:0] t2_r7_c3_rr2;
  wire [15:0] t2_r7_c3_rr3;
  wire [15:0] t3_r7_c3_rr0;
  wire [15:0] t3_r7_c3_rr1;
  wire [15:0] t4_r7_c3_rr0;
  wire [15:0] t0_r7_c4_rr0;
  wire [15:0] t0_r7_c4_rr1;
  wire [15:0] t0_r7_c4_rr2;
  wire [15:0] t0_r7_c4_rr3;
  wire [15:0] t0_r7_c4_rr4;
  wire [15:0] t0_r7_c4_rr5;
  wire [15:0] t0_r7_c4_rr6;
  wire [15:0] t0_r7_c4_rr7;
  wire [15:0] t0_r7_c4_rr8;
  wire [15:0] t0_r7_c4_rr9;
  wire [15:0] t0_r7_c4_rr10;
  wire [15:0] t0_r7_c4_rr11;
  wire [15:0] t0_r7_c4_rr12;
  wire [15:0] t0_r7_c4_rr13;
  wire [15:0] t0_r7_c4_rr14;
  wire [15:0] t1_r7_c4_rr0;
  wire [15:0] t1_r7_c4_rr1;
  wire [15:0] t1_r7_c4_rr2;
  wire [15:0] t1_r7_c4_rr3;
  wire [15:0] t1_r7_c4_rr4;
  wire [15:0] t1_r7_c4_rr5;
  wire [15:0] t1_r7_c4_rr6;
  wire [15:0] t1_r7_c4_rr7;
  wire [15:0] t2_r7_c4_rr0;
  wire [15:0] t2_r7_c4_rr1;
  wire [15:0] t2_r7_c4_rr2;
  wire [15:0] t2_r7_c4_rr3;
  wire [15:0] t3_r7_c4_rr0;
  wire [15:0] t3_r7_c4_rr1;
  wire [15:0] t4_r7_c4_rr0;
  wire [15:0] t0_r7_c5_rr0;
  wire [15:0] t0_r7_c5_rr1;
  wire [15:0] t0_r7_c5_rr2;
  wire [15:0] t0_r7_c5_rr3;
  wire [15:0] t0_r7_c5_rr4;
  wire [15:0] t0_r7_c5_rr5;
  wire [15:0] t0_r7_c5_rr6;
  wire [15:0] t0_r7_c5_rr7;
  wire [15:0] t0_r7_c5_rr8;
  wire [15:0] t0_r7_c5_rr9;
  wire [15:0] t0_r7_c5_rr10;
  wire [15:0] t0_r7_c5_rr11;
  wire [15:0] t0_r7_c5_rr12;
  wire [15:0] t0_r7_c5_rr13;
  wire [15:0] t0_r7_c5_rr14;
  wire [15:0] t1_r7_c5_rr0;
  wire [15:0] t1_r7_c5_rr1;
  wire [15:0] t1_r7_c5_rr2;
  wire [15:0] t1_r7_c5_rr3;
  wire [15:0] t1_r7_c5_rr4;
  wire [15:0] t1_r7_c5_rr5;
  wire [15:0] t1_r7_c5_rr6;
  wire [15:0] t1_r7_c5_rr7;
  wire [15:0] t2_r7_c5_rr0;
  wire [15:0] t2_r7_c5_rr1;
  wire [15:0] t2_r7_c5_rr2;
  wire [15:0] t2_r7_c5_rr3;
  wire [15:0] t3_r7_c5_rr0;
  wire [15:0] t3_r7_c5_rr1;
  wire [15:0] t4_r7_c5_rr0;
  wire [15:0] t0_r7_c6_rr0;
  wire [15:0] t0_r7_c6_rr1;
  wire [15:0] t0_r7_c6_rr2;
  wire [15:0] t0_r7_c6_rr3;
  wire [15:0] t0_r7_c6_rr4;
  wire [15:0] t0_r7_c6_rr5;
  wire [15:0] t0_r7_c6_rr6;
  wire [15:0] t0_r7_c6_rr7;
  wire [15:0] t0_r7_c6_rr8;
  wire [15:0] t0_r7_c6_rr9;
  wire [15:0] t0_r7_c6_rr10;
  wire [15:0] t0_r7_c6_rr11;
  wire [15:0] t0_r7_c6_rr12;
  wire [15:0] t0_r7_c6_rr13;
  wire [15:0] t0_r7_c6_rr14;
  wire [15:0] t1_r7_c6_rr0;
  wire [15:0] t1_r7_c6_rr1;
  wire [15:0] t1_r7_c6_rr2;
  wire [15:0] t1_r7_c6_rr3;
  wire [15:0] t1_r7_c6_rr4;
  wire [15:0] t1_r7_c6_rr5;
  wire [15:0] t1_r7_c6_rr6;
  wire [15:0] t1_r7_c6_rr7;
  wire [15:0] t2_r7_c6_rr0;
  wire [15:0] t2_r7_c6_rr1;
  wire [15:0] t2_r7_c6_rr2;
  wire [15:0] t2_r7_c6_rr3;
  wire [15:0] t3_r7_c6_rr0;
  wire [15:0] t3_r7_c6_rr1;
  wire [15:0] t4_r7_c6_rr0;
  wire [15:0] t0_r7_c7_rr0;
  wire [15:0] t0_r7_c7_rr1;
  wire [15:0] t0_r7_c7_rr2;
  wire [15:0] t0_r7_c7_rr3;
  wire [15:0] t0_r7_c7_rr4;
  wire [15:0] t0_r7_c7_rr5;
  wire [15:0] t0_r7_c7_rr6;
  wire [15:0] t0_r7_c7_rr7;
  wire [15:0] t0_r7_c7_rr8;
  wire [15:0] t0_r7_c7_rr9;
  wire [15:0] t0_r7_c7_rr10;
  wire [15:0] t0_r7_c7_rr11;
  wire [15:0] t0_r7_c7_rr12;
  wire [15:0] t0_r7_c7_rr13;
  wire [15:0] t0_r7_c7_rr14;
  wire [15:0] t1_r7_c7_rr0;
  wire [15:0] t1_r7_c7_rr1;
  wire [15:0] t1_r7_c7_rr2;
  wire [15:0] t1_r7_c7_rr3;
  wire [15:0] t1_r7_c7_rr4;
  wire [15:0] t1_r7_c7_rr5;
  wire [15:0] t1_r7_c7_rr6;
  wire [15:0] t1_r7_c7_rr7;
  wire [15:0] t2_r7_c7_rr0;
  wire [15:0] t2_r7_c7_rr1;
  wire [15:0] t2_r7_c7_rr2;
  wire [15:0] t2_r7_c7_rr3;
  wire [15:0] t3_r7_c7_rr0;
  wire [15:0] t3_r7_c7_rr1;
  wire [15:0] t4_r7_c7_rr0;
  wire [15:0] t0_r7_c8_rr0;
  wire [15:0] t0_r7_c8_rr1;
  wire [15:0] t0_r7_c8_rr2;
  wire [15:0] t0_r7_c8_rr3;
  wire [15:0] t0_r7_c8_rr4;
  wire [15:0] t0_r7_c8_rr5;
  wire [15:0] t0_r7_c8_rr6;
  wire [15:0] t0_r7_c8_rr7;
  wire [15:0] t0_r7_c8_rr8;
  wire [15:0] t0_r7_c8_rr9;
  wire [15:0] t0_r7_c8_rr10;
  wire [15:0] t0_r7_c8_rr11;
  wire [15:0] t0_r7_c8_rr12;
  wire [15:0] t0_r7_c8_rr13;
  wire [15:0] t0_r7_c8_rr14;
  wire [15:0] t1_r7_c8_rr0;
  wire [15:0] t1_r7_c8_rr1;
  wire [15:0] t1_r7_c8_rr2;
  wire [15:0] t1_r7_c8_rr3;
  wire [15:0] t1_r7_c8_rr4;
  wire [15:0] t1_r7_c8_rr5;
  wire [15:0] t1_r7_c8_rr6;
  wire [15:0] t1_r7_c8_rr7;
  wire [15:0] t2_r7_c8_rr0;
  wire [15:0] t2_r7_c8_rr1;
  wire [15:0] t2_r7_c8_rr2;
  wire [15:0] t2_r7_c8_rr3;
  wire [15:0] t3_r7_c8_rr0;
  wire [15:0] t3_r7_c8_rr1;
  wire [15:0] t4_r7_c8_rr0;
  wire [15:0] t0_r7_c9_rr0;
  wire [15:0] t0_r7_c9_rr1;
  wire [15:0] t0_r7_c9_rr2;
  wire [15:0] t0_r7_c9_rr3;
  wire [15:0] t0_r7_c9_rr4;
  wire [15:0] t0_r7_c9_rr5;
  wire [15:0] t0_r7_c9_rr6;
  wire [15:0] t0_r7_c9_rr7;
  wire [15:0] t0_r7_c9_rr8;
  wire [15:0] t0_r7_c9_rr9;
  wire [15:0] t0_r7_c9_rr10;
  wire [15:0] t0_r7_c9_rr11;
  wire [15:0] t0_r7_c9_rr12;
  wire [15:0] t0_r7_c9_rr13;
  wire [15:0] t0_r7_c9_rr14;
  wire [15:0] t1_r7_c9_rr0;
  wire [15:0] t1_r7_c9_rr1;
  wire [15:0] t1_r7_c9_rr2;
  wire [15:0] t1_r7_c9_rr3;
  wire [15:0] t1_r7_c9_rr4;
  wire [15:0] t1_r7_c9_rr5;
  wire [15:0] t1_r7_c9_rr6;
  wire [15:0] t1_r7_c9_rr7;
  wire [15:0] t2_r7_c9_rr0;
  wire [15:0] t2_r7_c9_rr1;
  wire [15:0] t2_r7_c9_rr2;
  wire [15:0] t2_r7_c9_rr3;
  wire [15:0] t3_r7_c9_rr0;
  wire [15:0] t3_r7_c9_rr1;
  wire [15:0] t4_r7_c9_rr0;
  wire [15:0] t0_r7_c10_rr0;
  wire [15:0] t0_r7_c10_rr1;
  wire [15:0] t0_r7_c10_rr2;
  wire [15:0] t0_r7_c10_rr3;
  wire [15:0] t0_r7_c10_rr4;
  wire [15:0] t0_r7_c10_rr5;
  wire [15:0] t0_r7_c10_rr6;
  wire [15:0] t0_r7_c10_rr7;
  wire [15:0] t0_r7_c10_rr8;
  wire [15:0] t0_r7_c10_rr9;
  wire [15:0] t0_r7_c10_rr10;
  wire [15:0] t0_r7_c10_rr11;
  wire [15:0] t0_r7_c10_rr12;
  wire [15:0] t0_r7_c10_rr13;
  wire [15:0] t0_r7_c10_rr14;
  wire [15:0] t1_r7_c10_rr0;
  wire [15:0] t1_r7_c10_rr1;
  wire [15:0] t1_r7_c10_rr2;
  wire [15:0] t1_r7_c10_rr3;
  wire [15:0] t1_r7_c10_rr4;
  wire [15:0] t1_r7_c10_rr5;
  wire [15:0] t1_r7_c10_rr6;
  wire [15:0] t1_r7_c10_rr7;
  wire [15:0] t2_r7_c10_rr0;
  wire [15:0] t2_r7_c10_rr1;
  wire [15:0] t2_r7_c10_rr2;
  wire [15:0] t2_r7_c10_rr3;
  wire [15:0] t3_r7_c10_rr0;
  wire [15:0] t3_r7_c10_rr1;
  wire [15:0] t4_r7_c10_rr0;
  wire [15:0] t0_r7_c11_rr0;
  wire [15:0] t0_r7_c11_rr1;
  wire [15:0] t0_r7_c11_rr2;
  wire [15:0] t0_r7_c11_rr3;
  wire [15:0] t0_r7_c11_rr4;
  wire [15:0] t0_r7_c11_rr5;
  wire [15:0] t0_r7_c11_rr6;
  wire [15:0] t0_r7_c11_rr7;
  wire [15:0] t0_r7_c11_rr8;
  wire [15:0] t0_r7_c11_rr9;
  wire [15:0] t0_r7_c11_rr10;
  wire [15:0] t0_r7_c11_rr11;
  wire [15:0] t0_r7_c11_rr12;
  wire [15:0] t0_r7_c11_rr13;
  wire [15:0] t0_r7_c11_rr14;
  wire [15:0] t1_r7_c11_rr0;
  wire [15:0] t1_r7_c11_rr1;
  wire [15:0] t1_r7_c11_rr2;
  wire [15:0] t1_r7_c11_rr3;
  wire [15:0] t1_r7_c11_rr4;
  wire [15:0] t1_r7_c11_rr5;
  wire [15:0] t1_r7_c11_rr6;
  wire [15:0] t1_r7_c11_rr7;
  wire [15:0] t2_r7_c11_rr0;
  wire [15:0] t2_r7_c11_rr1;
  wire [15:0] t2_r7_c11_rr2;
  wire [15:0] t2_r7_c11_rr3;
  wire [15:0] t3_r7_c11_rr0;
  wire [15:0] t3_r7_c11_rr1;
  wire [15:0] t4_r7_c11_rr0;
  wire [15:0] t0_r7_c12_rr0;
  wire [15:0] t0_r7_c12_rr1;
  wire [15:0] t0_r7_c12_rr2;
  wire [15:0] t0_r7_c12_rr3;
  wire [15:0] t0_r7_c12_rr4;
  wire [15:0] t0_r7_c12_rr5;
  wire [15:0] t0_r7_c12_rr6;
  wire [15:0] t0_r7_c12_rr7;
  wire [15:0] t0_r7_c12_rr8;
  wire [15:0] t0_r7_c12_rr9;
  wire [15:0] t0_r7_c12_rr10;
  wire [15:0] t0_r7_c12_rr11;
  wire [15:0] t0_r7_c12_rr12;
  wire [15:0] t0_r7_c12_rr13;
  wire [15:0] t0_r7_c12_rr14;
  wire [15:0] t1_r7_c12_rr0;
  wire [15:0] t1_r7_c12_rr1;
  wire [15:0] t1_r7_c12_rr2;
  wire [15:0] t1_r7_c12_rr3;
  wire [15:0] t1_r7_c12_rr4;
  wire [15:0] t1_r7_c12_rr5;
  wire [15:0] t1_r7_c12_rr6;
  wire [15:0] t1_r7_c12_rr7;
  wire [15:0] t2_r7_c12_rr0;
  wire [15:0] t2_r7_c12_rr1;
  wire [15:0] t2_r7_c12_rr2;
  wire [15:0] t2_r7_c12_rr3;
  wire [15:0] t3_r7_c12_rr0;
  wire [15:0] t3_r7_c12_rr1;
  wire [15:0] t4_r7_c12_rr0;
  wire [15:0] t0_r7_c13_rr0;
  wire [15:0] t0_r7_c13_rr1;
  wire [15:0] t0_r7_c13_rr2;
  wire [15:0] t0_r7_c13_rr3;
  wire [15:0] t0_r7_c13_rr4;
  wire [15:0] t0_r7_c13_rr5;
  wire [15:0] t0_r7_c13_rr6;
  wire [15:0] t0_r7_c13_rr7;
  wire [15:0] t0_r7_c13_rr8;
  wire [15:0] t0_r7_c13_rr9;
  wire [15:0] t0_r7_c13_rr10;
  wire [15:0] t0_r7_c13_rr11;
  wire [15:0] t0_r7_c13_rr12;
  wire [15:0] t0_r7_c13_rr13;
  wire [15:0] t0_r7_c13_rr14;
  wire [15:0] t1_r7_c13_rr0;
  wire [15:0] t1_r7_c13_rr1;
  wire [15:0] t1_r7_c13_rr2;
  wire [15:0] t1_r7_c13_rr3;
  wire [15:0] t1_r7_c13_rr4;
  wire [15:0] t1_r7_c13_rr5;
  wire [15:0] t1_r7_c13_rr6;
  wire [15:0] t1_r7_c13_rr7;
  wire [15:0] t2_r7_c13_rr0;
  wire [15:0] t2_r7_c13_rr1;
  wire [15:0] t2_r7_c13_rr2;
  wire [15:0] t2_r7_c13_rr3;
  wire [15:0] t3_r7_c13_rr0;
  wire [15:0] t3_r7_c13_rr1;
  wire [15:0] t4_r7_c13_rr0;
  wire [15:0] t0_r7_c14_rr0;
  wire [15:0] t0_r7_c14_rr1;
  wire [15:0] t0_r7_c14_rr2;
  wire [15:0] t0_r7_c14_rr3;
  wire [15:0] t0_r7_c14_rr4;
  wire [15:0] t0_r7_c14_rr5;
  wire [15:0] t0_r7_c14_rr6;
  wire [15:0] t0_r7_c14_rr7;
  wire [15:0] t0_r7_c14_rr8;
  wire [15:0] t0_r7_c14_rr9;
  wire [15:0] t0_r7_c14_rr10;
  wire [15:0] t0_r7_c14_rr11;
  wire [15:0] t0_r7_c14_rr12;
  wire [15:0] t0_r7_c14_rr13;
  wire [15:0] t0_r7_c14_rr14;
  wire [15:0] t1_r7_c14_rr0;
  wire [15:0] t1_r7_c14_rr1;
  wire [15:0] t1_r7_c14_rr2;
  wire [15:0] t1_r7_c14_rr3;
  wire [15:0] t1_r7_c14_rr4;
  wire [15:0] t1_r7_c14_rr5;
  wire [15:0] t1_r7_c14_rr6;
  wire [15:0] t1_r7_c14_rr7;
  wire [15:0] t2_r7_c14_rr0;
  wire [15:0] t2_r7_c14_rr1;
  wire [15:0] t2_r7_c14_rr2;
  wire [15:0] t2_r7_c14_rr3;
  wire [15:0] t3_r7_c14_rr0;
  wire [15:0] t3_r7_c14_rr1;
  wire [15:0] t4_r7_c14_rr0;
  wire [15:0] t0_r8_c0_rr0;
  wire [15:0] t0_r8_c0_rr1;
  wire [15:0] t0_r8_c0_rr2;
  wire [15:0] t0_r8_c0_rr3;
  wire [15:0] t0_r8_c0_rr4;
  wire [15:0] t0_r8_c0_rr5;
  wire [15:0] t0_r8_c0_rr6;
  wire [15:0] t0_r8_c0_rr7;
  wire [15:0] t0_r8_c0_rr8;
  wire [15:0] t0_r8_c0_rr9;
  wire [15:0] t0_r8_c0_rr10;
  wire [15:0] t0_r8_c0_rr11;
  wire [15:0] t0_r8_c0_rr12;
  wire [15:0] t0_r8_c0_rr13;
  wire [15:0] t0_r8_c0_rr14;
  wire [15:0] t1_r8_c0_rr0;
  wire [15:0] t1_r8_c0_rr1;
  wire [15:0] t1_r8_c0_rr2;
  wire [15:0] t1_r8_c0_rr3;
  wire [15:0] t1_r8_c0_rr4;
  wire [15:0] t1_r8_c0_rr5;
  wire [15:0] t1_r8_c0_rr6;
  wire [15:0] t1_r8_c0_rr7;
  wire [15:0] t2_r8_c0_rr0;
  wire [15:0] t2_r8_c0_rr1;
  wire [15:0] t2_r8_c0_rr2;
  wire [15:0] t2_r8_c0_rr3;
  wire [15:0] t3_r8_c0_rr0;
  wire [15:0] t3_r8_c0_rr1;
  wire [15:0] t4_r8_c0_rr0;
  wire [15:0] t0_r8_c1_rr0;
  wire [15:0] t0_r8_c1_rr1;
  wire [15:0] t0_r8_c1_rr2;
  wire [15:0] t0_r8_c1_rr3;
  wire [15:0] t0_r8_c1_rr4;
  wire [15:0] t0_r8_c1_rr5;
  wire [15:0] t0_r8_c1_rr6;
  wire [15:0] t0_r8_c1_rr7;
  wire [15:0] t0_r8_c1_rr8;
  wire [15:0] t0_r8_c1_rr9;
  wire [15:0] t0_r8_c1_rr10;
  wire [15:0] t0_r8_c1_rr11;
  wire [15:0] t0_r8_c1_rr12;
  wire [15:0] t0_r8_c1_rr13;
  wire [15:0] t0_r8_c1_rr14;
  wire [15:0] t1_r8_c1_rr0;
  wire [15:0] t1_r8_c1_rr1;
  wire [15:0] t1_r8_c1_rr2;
  wire [15:0] t1_r8_c1_rr3;
  wire [15:0] t1_r8_c1_rr4;
  wire [15:0] t1_r8_c1_rr5;
  wire [15:0] t1_r8_c1_rr6;
  wire [15:0] t1_r8_c1_rr7;
  wire [15:0] t2_r8_c1_rr0;
  wire [15:0] t2_r8_c1_rr1;
  wire [15:0] t2_r8_c1_rr2;
  wire [15:0] t2_r8_c1_rr3;
  wire [15:0] t3_r8_c1_rr0;
  wire [15:0] t3_r8_c1_rr1;
  wire [15:0] t4_r8_c1_rr0;
  wire [15:0] t0_r8_c2_rr0;
  wire [15:0] t0_r8_c2_rr1;
  wire [15:0] t0_r8_c2_rr2;
  wire [15:0] t0_r8_c2_rr3;
  wire [15:0] t0_r8_c2_rr4;
  wire [15:0] t0_r8_c2_rr5;
  wire [15:0] t0_r8_c2_rr6;
  wire [15:0] t0_r8_c2_rr7;
  wire [15:0] t0_r8_c2_rr8;
  wire [15:0] t0_r8_c2_rr9;
  wire [15:0] t0_r8_c2_rr10;
  wire [15:0] t0_r8_c2_rr11;
  wire [15:0] t0_r8_c2_rr12;
  wire [15:0] t0_r8_c2_rr13;
  wire [15:0] t0_r8_c2_rr14;
  wire [15:0] t1_r8_c2_rr0;
  wire [15:0] t1_r8_c2_rr1;
  wire [15:0] t1_r8_c2_rr2;
  wire [15:0] t1_r8_c2_rr3;
  wire [15:0] t1_r8_c2_rr4;
  wire [15:0] t1_r8_c2_rr5;
  wire [15:0] t1_r8_c2_rr6;
  wire [15:0] t1_r8_c2_rr7;
  wire [15:0] t2_r8_c2_rr0;
  wire [15:0] t2_r8_c2_rr1;
  wire [15:0] t2_r8_c2_rr2;
  wire [15:0] t2_r8_c2_rr3;
  wire [15:0] t3_r8_c2_rr0;
  wire [15:0] t3_r8_c2_rr1;
  wire [15:0] t4_r8_c2_rr0;
  wire [15:0] t0_r8_c3_rr0;
  wire [15:0] t0_r8_c3_rr1;
  wire [15:0] t0_r8_c3_rr2;
  wire [15:0] t0_r8_c3_rr3;
  wire [15:0] t0_r8_c3_rr4;
  wire [15:0] t0_r8_c3_rr5;
  wire [15:0] t0_r8_c3_rr6;
  wire [15:0] t0_r8_c3_rr7;
  wire [15:0] t0_r8_c3_rr8;
  wire [15:0] t0_r8_c3_rr9;
  wire [15:0] t0_r8_c3_rr10;
  wire [15:0] t0_r8_c3_rr11;
  wire [15:0] t0_r8_c3_rr12;
  wire [15:0] t0_r8_c3_rr13;
  wire [15:0] t0_r8_c3_rr14;
  wire [15:0] t1_r8_c3_rr0;
  wire [15:0] t1_r8_c3_rr1;
  wire [15:0] t1_r8_c3_rr2;
  wire [15:0] t1_r8_c3_rr3;
  wire [15:0] t1_r8_c3_rr4;
  wire [15:0] t1_r8_c3_rr5;
  wire [15:0] t1_r8_c3_rr6;
  wire [15:0] t1_r8_c3_rr7;
  wire [15:0] t2_r8_c3_rr0;
  wire [15:0] t2_r8_c3_rr1;
  wire [15:0] t2_r8_c3_rr2;
  wire [15:0] t2_r8_c3_rr3;
  wire [15:0] t3_r8_c3_rr0;
  wire [15:0] t3_r8_c3_rr1;
  wire [15:0] t4_r8_c3_rr0;
  wire [15:0] t0_r8_c4_rr0;
  wire [15:0] t0_r8_c4_rr1;
  wire [15:0] t0_r8_c4_rr2;
  wire [15:0] t0_r8_c4_rr3;
  wire [15:0] t0_r8_c4_rr4;
  wire [15:0] t0_r8_c4_rr5;
  wire [15:0] t0_r8_c4_rr6;
  wire [15:0] t0_r8_c4_rr7;
  wire [15:0] t0_r8_c4_rr8;
  wire [15:0] t0_r8_c4_rr9;
  wire [15:0] t0_r8_c4_rr10;
  wire [15:0] t0_r8_c4_rr11;
  wire [15:0] t0_r8_c4_rr12;
  wire [15:0] t0_r8_c4_rr13;
  wire [15:0] t0_r8_c4_rr14;
  wire [15:0] t1_r8_c4_rr0;
  wire [15:0] t1_r8_c4_rr1;
  wire [15:0] t1_r8_c4_rr2;
  wire [15:0] t1_r8_c4_rr3;
  wire [15:0] t1_r8_c4_rr4;
  wire [15:0] t1_r8_c4_rr5;
  wire [15:0] t1_r8_c4_rr6;
  wire [15:0] t1_r8_c4_rr7;
  wire [15:0] t2_r8_c4_rr0;
  wire [15:0] t2_r8_c4_rr1;
  wire [15:0] t2_r8_c4_rr2;
  wire [15:0] t2_r8_c4_rr3;
  wire [15:0] t3_r8_c4_rr0;
  wire [15:0] t3_r8_c4_rr1;
  wire [15:0] t4_r8_c4_rr0;
  wire [15:0] t0_r8_c5_rr0;
  wire [15:0] t0_r8_c5_rr1;
  wire [15:0] t0_r8_c5_rr2;
  wire [15:0] t0_r8_c5_rr3;
  wire [15:0] t0_r8_c5_rr4;
  wire [15:0] t0_r8_c5_rr5;
  wire [15:0] t0_r8_c5_rr6;
  wire [15:0] t0_r8_c5_rr7;
  wire [15:0] t0_r8_c5_rr8;
  wire [15:0] t0_r8_c5_rr9;
  wire [15:0] t0_r8_c5_rr10;
  wire [15:0] t0_r8_c5_rr11;
  wire [15:0] t0_r8_c5_rr12;
  wire [15:0] t0_r8_c5_rr13;
  wire [15:0] t0_r8_c5_rr14;
  wire [15:0] t1_r8_c5_rr0;
  wire [15:0] t1_r8_c5_rr1;
  wire [15:0] t1_r8_c5_rr2;
  wire [15:0] t1_r8_c5_rr3;
  wire [15:0] t1_r8_c5_rr4;
  wire [15:0] t1_r8_c5_rr5;
  wire [15:0] t1_r8_c5_rr6;
  wire [15:0] t1_r8_c5_rr7;
  wire [15:0] t2_r8_c5_rr0;
  wire [15:0] t2_r8_c5_rr1;
  wire [15:0] t2_r8_c5_rr2;
  wire [15:0] t2_r8_c5_rr3;
  wire [15:0] t3_r8_c5_rr0;
  wire [15:0] t3_r8_c5_rr1;
  wire [15:0] t4_r8_c5_rr0;
  wire [15:0] t0_r8_c6_rr0;
  wire [15:0] t0_r8_c6_rr1;
  wire [15:0] t0_r8_c6_rr2;
  wire [15:0] t0_r8_c6_rr3;
  wire [15:0] t0_r8_c6_rr4;
  wire [15:0] t0_r8_c6_rr5;
  wire [15:0] t0_r8_c6_rr6;
  wire [15:0] t0_r8_c6_rr7;
  wire [15:0] t0_r8_c6_rr8;
  wire [15:0] t0_r8_c6_rr9;
  wire [15:0] t0_r8_c6_rr10;
  wire [15:0] t0_r8_c6_rr11;
  wire [15:0] t0_r8_c6_rr12;
  wire [15:0] t0_r8_c6_rr13;
  wire [15:0] t0_r8_c6_rr14;
  wire [15:0] t1_r8_c6_rr0;
  wire [15:0] t1_r8_c6_rr1;
  wire [15:0] t1_r8_c6_rr2;
  wire [15:0] t1_r8_c6_rr3;
  wire [15:0] t1_r8_c6_rr4;
  wire [15:0] t1_r8_c6_rr5;
  wire [15:0] t1_r8_c6_rr6;
  wire [15:0] t1_r8_c6_rr7;
  wire [15:0] t2_r8_c6_rr0;
  wire [15:0] t2_r8_c6_rr1;
  wire [15:0] t2_r8_c6_rr2;
  wire [15:0] t2_r8_c6_rr3;
  wire [15:0] t3_r8_c6_rr0;
  wire [15:0] t3_r8_c6_rr1;
  wire [15:0] t4_r8_c6_rr0;
  wire [15:0] t0_r8_c7_rr0;
  wire [15:0] t0_r8_c7_rr1;
  wire [15:0] t0_r8_c7_rr2;
  wire [15:0] t0_r8_c7_rr3;
  wire [15:0] t0_r8_c7_rr4;
  wire [15:0] t0_r8_c7_rr5;
  wire [15:0] t0_r8_c7_rr6;
  wire [15:0] t0_r8_c7_rr7;
  wire [15:0] t0_r8_c7_rr8;
  wire [15:0] t0_r8_c7_rr9;
  wire [15:0] t0_r8_c7_rr10;
  wire [15:0] t0_r8_c7_rr11;
  wire [15:0] t0_r8_c7_rr12;
  wire [15:0] t0_r8_c7_rr13;
  wire [15:0] t0_r8_c7_rr14;
  wire [15:0] t1_r8_c7_rr0;
  wire [15:0] t1_r8_c7_rr1;
  wire [15:0] t1_r8_c7_rr2;
  wire [15:0] t1_r8_c7_rr3;
  wire [15:0] t1_r8_c7_rr4;
  wire [15:0] t1_r8_c7_rr5;
  wire [15:0] t1_r8_c7_rr6;
  wire [15:0] t1_r8_c7_rr7;
  wire [15:0] t2_r8_c7_rr0;
  wire [15:0] t2_r8_c7_rr1;
  wire [15:0] t2_r8_c7_rr2;
  wire [15:0] t2_r8_c7_rr3;
  wire [15:0] t3_r8_c7_rr0;
  wire [15:0] t3_r8_c7_rr1;
  wire [15:0] t4_r8_c7_rr0;
  wire [15:0] t0_r8_c8_rr0;
  wire [15:0] t0_r8_c8_rr1;
  wire [15:0] t0_r8_c8_rr2;
  wire [15:0] t0_r8_c8_rr3;
  wire [15:0] t0_r8_c8_rr4;
  wire [15:0] t0_r8_c8_rr5;
  wire [15:0] t0_r8_c8_rr6;
  wire [15:0] t0_r8_c8_rr7;
  wire [15:0] t0_r8_c8_rr8;
  wire [15:0] t0_r8_c8_rr9;
  wire [15:0] t0_r8_c8_rr10;
  wire [15:0] t0_r8_c8_rr11;
  wire [15:0] t0_r8_c8_rr12;
  wire [15:0] t0_r8_c8_rr13;
  wire [15:0] t0_r8_c8_rr14;
  wire [15:0] t1_r8_c8_rr0;
  wire [15:0] t1_r8_c8_rr1;
  wire [15:0] t1_r8_c8_rr2;
  wire [15:0] t1_r8_c8_rr3;
  wire [15:0] t1_r8_c8_rr4;
  wire [15:0] t1_r8_c8_rr5;
  wire [15:0] t1_r8_c8_rr6;
  wire [15:0] t1_r8_c8_rr7;
  wire [15:0] t2_r8_c8_rr0;
  wire [15:0] t2_r8_c8_rr1;
  wire [15:0] t2_r8_c8_rr2;
  wire [15:0] t2_r8_c8_rr3;
  wire [15:0] t3_r8_c8_rr0;
  wire [15:0] t3_r8_c8_rr1;
  wire [15:0] t4_r8_c8_rr0;
  wire [15:0] t0_r8_c9_rr0;
  wire [15:0] t0_r8_c9_rr1;
  wire [15:0] t0_r8_c9_rr2;
  wire [15:0] t0_r8_c9_rr3;
  wire [15:0] t0_r8_c9_rr4;
  wire [15:0] t0_r8_c9_rr5;
  wire [15:0] t0_r8_c9_rr6;
  wire [15:0] t0_r8_c9_rr7;
  wire [15:0] t0_r8_c9_rr8;
  wire [15:0] t0_r8_c9_rr9;
  wire [15:0] t0_r8_c9_rr10;
  wire [15:0] t0_r8_c9_rr11;
  wire [15:0] t0_r8_c9_rr12;
  wire [15:0] t0_r8_c9_rr13;
  wire [15:0] t0_r8_c9_rr14;
  wire [15:0] t1_r8_c9_rr0;
  wire [15:0] t1_r8_c9_rr1;
  wire [15:0] t1_r8_c9_rr2;
  wire [15:0] t1_r8_c9_rr3;
  wire [15:0] t1_r8_c9_rr4;
  wire [15:0] t1_r8_c9_rr5;
  wire [15:0] t1_r8_c9_rr6;
  wire [15:0] t1_r8_c9_rr7;
  wire [15:0] t2_r8_c9_rr0;
  wire [15:0] t2_r8_c9_rr1;
  wire [15:0] t2_r8_c9_rr2;
  wire [15:0] t2_r8_c9_rr3;
  wire [15:0] t3_r8_c9_rr0;
  wire [15:0] t3_r8_c9_rr1;
  wire [15:0] t4_r8_c9_rr0;
  wire [15:0] t0_r8_c10_rr0;
  wire [15:0] t0_r8_c10_rr1;
  wire [15:0] t0_r8_c10_rr2;
  wire [15:0] t0_r8_c10_rr3;
  wire [15:0] t0_r8_c10_rr4;
  wire [15:0] t0_r8_c10_rr5;
  wire [15:0] t0_r8_c10_rr6;
  wire [15:0] t0_r8_c10_rr7;
  wire [15:0] t0_r8_c10_rr8;
  wire [15:0] t0_r8_c10_rr9;
  wire [15:0] t0_r8_c10_rr10;
  wire [15:0] t0_r8_c10_rr11;
  wire [15:0] t0_r8_c10_rr12;
  wire [15:0] t0_r8_c10_rr13;
  wire [15:0] t0_r8_c10_rr14;
  wire [15:0] t1_r8_c10_rr0;
  wire [15:0] t1_r8_c10_rr1;
  wire [15:0] t1_r8_c10_rr2;
  wire [15:0] t1_r8_c10_rr3;
  wire [15:0] t1_r8_c10_rr4;
  wire [15:0] t1_r8_c10_rr5;
  wire [15:0] t1_r8_c10_rr6;
  wire [15:0] t1_r8_c10_rr7;
  wire [15:0] t2_r8_c10_rr0;
  wire [15:0] t2_r8_c10_rr1;
  wire [15:0] t2_r8_c10_rr2;
  wire [15:0] t2_r8_c10_rr3;
  wire [15:0] t3_r8_c10_rr0;
  wire [15:0] t3_r8_c10_rr1;
  wire [15:0] t4_r8_c10_rr0;
  wire [15:0] t0_r8_c11_rr0;
  wire [15:0] t0_r8_c11_rr1;
  wire [15:0] t0_r8_c11_rr2;
  wire [15:0] t0_r8_c11_rr3;
  wire [15:0] t0_r8_c11_rr4;
  wire [15:0] t0_r8_c11_rr5;
  wire [15:0] t0_r8_c11_rr6;
  wire [15:0] t0_r8_c11_rr7;
  wire [15:0] t0_r8_c11_rr8;
  wire [15:0] t0_r8_c11_rr9;
  wire [15:0] t0_r8_c11_rr10;
  wire [15:0] t0_r8_c11_rr11;
  wire [15:0] t0_r8_c11_rr12;
  wire [15:0] t0_r8_c11_rr13;
  wire [15:0] t0_r8_c11_rr14;
  wire [15:0] t1_r8_c11_rr0;
  wire [15:0] t1_r8_c11_rr1;
  wire [15:0] t1_r8_c11_rr2;
  wire [15:0] t1_r8_c11_rr3;
  wire [15:0] t1_r8_c11_rr4;
  wire [15:0] t1_r8_c11_rr5;
  wire [15:0] t1_r8_c11_rr6;
  wire [15:0] t1_r8_c11_rr7;
  wire [15:0] t2_r8_c11_rr0;
  wire [15:0] t2_r8_c11_rr1;
  wire [15:0] t2_r8_c11_rr2;
  wire [15:0] t2_r8_c11_rr3;
  wire [15:0] t3_r8_c11_rr0;
  wire [15:0] t3_r8_c11_rr1;
  wire [15:0] t4_r8_c11_rr0;
  wire [15:0] t0_r8_c12_rr0;
  wire [15:0] t0_r8_c12_rr1;
  wire [15:0] t0_r8_c12_rr2;
  wire [15:0] t0_r8_c12_rr3;
  wire [15:0] t0_r8_c12_rr4;
  wire [15:0] t0_r8_c12_rr5;
  wire [15:0] t0_r8_c12_rr6;
  wire [15:0] t0_r8_c12_rr7;
  wire [15:0] t0_r8_c12_rr8;
  wire [15:0] t0_r8_c12_rr9;
  wire [15:0] t0_r8_c12_rr10;
  wire [15:0] t0_r8_c12_rr11;
  wire [15:0] t0_r8_c12_rr12;
  wire [15:0] t0_r8_c12_rr13;
  wire [15:0] t0_r8_c12_rr14;
  wire [15:0] t1_r8_c12_rr0;
  wire [15:0] t1_r8_c12_rr1;
  wire [15:0] t1_r8_c12_rr2;
  wire [15:0] t1_r8_c12_rr3;
  wire [15:0] t1_r8_c12_rr4;
  wire [15:0] t1_r8_c12_rr5;
  wire [15:0] t1_r8_c12_rr6;
  wire [15:0] t1_r8_c12_rr7;
  wire [15:0] t2_r8_c12_rr0;
  wire [15:0] t2_r8_c12_rr1;
  wire [15:0] t2_r8_c12_rr2;
  wire [15:0] t2_r8_c12_rr3;
  wire [15:0] t3_r8_c12_rr0;
  wire [15:0] t3_r8_c12_rr1;
  wire [15:0] t4_r8_c12_rr0;
  wire [15:0] t0_r8_c13_rr0;
  wire [15:0] t0_r8_c13_rr1;
  wire [15:0] t0_r8_c13_rr2;
  wire [15:0] t0_r8_c13_rr3;
  wire [15:0] t0_r8_c13_rr4;
  wire [15:0] t0_r8_c13_rr5;
  wire [15:0] t0_r8_c13_rr6;
  wire [15:0] t0_r8_c13_rr7;
  wire [15:0] t0_r8_c13_rr8;
  wire [15:0] t0_r8_c13_rr9;
  wire [15:0] t0_r8_c13_rr10;
  wire [15:0] t0_r8_c13_rr11;
  wire [15:0] t0_r8_c13_rr12;
  wire [15:0] t0_r8_c13_rr13;
  wire [15:0] t0_r8_c13_rr14;
  wire [15:0] t1_r8_c13_rr0;
  wire [15:0] t1_r8_c13_rr1;
  wire [15:0] t1_r8_c13_rr2;
  wire [15:0] t1_r8_c13_rr3;
  wire [15:0] t1_r8_c13_rr4;
  wire [15:0] t1_r8_c13_rr5;
  wire [15:0] t1_r8_c13_rr6;
  wire [15:0] t1_r8_c13_rr7;
  wire [15:0] t2_r8_c13_rr0;
  wire [15:0] t2_r8_c13_rr1;
  wire [15:0] t2_r8_c13_rr2;
  wire [15:0] t2_r8_c13_rr3;
  wire [15:0] t3_r8_c13_rr0;
  wire [15:0] t3_r8_c13_rr1;
  wire [15:0] t4_r8_c13_rr0;
  wire [15:0] t0_r8_c14_rr0;
  wire [15:0] t0_r8_c14_rr1;
  wire [15:0] t0_r8_c14_rr2;
  wire [15:0] t0_r8_c14_rr3;
  wire [15:0] t0_r8_c14_rr4;
  wire [15:0] t0_r8_c14_rr5;
  wire [15:0] t0_r8_c14_rr6;
  wire [15:0] t0_r8_c14_rr7;
  wire [15:0] t0_r8_c14_rr8;
  wire [15:0] t0_r8_c14_rr9;
  wire [15:0] t0_r8_c14_rr10;
  wire [15:0] t0_r8_c14_rr11;
  wire [15:0] t0_r8_c14_rr12;
  wire [15:0] t0_r8_c14_rr13;
  wire [15:0] t0_r8_c14_rr14;
  wire [15:0] t1_r8_c14_rr0;
  wire [15:0] t1_r8_c14_rr1;
  wire [15:0] t1_r8_c14_rr2;
  wire [15:0] t1_r8_c14_rr3;
  wire [15:0] t1_r8_c14_rr4;
  wire [15:0] t1_r8_c14_rr5;
  wire [15:0] t1_r8_c14_rr6;
  wire [15:0] t1_r8_c14_rr7;
  wire [15:0] t2_r8_c14_rr0;
  wire [15:0] t2_r8_c14_rr1;
  wire [15:0] t2_r8_c14_rr2;
  wire [15:0] t2_r8_c14_rr3;
  wire [15:0] t3_r8_c14_rr0;
  wire [15:0] t3_r8_c14_rr1;
  wire [15:0] t4_r8_c14_rr0;
  wire [15:0] t0_r9_c0_rr0;
  wire [15:0] t0_r9_c0_rr1;
  wire [15:0] t0_r9_c0_rr2;
  wire [15:0] t0_r9_c0_rr3;
  wire [15:0] t0_r9_c0_rr4;
  wire [15:0] t0_r9_c0_rr5;
  wire [15:0] t0_r9_c0_rr6;
  wire [15:0] t0_r9_c0_rr7;
  wire [15:0] t0_r9_c0_rr8;
  wire [15:0] t0_r9_c0_rr9;
  wire [15:0] t0_r9_c0_rr10;
  wire [15:0] t0_r9_c0_rr11;
  wire [15:0] t0_r9_c0_rr12;
  wire [15:0] t0_r9_c0_rr13;
  wire [15:0] t0_r9_c0_rr14;
  wire [15:0] t1_r9_c0_rr0;
  wire [15:0] t1_r9_c0_rr1;
  wire [15:0] t1_r9_c0_rr2;
  wire [15:0] t1_r9_c0_rr3;
  wire [15:0] t1_r9_c0_rr4;
  wire [15:0] t1_r9_c0_rr5;
  wire [15:0] t1_r9_c0_rr6;
  wire [15:0] t1_r9_c0_rr7;
  wire [15:0] t2_r9_c0_rr0;
  wire [15:0] t2_r9_c0_rr1;
  wire [15:0] t2_r9_c0_rr2;
  wire [15:0] t2_r9_c0_rr3;
  wire [15:0] t3_r9_c0_rr0;
  wire [15:0] t3_r9_c0_rr1;
  wire [15:0] t4_r9_c0_rr0;
  wire [15:0] t0_r9_c1_rr0;
  wire [15:0] t0_r9_c1_rr1;
  wire [15:0] t0_r9_c1_rr2;
  wire [15:0] t0_r9_c1_rr3;
  wire [15:0] t0_r9_c1_rr4;
  wire [15:0] t0_r9_c1_rr5;
  wire [15:0] t0_r9_c1_rr6;
  wire [15:0] t0_r9_c1_rr7;
  wire [15:0] t0_r9_c1_rr8;
  wire [15:0] t0_r9_c1_rr9;
  wire [15:0] t0_r9_c1_rr10;
  wire [15:0] t0_r9_c1_rr11;
  wire [15:0] t0_r9_c1_rr12;
  wire [15:0] t0_r9_c1_rr13;
  wire [15:0] t0_r9_c1_rr14;
  wire [15:0] t1_r9_c1_rr0;
  wire [15:0] t1_r9_c1_rr1;
  wire [15:0] t1_r9_c1_rr2;
  wire [15:0] t1_r9_c1_rr3;
  wire [15:0] t1_r9_c1_rr4;
  wire [15:0] t1_r9_c1_rr5;
  wire [15:0] t1_r9_c1_rr6;
  wire [15:0] t1_r9_c1_rr7;
  wire [15:0] t2_r9_c1_rr0;
  wire [15:0] t2_r9_c1_rr1;
  wire [15:0] t2_r9_c1_rr2;
  wire [15:0] t2_r9_c1_rr3;
  wire [15:0] t3_r9_c1_rr0;
  wire [15:0] t3_r9_c1_rr1;
  wire [15:0] t4_r9_c1_rr0;
  wire [15:0] t0_r9_c2_rr0;
  wire [15:0] t0_r9_c2_rr1;
  wire [15:0] t0_r9_c2_rr2;
  wire [15:0] t0_r9_c2_rr3;
  wire [15:0] t0_r9_c2_rr4;
  wire [15:0] t0_r9_c2_rr5;
  wire [15:0] t0_r9_c2_rr6;
  wire [15:0] t0_r9_c2_rr7;
  wire [15:0] t0_r9_c2_rr8;
  wire [15:0] t0_r9_c2_rr9;
  wire [15:0] t0_r9_c2_rr10;
  wire [15:0] t0_r9_c2_rr11;
  wire [15:0] t0_r9_c2_rr12;
  wire [15:0] t0_r9_c2_rr13;
  wire [15:0] t0_r9_c2_rr14;
  wire [15:0] t1_r9_c2_rr0;
  wire [15:0] t1_r9_c2_rr1;
  wire [15:0] t1_r9_c2_rr2;
  wire [15:0] t1_r9_c2_rr3;
  wire [15:0] t1_r9_c2_rr4;
  wire [15:0] t1_r9_c2_rr5;
  wire [15:0] t1_r9_c2_rr6;
  wire [15:0] t1_r9_c2_rr7;
  wire [15:0] t2_r9_c2_rr0;
  wire [15:0] t2_r9_c2_rr1;
  wire [15:0] t2_r9_c2_rr2;
  wire [15:0] t2_r9_c2_rr3;
  wire [15:0] t3_r9_c2_rr0;
  wire [15:0] t3_r9_c2_rr1;
  wire [15:0] t4_r9_c2_rr0;
  wire [15:0] t0_r9_c3_rr0;
  wire [15:0] t0_r9_c3_rr1;
  wire [15:0] t0_r9_c3_rr2;
  wire [15:0] t0_r9_c3_rr3;
  wire [15:0] t0_r9_c3_rr4;
  wire [15:0] t0_r9_c3_rr5;
  wire [15:0] t0_r9_c3_rr6;
  wire [15:0] t0_r9_c3_rr7;
  wire [15:0] t0_r9_c3_rr8;
  wire [15:0] t0_r9_c3_rr9;
  wire [15:0] t0_r9_c3_rr10;
  wire [15:0] t0_r9_c3_rr11;
  wire [15:0] t0_r9_c3_rr12;
  wire [15:0] t0_r9_c3_rr13;
  wire [15:0] t0_r9_c3_rr14;
  wire [15:0] t1_r9_c3_rr0;
  wire [15:0] t1_r9_c3_rr1;
  wire [15:0] t1_r9_c3_rr2;
  wire [15:0] t1_r9_c3_rr3;
  wire [15:0] t1_r9_c3_rr4;
  wire [15:0] t1_r9_c3_rr5;
  wire [15:0] t1_r9_c3_rr6;
  wire [15:0] t1_r9_c3_rr7;
  wire [15:0] t2_r9_c3_rr0;
  wire [15:0] t2_r9_c3_rr1;
  wire [15:0] t2_r9_c3_rr2;
  wire [15:0] t2_r9_c3_rr3;
  wire [15:0] t3_r9_c3_rr0;
  wire [15:0] t3_r9_c3_rr1;
  wire [15:0] t4_r9_c3_rr0;
  wire [15:0] t0_r9_c4_rr0;
  wire [15:0] t0_r9_c4_rr1;
  wire [15:0] t0_r9_c4_rr2;
  wire [15:0] t0_r9_c4_rr3;
  wire [15:0] t0_r9_c4_rr4;
  wire [15:0] t0_r9_c4_rr5;
  wire [15:0] t0_r9_c4_rr6;
  wire [15:0] t0_r9_c4_rr7;
  wire [15:0] t0_r9_c4_rr8;
  wire [15:0] t0_r9_c4_rr9;
  wire [15:0] t0_r9_c4_rr10;
  wire [15:0] t0_r9_c4_rr11;
  wire [15:0] t0_r9_c4_rr12;
  wire [15:0] t0_r9_c4_rr13;
  wire [15:0] t0_r9_c4_rr14;
  wire [15:0] t1_r9_c4_rr0;
  wire [15:0] t1_r9_c4_rr1;
  wire [15:0] t1_r9_c4_rr2;
  wire [15:0] t1_r9_c4_rr3;
  wire [15:0] t1_r9_c4_rr4;
  wire [15:0] t1_r9_c4_rr5;
  wire [15:0] t1_r9_c4_rr6;
  wire [15:0] t1_r9_c4_rr7;
  wire [15:0] t2_r9_c4_rr0;
  wire [15:0] t2_r9_c4_rr1;
  wire [15:0] t2_r9_c4_rr2;
  wire [15:0] t2_r9_c4_rr3;
  wire [15:0] t3_r9_c4_rr0;
  wire [15:0] t3_r9_c4_rr1;
  wire [15:0] t4_r9_c4_rr0;
  wire [15:0] t0_r9_c5_rr0;
  wire [15:0] t0_r9_c5_rr1;
  wire [15:0] t0_r9_c5_rr2;
  wire [15:0] t0_r9_c5_rr3;
  wire [15:0] t0_r9_c5_rr4;
  wire [15:0] t0_r9_c5_rr5;
  wire [15:0] t0_r9_c5_rr6;
  wire [15:0] t0_r9_c5_rr7;
  wire [15:0] t0_r9_c5_rr8;
  wire [15:0] t0_r9_c5_rr9;
  wire [15:0] t0_r9_c5_rr10;
  wire [15:0] t0_r9_c5_rr11;
  wire [15:0] t0_r9_c5_rr12;
  wire [15:0] t0_r9_c5_rr13;
  wire [15:0] t0_r9_c5_rr14;
  wire [15:0] t1_r9_c5_rr0;
  wire [15:0] t1_r9_c5_rr1;
  wire [15:0] t1_r9_c5_rr2;
  wire [15:0] t1_r9_c5_rr3;
  wire [15:0] t1_r9_c5_rr4;
  wire [15:0] t1_r9_c5_rr5;
  wire [15:0] t1_r9_c5_rr6;
  wire [15:0] t1_r9_c5_rr7;
  wire [15:0] t2_r9_c5_rr0;
  wire [15:0] t2_r9_c5_rr1;
  wire [15:0] t2_r9_c5_rr2;
  wire [15:0] t2_r9_c5_rr3;
  wire [15:0] t3_r9_c5_rr0;
  wire [15:0] t3_r9_c5_rr1;
  wire [15:0] t4_r9_c5_rr0;
  wire [15:0] t0_r9_c6_rr0;
  wire [15:0] t0_r9_c6_rr1;
  wire [15:0] t0_r9_c6_rr2;
  wire [15:0] t0_r9_c6_rr3;
  wire [15:0] t0_r9_c6_rr4;
  wire [15:0] t0_r9_c6_rr5;
  wire [15:0] t0_r9_c6_rr6;
  wire [15:0] t0_r9_c6_rr7;
  wire [15:0] t0_r9_c6_rr8;
  wire [15:0] t0_r9_c6_rr9;
  wire [15:0] t0_r9_c6_rr10;
  wire [15:0] t0_r9_c6_rr11;
  wire [15:0] t0_r9_c6_rr12;
  wire [15:0] t0_r9_c6_rr13;
  wire [15:0] t0_r9_c6_rr14;
  wire [15:0] t1_r9_c6_rr0;
  wire [15:0] t1_r9_c6_rr1;
  wire [15:0] t1_r9_c6_rr2;
  wire [15:0] t1_r9_c6_rr3;
  wire [15:0] t1_r9_c6_rr4;
  wire [15:0] t1_r9_c6_rr5;
  wire [15:0] t1_r9_c6_rr6;
  wire [15:0] t1_r9_c6_rr7;
  wire [15:0] t2_r9_c6_rr0;
  wire [15:0] t2_r9_c6_rr1;
  wire [15:0] t2_r9_c6_rr2;
  wire [15:0] t2_r9_c6_rr3;
  wire [15:0] t3_r9_c6_rr0;
  wire [15:0] t3_r9_c6_rr1;
  wire [15:0] t4_r9_c6_rr0;
  wire [15:0] t0_r9_c7_rr0;
  wire [15:0] t0_r9_c7_rr1;
  wire [15:0] t0_r9_c7_rr2;
  wire [15:0] t0_r9_c7_rr3;
  wire [15:0] t0_r9_c7_rr4;
  wire [15:0] t0_r9_c7_rr5;
  wire [15:0] t0_r9_c7_rr6;
  wire [15:0] t0_r9_c7_rr7;
  wire [15:0] t0_r9_c7_rr8;
  wire [15:0] t0_r9_c7_rr9;
  wire [15:0] t0_r9_c7_rr10;
  wire [15:0] t0_r9_c7_rr11;
  wire [15:0] t0_r9_c7_rr12;
  wire [15:0] t0_r9_c7_rr13;
  wire [15:0] t0_r9_c7_rr14;
  wire [15:0] t1_r9_c7_rr0;
  wire [15:0] t1_r9_c7_rr1;
  wire [15:0] t1_r9_c7_rr2;
  wire [15:0] t1_r9_c7_rr3;
  wire [15:0] t1_r9_c7_rr4;
  wire [15:0] t1_r9_c7_rr5;
  wire [15:0] t1_r9_c7_rr6;
  wire [15:0] t1_r9_c7_rr7;
  wire [15:0] t2_r9_c7_rr0;
  wire [15:0] t2_r9_c7_rr1;
  wire [15:0] t2_r9_c7_rr2;
  wire [15:0] t2_r9_c7_rr3;
  wire [15:0] t3_r9_c7_rr0;
  wire [15:0] t3_r9_c7_rr1;
  wire [15:0] t4_r9_c7_rr0;
  wire [15:0] t0_r9_c8_rr0;
  wire [15:0] t0_r9_c8_rr1;
  wire [15:0] t0_r9_c8_rr2;
  wire [15:0] t0_r9_c8_rr3;
  wire [15:0] t0_r9_c8_rr4;
  wire [15:0] t0_r9_c8_rr5;
  wire [15:0] t0_r9_c8_rr6;
  wire [15:0] t0_r9_c8_rr7;
  wire [15:0] t0_r9_c8_rr8;
  wire [15:0] t0_r9_c8_rr9;
  wire [15:0] t0_r9_c8_rr10;
  wire [15:0] t0_r9_c8_rr11;
  wire [15:0] t0_r9_c8_rr12;
  wire [15:0] t0_r9_c8_rr13;
  wire [15:0] t0_r9_c8_rr14;
  wire [15:0] t1_r9_c8_rr0;
  wire [15:0] t1_r9_c8_rr1;
  wire [15:0] t1_r9_c8_rr2;
  wire [15:0] t1_r9_c8_rr3;
  wire [15:0] t1_r9_c8_rr4;
  wire [15:0] t1_r9_c8_rr5;
  wire [15:0] t1_r9_c8_rr6;
  wire [15:0] t1_r9_c8_rr7;
  wire [15:0] t2_r9_c8_rr0;
  wire [15:0] t2_r9_c8_rr1;
  wire [15:0] t2_r9_c8_rr2;
  wire [15:0] t2_r9_c8_rr3;
  wire [15:0] t3_r9_c8_rr0;
  wire [15:0] t3_r9_c8_rr1;
  wire [15:0] t4_r9_c8_rr0;
  wire [15:0] t0_r9_c9_rr0;
  wire [15:0] t0_r9_c9_rr1;
  wire [15:0] t0_r9_c9_rr2;
  wire [15:0] t0_r9_c9_rr3;
  wire [15:0] t0_r9_c9_rr4;
  wire [15:0] t0_r9_c9_rr5;
  wire [15:0] t0_r9_c9_rr6;
  wire [15:0] t0_r9_c9_rr7;
  wire [15:0] t0_r9_c9_rr8;
  wire [15:0] t0_r9_c9_rr9;
  wire [15:0] t0_r9_c9_rr10;
  wire [15:0] t0_r9_c9_rr11;
  wire [15:0] t0_r9_c9_rr12;
  wire [15:0] t0_r9_c9_rr13;
  wire [15:0] t0_r9_c9_rr14;
  wire [15:0] t1_r9_c9_rr0;
  wire [15:0] t1_r9_c9_rr1;
  wire [15:0] t1_r9_c9_rr2;
  wire [15:0] t1_r9_c9_rr3;
  wire [15:0] t1_r9_c9_rr4;
  wire [15:0] t1_r9_c9_rr5;
  wire [15:0] t1_r9_c9_rr6;
  wire [15:0] t1_r9_c9_rr7;
  wire [15:0] t2_r9_c9_rr0;
  wire [15:0] t2_r9_c9_rr1;
  wire [15:0] t2_r9_c9_rr2;
  wire [15:0] t2_r9_c9_rr3;
  wire [15:0] t3_r9_c9_rr0;
  wire [15:0] t3_r9_c9_rr1;
  wire [15:0] t4_r9_c9_rr0;
  wire [15:0] t0_r9_c10_rr0;
  wire [15:0] t0_r9_c10_rr1;
  wire [15:0] t0_r9_c10_rr2;
  wire [15:0] t0_r9_c10_rr3;
  wire [15:0] t0_r9_c10_rr4;
  wire [15:0] t0_r9_c10_rr5;
  wire [15:0] t0_r9_c10_rr6;
  wire [15:0] t0_r9_c10_rr7;
  wire [15:0] t0_r9_c10_rr8;
  wire [15:0] t0_r9_c10_rr9;
  wire [15:0] t0_r9_c10_rr10;
  wire [15:0] t0_r9_c10_rr11;
  wire [15:0] t0_r9_c10_rr12;
  wire [15:0] t0_r9_c10_rr13;
  wire [15:0] t0_r9_c10_rr14;
  wire [15:0] t1_r9_c10_rr0;
  wire [15:0] t1_r9_c10_rr1;
  wire [15:0] t1_r9_c10_rr2;
  wire [15:0] t1_r9_c10_rr3;
  wire [15:0] t1_r9_c10_rr4;
  wire [15:0] t1_r9_c10_rr5;
  wire [15:0] t1_r9_c10_rr6;
  wire [15:0] t1_r9_c10_rr7;
  wire [15:0] t2_r9_c10_rr0;
  wire [15:0] t2_r9_c10_rr1;
  wire [15:0] t2_r9_c10_rr2;
  wire [15:0] t2_r9_c10_rr3;
  wire [15:0] t3_r9_c10_rr0;
  wire [15:0] t3_r9_c10_rr1;
  wire [15:0] t4_r9_c10_rr0;
  wire [15:0] t0_r9_c11_rr0;
  wire [15:0] t0_r9_c11_rr1;
  wire [15:0] t0_r9_c11_rr2;
  wire [15:0] t0_r9_c11_rr3;
  wire [15:0] t0_r9_c11_rr4;
  wire [15:0] t0_r9_c11_rr5;
  wire [15:0] t0_r9_c11_rr6;
  wire [15:0] t0_r9_c11_rr7;
  wire [15:0] t0_r9_c11_rr8;
  wire [15:0] t0_r9_c11_rr9;
  wire [15:0] t0_r9_c11_rr10;
  wire [15:0] t0_r9_c11_rr11;
  wire [15:0] t0_r9_c11_rr12;
  wire [15:0] t0_r9_c11_rr13;
  wire [15:0] t0_r9_c11_rr14;
  wire [15:0] t1_r9_c11_rr0;
  wire [15:0] t1_r9_c11_rr1;
  wire [15:0] t1_r9_c11_rr2;
  wire [15:0] t1_r9_c11_rr3;
  wire [15:0] t1_r9_c11_rr4;
  wire [15:0] t1_r9_c11_rr5;
  wire [15:0] t1_r9_c11_rr6;
  wire [15:0] t1_r9_c11_rr7;
  wire [15:0] t2_r9_c11_rr0;
  wire [15:0] t2_r9_c11_rr1;
  wire [15:0] t2_r9_c11_rr2;
  wire [15:0] t2_r9_c11_rr3;
  wire [15:0] t3_r9_c11_rr0;
  wire [15:0] t3_r9_c11_rr1;
  wire [15:0] t4_r9_c11_rr0;
  wire [15:0] t0_r9_c12_rr0;
  wire [15:0] t0_r9_c12_rr1;
  wire [15:0] t0_r9_c12_rr2;
  wire [15:0] t0_r9_c12_rr3;
  wire [15:0] t0_r9_c12_rr4;
  wire [15:0] t0_r9_c12_rr5;
  wire [15:0] t0_r9_c12_rr6;
  wire [15:0] t0_r9_c12_rr7;
  wire [15:0] t0_r9_c12_rr8;
  wire [15:0] t0_r9_c12_rr9;
  wire [15:0] t0_r9_c12_rr10;
  wire [15:0] t0_r9_c12_rr11;
  wire [15:0] t0_r9_c12_rr12;
  wire [15:0] t0_r9_c12_rr13;
  wire [15:0] t0_r9_c12_rr14;
  wire [15:0] t1_r9_c12_rr0;
  wire [15:0] t1_r9_c12_rr1;
  wire [15:0] t1_r9_c12_rr2;
  wire [15:0] t1_r9_c12_rr3;
  wire [15:0] t1_r9_c12_rr4;
  wire [15:0] t1_r9_c12_rr5;
  wire [15:0] t1_r9_c12_rr6;
  wire [15:0] t1_r9_c12_rr7;
  wire [15:0] t2_r9_c12_rr0;
  wire [15:0] t2_r9_c12_rr1;
  wire [15:0] t2_r9_c12_rr2;
  wire [15:0] t2_r9_c12_rr3;
  wire [15:0] t3_r9_c12_rr0;
  wire [15:0] t3_r9_c12_rr1;
  wire [15:0] t4_r9_c12_rr0;
  wire [15:0] t0_r9_c13_rr0;
  wire [15:0] t0_r9_c13_rr1;
  wire [15:0] t0_r9_c13_rr2;
  wire [15:0] t0_r9_c13_rr3;
  wire [15:0] t0_r9_c13_rr4;
  wire [15:0] t0_r9_c13_rr5;
  wire [15:0] t0_r9_c13_rr6;
  wire [15:0] t0_r9_c13_rr7;
  wire [15:0] t0_r9_c13_rr8;
  wire [15:0] t0_r9_c13_rr9;
  wire [15:0] t0_r9_c13_rr10;
  wire [15:0] t0_r9_c13_rr11;
  wire [15:0] t0_r9_c13_rr12;
  wire [15:0] t0_r9_c13_rr13;
  wire [15:0] t0_r9_c13_rr14;
  wire [15:0] t1_r9_c13_rr0;
  wire [15:0] t1_r9_c13_rr1;
  wire [15:0] t1_r9_c13_rr2;
  wire [15:0] t1_r9_c13_rr3;
  wire [15:0] t1_r9_c13_rr4;
  wire [15:0] t1_r9_c13_rr5;
  wire [15:0] t1_r9_c13_rr6;
  wire [15:0] t1_r9_c13_rr7;
  wire [15:0] t2_r9_c13_rr0;
  wire [15:0] t2_r9_c13_rr1;
  wire [15:0] t2_r9_c13_rr2;
  wire [15:0] t2_r9_c13_rr3;
  wire [15:0] t3_r9_c13_rr0;
  wire [15:0] t3_r9_c13_rr1;
  wire [15:0] t4_r9_c13_rr0;
  wire [15:0] t0_r9_c14_rr0;
  wire [15:0] t0_r9_c14_rr1;
  wire [15:0] t0_r9_c14_rr2;
  wire [15:0] t0_r9_c14_rr3;
  wire [15:0] t0_r9_c14_rr4;
  wire [15:0] t0_r9_c14_rr5;
  wire [15:0] t0_r9_c14_rr6;
  wire [15:0] t0_r9_c14_rr7;
  wire [15:0] t0_r9_c14_rr8;
  wire [15:0] t0_r9_c14_rr9;
  wire [15:0] t0_r9_c14_rr10;
  wire [15:0] t0_r9_c14_rr11;
  wire [15:0] t0_r9_c14_rr12;
  wire [15:0] t0_r9_c14_rr13;
  wire [15:0] t0_r9_c14_rr14;
  wire [15:0] t1_r9_c14_rr0;
  wire [15:0] t1_r9_c14_rr1;
  wire [15:0] t1_r9_c14_rr2;
  wire [15:0] t1_r9_c14_rr3;
  wire [15:0] t1_r9_c14_rr4;
  wire [15:0] t1_r9_c14_rr5;
  wire [15:0] t1_r9_c14_rr6;
  wire [15:0] t1_r9_c14_rr7;
  wire [15:0] t2_r9_c14_rr0;
  wire [15:0] t2_r9_c14_rr1;
  wire [15:0] t2_r9_c14_rr2;
  wire [15:0] t2_r9_c14_rr3;
  wire [15:0] t3_r9_c14_rr0;
  wire [15:0] t3_r9_c14_rr1;
  wire [15:0] t4_r9_c14_rr0;
  wire [15:0] t0_r10_c0_rr0;
  wire [15:0] t0_r10_c0_rr1;
  wire [15:0] t0_r10_c0_rr2;
  wire [15:0] t0_r10_c0_rr3;
  wire [15:0] t0_r10_c0_rr4;
  wire [15:0] t0_r10_c0_rr5;
  wire [15:0] t0_r10_c0_rr6;
  wire [15:0] t0_r10_c0_rr7;
  wire [15:0] t0_r10_c0_rr8;
  wire [15:0] t0_r10_c0_rr9;
  wire [15:0] t0_r10_c0_rr10;
  wire [15:0] t0_r10_c0_rr11;
  wire [15:0] t0_r10_c0_rr12;
  wire [15:0] t0_r10_c0_rr13;
  wire [15:0] t0_r10_c0_rr14;
  wire [15:0] t1_r10_c0_rr0;
  wire [15:0] t1_r10_c0_rr1;
  wire [15:0] t1_r10_c0_rr2;
  wire [15:0] t1_r10_c0_rr3;
  wire [15:0] t1_r10_c0_rr4;
  wire [15:0] t1_r10_c0_rr5;
  wire [15:0] t1_r10_c0_rr6;
  wire [15:0] t1_r10_c0_rr7;
  wire [15:0] t2_r10_c0_rr0;
  wire [15:0] t2_r10_c0_rr1;
  wire [15:0] t2_r10_c0_rr2;
  wire [15:0] t2_r10_c0_rr3;
  wire [15:0] t3_r10_c0_rr0;
  wire [15:0] t3_r10_c0_rr1;
  wire [15:0] t4_r10_c0_rr0;
  wire [15:0] t0_r10_c1_rr0;
  wire [15:0] t0_r10_c1_rr1;
  wire [15:0] t0_r10_c1_rr2;
  wire [15:0] t0_r10_c1_rr3;
  wire [15:0] t0_r10_c1_rr4;
  wire [15:0] t0_r10_c1_rr5;
  wire [15:0] t0_r10_c1_rr6;
  wire [15:0] t0_r10_c1_rr7;
  wire [15:0] t0_r10_c1_rr8;
  wire [15:0] t0_r10_c1_rr9;
  wire [15:0] t0_r10_c1_rr10;
  wire [15:0] t0_r10_c1_rr11;
  wire [15:0] t0_r10_c1_rr12;
  wire [15:0] t0_r10_c1_rr13;
  wire [15:0] t0_r10_c1_rr14;
  wire [15:0] t1_r10_c1_rr0;
  wire [15:0] t1_r10_c1_rr1;
  wire [15:0] t1_r10_c1_rr2;
  wire [15:0] t1_r10_c1_rr3;
  wire [15:0] t1_r10_c1_rr4;
  wire [15:0] t1_r10_c1_rr5;
  wire [15:0] t1_r10_c1_rr6;
  wire [15:0] t1_r10_c1_rr7;
  wire [15:0] t2_r10_c1_rr0;
  wire [15:0] t2_r10_c1_rr1;
  wire [15:0] t2_r10_c1_rr2;
  wire [15:0] t2_r10_c1_rr3;
  wire [15:0] t3_r10_c1_rr0;
  wire [15:0] t3_r10_c1_rr1;
  wire [15:0] t4_r10_c1_rr0;
  wire [15:0] t0_r10_c2_rr0;
  wire [15:0] t0_r10_c2_rr1;
  wire [15:0] t0_r10_c2_rr2;
  wire [15:0] t0_r10_c2_rr3;
  wire [15:0] t0_r10_c2_rr4;
  wire [15:0] t0_r10_c2_rr5;
  wire [15:0] t0_r10_c2_rr6;
  wire [15:0] t0_r10_c2_rr7;
  wire [15:0] t0_r10_c2_rr8;
  wire [15:0] t0_r10_c2_rr9;
  wire [15:0] t0_r10_c2_rr10;
  wire [15:0] t0_r10_c2_rr11;
  wire [15:0] t0_r10_c2_rr12;
  wire [15:0] t0_r10_c2_rr13;
  wire [15:0] t0_r10_c2_rr14;
  wire [15:0] t1_r10_c2_rr0;
  wire [15:0] t1_r10_c2_rr1;
  wire [15:0] t1_r10_c2_rr2;
  wire [15:0] t1_r10_c2_rr3;
  wire [15:0] t1_r10_c2_rr4;
  wire [15:0] t1_r10_c2_rr5;
  wire [15:0] t1_r10_c2_rr6;
  wire [15:0] t1_r10_c2_rr7;
  wire [15:0] t2_r10_c2_rr0;
  wire [15:0] t2_r10_c2_rr1;
  wire [15:0] t2_r10_c2_rr2;
  wire [15:0] t2_r10_c2_rr3;
  wire [15:0] t3_r10_c2_rr0;
  wire [15:0] t3_r10_c2_rr1;
  wire [15:0] t4_r10_c2_rr0;
  wire [15:0] t0_r10_c3_rr0;
  wire [15:0] t0_r10_c3_rr1;
  wire [15:0] t0_r10_c3_rr2;
  wire [15:0] t0_r10_c3_rr3;
  wire [15:0] t0_r10_c3_rr4;
  wire [15:0] t0_r10_c3_rr5;
  wire [15:0] t0_r10_c3_rr6;
  wire [15:0] t0_r10_c3_rr7;
  wire [15:0] t0_r10_c3_rr8;
  wire [15:0] t0_r10_c3_rr9;
  wire [15:0] t0_r10_c3_rr10;
  wire [15:0] t0_r10_c3_rr11;
  wire [15:0] t0_r10_c3_rr12;
  wire [15:0] t0_r10_c3_rr13;
  wire [15:0] t0_r10_c3_rr14;
  wire [15:0] t1_r10_c3_rr0;
  wire [15:0] t1_r10_c3_rr1;
  wire [15:0] t1_r10_c3_rr2;
  wire [15:0] t1_r10_c3_rr3;
  wire [15:0] t1_r10_c3_rr4;
  wire [15:0] t1_r10_c3_rr5;
  wire [15:0] t1_r10_c3_rr6;
  wire [15:0] t1_r10_c3_rr7;
  wire [15:0] t2_r10_c3_rr0;
  wire [15:0] t2_r10_c3_rr1;
  wire [15:0] t2_r10_c3_rr2;
  wire [15:0] t2_r10_c3_rr3;
  wire [15:0] t3_r10_c3_rr0;
  wire [15:0] t3_r10_c3_rr1;
  wire [15:0] t4_r10_c3_rr0;
  wire [15:0] t0_r10_c4_rr0;
  wire [15:0] t0_r10_c4_rr1;
  wire [15:0] t0_r10_c4_rr2;
  wire [15:0] t0_r10_c4_rr3;
  wire [15:0] t0_r10_c4_rr4;
  wire [15:0] t0_r10_c4_rr5;
  wire [15:0] t0_r10_c4_rr6;
  wire [15:0] t0_r10_c4_rr7;
  wire [15:0] t0_r10_c4_rr8;
  wire [15:0] t0_r10_c4_rr9;
  wire [15:0] t0_r10_c4_rr10;
  wire [15:0] t0_r10_c4_rr11;
  wire [15:0] t0_r10_c4_rr12;
  wire [15:0] t0_r10_c4_rr13;
  wire [15:0] t0_r10_c4_rr14;
  wire [15:0] t1_r10_c4_rr0;
  wire [15:0] t1_r10_c4_rr1;
  wire [15:0] t1_r10_c4_rr2;
  wire [15:0] t1_r10_c4_rr3;
  wire [15:0] t1_r10_c4_rr4;
  wire [15:0] t1_r10_c4_rr5;
  wire [15:0] t1_r10_c4_rr6;
  wire [15:0] t1_r10_c4_rr7;
  wire [15:0] t2_r10_c4_rr0;
  wire [15:0] t2_r10_c4_rr1;
  wire [15:0] t2_r10_c4_rr2;
  wire [15:0] t2_r10_c4_rr3;
  wire [15:0] t3_r10_c4_rr0;
  wire [15:0] t3_r10_c4_rr1;
  wire [15:0] t4_r10_c4_rr0;
  wire [15:0] t0_r10_c5_rr0;
  wire [15:0] t0_r10_c5_rr1;
  wire [15:0] t0_r10_c5_rr2;
  wire [15:0] t0_r10_c5_rr3;
  wire [15:0] t0_r10_c5_rr4;
  wire [15:0] t0_r10_c5_rr5;
  wire [15:0] t0_r10_c5_rr6;
  wire [15:0] t0_r10_c5_rr7;
  wire [15:0] t0_r10_c5_rr8;
  wire [15:0] t0_r10_c5_rr9;
  wire [15:0] t0_r10_c5_rr10;
  wire [15:0] t0_r10_c5_rr11;
  wire [15:0] t0_r10_c5_rr12;
  wire [15:0] t0_r10_c5_rr13;
  wire [15:0] t0_r10_c5_rr14;
  wire [15:0] t1_r10_c5_rr0;
  wire [15:0] t1_r10_c5_rr1;
  wire [15:0] t1_r10_c5_rr2;
  wire [15:0] t1_r10_c5_rr3;
  wire [15:0] t1_r10_c5_rr4;
  wire [15:0] t1_r10_c5_rr5;
  wire [15:0] t1_r10_c5_rr6;
  wire [15:0] t1_r10_c5_rr7;
  wire [15:0] t2_r10_c5_rr0;
  wire [15:0] t2_r10_c5_rr1;
  wire [15:0] t2_r10_c5_rr2;
  wire [15:0] t2_r10_c5_rr3;
  wire [15:0] t3_r10_c5_rr0;
  wire [15:0] t3_r10_c5_rr1;
  wire [15:0] t4_r10_c5_rr0;
  wire [15:0] t0_r10_c6_rr0;
  wire [15:0] t0_r10_c6_rr1;
  wire [15:0] t0_r10_c6_rr2;
  wire [15:0] t0_r10_c6_rr3;
  wire [15:0] t0_r10_c6_rr4;
  wire [15:0] t0_r10_c6_rr5;
  wire [15:0] t0_r10_c6_rr6;
  wire [15:0] t0_r10_c6_rr7;
  wire [15:0] t0_r10_c6_rr8;
  wire [15:0] t0_r10_c6_rr9;
  wire [15:0] t0_r10_c6_rr10;
  wire [15:0] t0_r10_c6_rr11;
  wire [15:0] t0_r10_c6_rr12;
  wire [15:0] t0_r10_c6_rr13;
  wire [15:0] t0_r10_c6_rr14;
  wire [15:0] t1_r10_c6_rr0;
  wire [15:0] t1_r10_c6_rr1;
  wire [15:0] t1_r10_c6_rr2;
  wire [15:0] t1_r10_c6_rr3;
  wire [15:0] t1_r10_c6_rr4;
  wire [15:0] t1_r10_c6_rr5;
  wire [15:0] t1_r10_c6_rr6;
  wire [15:0] t1_r10_c6_rr7;
  wire [15:0] t2_r10_c6_rr0;
  wire [15:0] t2_r10_c6_rr1;
  wire [15:0] t2_r10_c6_rr2;
  wire [15:0] t2_r10_c6_rr3;
  wire [15:0] t3_r10_c6_rr0;
  wire [15:0] t3_r10_c6_rr1;
  wire [15:0] t4_r10_c6_rr0;
  wire [15:0] t0_r10_c7_rr0;
  wire [15:0] t0_r10_c7_rr1;
  wire [15:0] t0_r10_c7_rr2;
  wire [15:0] t0_r10_c7_rr3;
  wire [15:0] t0_r10_c7_rr4;
  wire [15:0] t0_r10_c7_rr5;
  wire [15:0] t0_r10_c7_rr6;
  wire [15:0] t0_r10_c7_rr7;
  wire [15:0] t0_r10_c7_rr8;
  wire [15:0] t0_r10_c7_rr9;
  wire [15:0] t0_r10_c7_rr10;
  wire [15:0] t0_r10_c7_rr11;
  wire [15:0] t0_r10_c7_rr12;
  wire [15:0] t0_r10_c7_rr13;
  wire [15:0] t0_r10_c7_rr14;
  wire [15:0] t1_r10_c7_rr0;
  wire [15:0] t1_r10_c7_rr1;
  wire [15:0] t1_r10_c7_rr2;
  wire [15:0] t1_r10_c7_rr3;
  wire [15:0] t1_r10_c7_rr4;
  wire [15:0] t1_r10_c7_rr5;
  wire [15:0] t1_r10_c7_rr6;
  wire [15:0] t1_r10_c7_rr7;
  wire [15:0] t2_r10_c7_rr0;
  wire [15:0] t2_r10_c7_rr1;
  wire [15:0] t2_r10_c7_rr2;
  wire [15:0] t2_r10_c7_rr3;
  wire [15:0] t3_r10_c7_rr0;
  wire [15:0] t3_r10_c7_rr1;
  wire [15:0] t4_r10_c7_rr0;
  wire [15:0] t0_r10_c8_rr0;
  wire [15:0] t0_r10_c8_rr1;
  wire [15:0] t0_r10_c8_rr2;
  wire [15:0] t0_r10_c8_rr3;
  wire [15:0] t0_r10_c8_rr4;
  wire [15:0] t0_r10_c8_rr5;
  wire [15:0] t0_r10_c8_rr6;
  wire [15:0] t0_r10_c8_rr7;
  wire [15:0] t0_r10_c8_rr8;
  wire [15:0] t0_r10_c8_rr9;
  wire [15:0] t0_r10_c8_rr10;
  wire [15:0] t0_r10_c8_rr11;
  wire [15:0] t0_r10_c8_rr12;
  wire [15:0] t0_r10_c8_rr13;
  wire [15:0] t0_r10_c8_rr14;
  wire [15:0] t1_r10_c8_rr0;
  wire [15:0] t1_r10_c8_rr1;
  wire [15:0] t1_r10_c8_rr2;
  wire [15:0] t1_r10_c8_rr3;
  wire [15:0] t1_r10_c8_rr4;
  wire [15:0] t1_r10_c8_rr5;
  wire [15:0] t1_r10_c8_rr6;
  wire [15:0] t1_r10_c8_rr7;
  wire [15:0] t2_r10_c8_rr0;
  wire [15:0] t2_r10_c8_rr1;
  wire [15:0] t2_r10_c8_rr2;
  wire [15:0] t2_r10_c8_rr3;
  wire [15:0] t3_r10_c8_rr0;
  wire [15:0] t3_r10_c8_rr1;
  wire [15:0] t4_r10_c8_rr0;
  wire [15:0] t0_r10_c9_rr0;
  wire [15:0] t0_r10_c9_rr1;
  wire [15:0] t0_r10_c9_rr2;
  wire [15:0] t0_r10_c9_rr3;
  wire [15:0] t0_r10_c9_rr4;
  wire [15:0] t0_r10_c9_rr5;
  wire [15:0] t0_r10_c9_rr6;
  wire [15:0] t0_r10_c9_rr7;
  wire [15:0] t0_r10_c9_rr8;
  wire [15:0] t0_r10_c9_rr9;
  wire [15:0] t0_r10_c9_rr10;
  wire [15:0] t0_r10_c9_rr11;
  wire [15:0] t0_r10_c9_rr12;
  wire [15:0] t0_r10_c9_rr13;
  wire [15:0] t0_r10_c9_rr14;
  wire [15:0] t1_r10_c9_rr0;
  wire [15:0] t1_r10_c9_rr1;
  wire [15:0] t1_r10_c9_rr2;
  wire [15:0] t1_r10_c9_rr3;
  wire [15:0] t1_r10_c9_rr4;
  wire [15:0] t1_r10_c9_rr5;
  wire [15:0] t1_r10_c9_rr6;
  wire [15:0] t1_r10_c9_rr7;
  wire [15:0] t2_r10_c9_rr0;
  wire [15:0] t2_r10_c9_rr1;
  wire [15:0] t2_r10_c9_rr2;
  wire [15:0] t2_r10_c9_rr3;
  wire [15:0] t3_r10_c9_rr0;
  wire [15:0] t3_r10_c9_rr1;
  wire [15:0] t4_r10_c9_rr0;
  wire [15:0] t0_r10_c10_rr0;
  wire [15:0] t0_r10_c10_rr1;
  wire [15:0] t0_r10_c10_rr2;
  wire [15:0] t0_r10_c10_rr3;
  wire [15:0] t0_r10_c10_rr4;
  wire [15:0] t0_r10_c10_rr5;
  wire [15:0] t0_r10_c10_rr6;
  wire [15:0] t0_r10_c10_rr7;
  wire [15:0] t0_r10_c10_rr8;
  wire [15:0] t0_r10_c10_rr9;
  wire [15:0] t0_r10_c10_rr10;
  wire [15:0] t0_r10_c10_rr11;
  wire [15:0] t0_r10_c10_rr12;
  wire [15:0] t0_r10_c10_rr13;
  wire [15:0] t0_r10_c10_rr14;
  wire [15:0] t1_r10_c10_rr0;
  wire [15:0] t1_r10_c10_rr1;
  wire [15:0] t1_r10_c10_rr2;
  wire [15:0] t1_r10_c10_rr3;
  wire [15:0] t1_r10_c10_rr4;
  wire [15:0] t1_r10_c10_rr5;
  wire [15:0] t1_r10_c10_rr6;
  wire [15:0] t1_r10_c10_rr7;
  wire [15:0] t2_r10_c10_rr0;
  wire [15:0] t2_r10_c10_rr1;
  wire [15:0] t2_r10_c10_rr2;
  wire [15:0] t2_r10_c10_rr3;
  wire [15:0] t3_r10_c10_rr0;
  wire [15:0] t3_r10_c10_rr1;
  wire [15:0] t4_r10_c10_rr0;
  wire [15:0] t0_r10_c11_rr0;
  wire [15:0] t0_r10_c11_rr1;
  wire [15:0] t0_r10_c11_rr2;
  wire [15:0] t0_r10_c11_rr3;
  wire [15:0] t0_r10_c11_rr4;
  wire [15:0] t0_r10_c11_rr5;
  wire [15:0] t0_r10_c11_rr6;
  wire [15:0] t0_r10_c11_rr7;
  wire [15:0] t0_r10_c11_rr8;
  wire [15:0] t0_r10_c11_rr9;
  wire [15:0] t0_r10_c11_rr10;
  wire [15:0] t0_r10_c11_rr11;
  wire [15:0] t0_r10_c11_rr12;
  wire [15:0] t0_r10_c11_rr13;
  wire [15:0] t0_r10_c11_rr14;
  wire [15:0] t1_r10_c11_rr0;
  wire [15:0] t1_r10_c11_rr1;
  wire [15:0] t1_r10_c11_rr2;
  wire [15:0] t1_r10_c11_rr3;
  wire [15:0] t1_r10_c11_rr4;
  wire [15:0] t1_r10_c11_rr5;
  wire [15:0] t1_r10_c11_rr6;
  wire [15:0] t1_r10_c11_rr7;
  wire [15:0] t2_r10_c11_rr0;
  wire [15:0] t2_r10_c11_rr1;
  wire [15:0] t2_r10_c11_rr2;
  wire [15:0] t2_r10_c11_rr3;
  wire [15:0] t3_r10_c11_rr0;
  wire [15:0] t3_r10_c11_rr1;
  wire [15:0] t4_r10_c11_rr0;
  wire [15:0] t0_r10_c12_rr0;
  wire [15:0] t0_r10_c12_rr1;
  wire [15:0] t0_r10_c12_rr2;
  wire [15:0] t0_r10_c12_rr3;
  wire [15:0] t0_r10_c12_rr4;
  wire [15:0] t0_r10_c12_rr5;
  wire [15:0] t0_r10_c12_rr6;
  wire [15:0] t0_r10_c12_rr7;
  wire [15:0] t0_r10_c12_rr8;
  wire [15:0] t0_r10_c12_rr9;
  wire [15:0] t0_r10_c12_rr10;
  wire [15:0] t0_r10_c12_rr11;
  wire [15:0] t0_r10_c12_rr12;
  wire [15:0] t0_r10_c12_rr13;
  wire [15:0] t0_r10_c12_rr14;
  wire [15:0] t1_r10_c12_rr0;
  wire [15:0] t1_r10_c12_rr1;
  wire [15:0] t1_r10_c12_rr2;
  wire [15:0] t1_r10_c12_rr3;
  wire [15:0] t1_r10_c12_rr4;
  wire [15:0] t1_r10_c12_rr5;
  wire [15:0] t1_r10_c12_rr6;
  wire [15:0] t1_r10_c12_rr7;
  wire [15:0] t2_r10_c12_rr0;
  wire [15:0] t2_r10_c12_rr1;
  wire [15:0] t2_r10_c12_rr2;
  wire [15:0] t2_r10_c12_rr3;
  wire [15:0] t3_r10_c12_rr0;
  wire [15:0] t3_r10_c12_rr1;
  wire [15:0] t4_r10_c12_rr0;
  wire [15:0] t0_r10_c13_rr0;
  wire [15:0] t0_r10_c13_rr1;
  wire [15:0] t0_r10_c13_rr2;
  wire [15:0] t0_r10_c13_rr3;
  wire [15:0] t0_r10_c13_rr4;
  wire [15:0] t0_r10_c13_rr5;
  wire [15:0] t0_r10_c13_rr6;
  wire [15:0] t0_r10_c13_rr7;
  wire [15:0] t0_r10_c13_rr8;
  wire [15:0] t0_r10_c13_rr9;
  wire [15:0] t0_r10_c13_rr10;
  wire [15:0] t0_r10_c13_rr11;
  wire [15:0] t0_r10_c13_rr12;
  wire [15:0] t0_r10_c13_rr13;
  wire [15:0] t0_r10_c13_rr14;
  wire [15:0] t1_r10_c13_rr0;
  wire [15:0] t1_r10_c13_rr1;
  wire [15:0] t1_r10_c13_rr2;
  wire [15:0] t1_r10_c13_rr3;
  wire [15:0] t1_r10_c13_rr4;
  wire [15:0] t1_r10_c13_rr5;
  wire [15:0] t1_r10_c13_rr6;
  wire [15:0] t1_r10_c13_rr7;
  wire [15:0] t2_r10_c13_rr0;
  wire [15:0] t2_r10_c13_rr1;
  wire [15:0] t2_r10_c13_rr2;
  wire [15:0] t2_r10_c13_rr3;
  wire [15:0] t3_r10_c13_rr0;
  wire [15:0] t3_r10_c13_rr1;
  wire [15:0] t4_r10_c13_rr0;
  wire [15:0] t0_r10_c14_rr0;
  wire [15:0] t0_r10_c14_rr1;
  wire [15:0] t0_r10_c14_rr2;
  wire [15:0] t0_r10_c14_rr3;
  wire [15:0] t0_r10_c14_rr4;
  wire [15:0] t0_r10_c14_rr5;
  wire [15:0] t0_r10_c14_rr6;
  wire [15:0] t0_r10_c14_rr7;
  wire [15:0] t0_r10_c14_rr8;
  wire [15:0] t0_r10_c14_rr9;
  wire [15:0] t0_r10_c14_rr10;
  wire [15:0] t0_r10_c14_rr11;
  wire [15:0] t0_r10_c14_rr12;
  wire [15:0] t0_r10_c14_rr13;
  wire [15:0] t0_r10_c14_rr14;
  wire [15:0] t1_r10_c14_rr0;
  wire [15:0] t1_r10_c14_rr1;
  wire [15:0] t1_r10_c14_rr2;
  wire [15:0] t1_r10_c14_rr3;
  wire [15:0] t1_r10_c14_rr4;
  wire [15:0] t1_r10_c14_rr5;
  wire [15:0] t1_r10_c14_rr6;
  wire [15:0] t1_r10_c14_rr7;
  wire [15:0] t2_r10_c14_rr0;
  wire [15:0] t2_r10_c14_rr1;
  wire [15:0] t2_r10_c14_rr2;
  wire [15:0] t2_r10_c14_rr3;
  wire [15:0] t3_r10_c14_rr0;
  wire [15:0] t3_r10_c14_rr1;
  wire [15:0] t4_r10_c14_rr0;
  wire [15:0] t0_r11_c0_rr0;
  wire [15:0] t0_r11_c0_rr1;
  wire [15:0] t0_r11_c0_rr2;
  wire [15:0] t0_r11_c0_rr3;
  wire [15:0] t0_r11_c0_rr4;
  wire [15:0] t0_r11_c0_rr5;
  wire [15:0] t0_r11_c0_rr6;
  wire [15:0] t0_r11_c0_rr7;
  wire [15:0] t0_r11_c0_rr8;
  wire [15:0] t0_r11_c0_rr9;
  wire [15:0] t0_r11_c0_rr10;
  wire [15:0] t0_r11_c0_rr11;
  wire [15:0] t0_r11_c0_rr12;
  wire [15:0] t0_r11_c0_rr13;
  wire [15:0] t0_r11_c0_rr14;
  wire [15:0] t1_r11_c0_rr0;
  wire [15:0] t1_r11_c0_rr1;
  wire [15:0] t1_r11_c0_rr2;
  wire [15:0] t1_r11_c0_rr3;
  wire [15:0] t1_r11_c0_rr4;
  wire [15:0] t1_r11_c0_rr5;
  wire [15:0] t1_r11_c0_rr6;
  wire [15:0] t1_r11_c0_rr7;
  wire [15:0] t2_r11_c0_rr0;
  wire [15:0] t2_r11_c0_rr1;
  wire [15:0] t2_r11_c0_rr2;
  wire [15:0] t2_r11_c0_rr3;
  wire [15:0] t3_r11_c0_rr0;
  wire [15:0] t3_r11_c0_rr1;
  wire [15:0] t4_r11_c0_rr0;
  wire [15:0] t0_r11_c1_rr0;
  wire [15:0] t0_r11_c1_rr1;
  wire [15:0] t0_r11_c1_rr2;
  wire [15:0] t0_r11_c1_rr3;
  wire [15:0] t0_r11_c1_rr4;
  wire [15:0] t0_r11_c1_rr5;
  wire [15:0] t0_r11_c1_rr6;
  wire [15:0] t0_r11_c1_rr7;
  wire [15:0] t0_r11_c1_rr8;
  wire [15:0] t0_r11_c1_rr9;
  wire [15:0] t0_r11_c1_rr10;
  wire [15:0] t0_r11_c1_rr11;
  wire [15:0] t0_r11_c1_rr12;
  wire [15:0] t0_r11_c1_rr13;
  wire [15:0] t0_r11_c1_rr14;
  wire [15:0] t1_r11_c1_rr0;
  wire [15:0] t1_r11_c1_rr1;
  wire [15:0] t1_r11_c1_rr2;
  wire [15:0] t1_r11_c1_rr3;
  wire [15:0] t1_r11_c1_rr4;
  wire [15:0] t1_r11_c1_rr5;
  wire [15:0] t1_r11_c1_rr6;
  wire [15:0] t1_r11_c1_rr7;
  wire [15:0] t2_r11_c1_rr0;
  wire [15:0] t2_r11_c1_rr1;
  wire [15:0] t2_r11_c1_rr2;
  wire [15:0] t2_r11_c1_rr3;
  wire [15:0] t3_r11_c1_rr0;
  wire [15:0] t3_r11_c1_rr1;
  wire [15:0] t4_r11_c1_rr0;
  wire [15:0] t0_r11_c2_rr0;
  wire [15:0] t0_r11_c2_rr1;
  wire [15:0] t0_r11_c2_rr2;
  wire [15:0] t0_r11_c2_rr3;
  wire [15:0] t0_r11_c2_rr4;
  wire [15:0] t0_r11_c2_rr5;
  wire [15:0] t0_r11_c2_rr6;
  wire [15:0] t0_r11_c2_rr7;
  wire [15:0] t0_r11_c2_rr8;
  wire [15:0] t0_r11_c2_rr9;
  wire [15:0] t0_r11_c2_rr10;
  wire [15:0] t0_r11_c2_rr11;
  wire [15:0] t0_r11_c2_rr12;
  wire [15:0] t0_r11_c2_rr13;
  wire [15:0] t0_r11_c2_rr14;
  wire [15:0] t1_r11_c2_rr0;
  wire [15:0] t1_r11_c2_rr1;
  wire [15:0] t1_r11_c2_rr2;
  wire [15:0] t1_r11_c2_rr3;
  wire [15:0] t1_r11_c2_rr4;
  wire [15:0] t1_r11_c2_rr5;
  wire [15:0] t1_r11_c2_rr6;
  wire [15:0] t1_r11_c2_rr7;
  wire [15:0] t2_r11_c2_rr0;
  wire [15:0] t2_r11_c2_rr1;
  wire [15:0] t2_r11_c2_rr2;
  wire [15:0] t2_r11_c2_rr3;
  wire [15:0] t3_r11_c2_rr0;
  wire [15:0] t3_r11_c2_rr1;
  wire [15:0] t4_r11_c2_rr0;
  wire [15:0] t0_r11_c3_rr0;
  wire [15:0] t0_r11_c3_rr1;
  wire [15:0] t0_r11_c3_rr2;
  wire [15:0] t0_r11_c3_rr3;
  wire [15:0] t0_r11_c3_rr4;
  wire [15:0] t0_r11_c3_rr5;
  wire [15:0] t0_r11_c3_rr6;
  wire [15:0] t0_r11_c3_rr7;
  wire [15:0] t0_r11_c3_rr8;
  wire [15:0] t0_r11_c3_rr9;
  wire [15:0] t0_r11_c3_rr10;
  wire [15:0] t0_r11_c3_rr11;
  wire [15:0] t0_r11_c3_rr12;
  wire [15:0] t0_r11_c3_rr13;
  wire [15:0] t0_r11_c3_rr14;
  wire [15:0] t1_r11_c3_rr0;
  wire [15:0] t1_r11_c3_rr1;
  wire [15:0] t1_r11_c3_rr2;
  wire [15:0] t1_r11_c3_rr3;
  wire [15:0] t1_r11_c3_rr4;
  wire [15:0] t1_r11_c3_rr5;
  wire [15:0] t1_r11_c3_rr6;
  wire [15:0] t1_r11_c3_rr7;
  wire [15:0] t2_r11_c3_rr0;
  wire [15:0] t2_r11_c3_rr1;
  wire [15:0] t2_r11_c3_rr2;
  wire [15:0] t2_r11_c3_rr3;
  wire [15:0] t3_r11_c3_rr0;
  wire [15:0] t3_r11_c3_rr1;
  wire [15:0] t4_r11_c3_rr0;
  wire [15:0] t0_r11_c4_rr0;
  wire [15:0] t0_r11_c4_rr1;
  wire [15:0] t0_r11_c4_rr2;
  wire [15:0] t0_r11_c4_rr3;
  wire [15:0] t0_r11_c4_rr4;
  wire [15:0] t0_r11_c4_rr5;
  wire [15:0] t0_r11_c4_rr6;
  wire [15:0] t0_r11_c4_rr7;
  wire [15:0] t0_r11_c4_rr8;
  wire [15:0] t0_r11_c4_rr9;
  wire [15:0] t0_r11_c4_rr10;
  wire [15:0] t0_r11_c4_rr11;
  wire [15:0] t0_r11_c4_rr12;
  wire [15:0] t0_r11_c4_rr13;
  wire [15:0] t0_r11_c4_rr14;
  wire [15:0] t1_r11_c4_rr0;
  wire [15:0] t1_r11_c4_rr1;
  wire [15:0] t1_r11_c4_rr2;
  wire [15:0] t1_r11_c4_rr3;
  wire [15:0] t1_r11_c4_rr4;
  wire [15:0] t1_r11_c4_rr5;
  wire [15:0] t1_r11_c4_rr6;
  wire [15:0] t1_r11_c4_rr7;
  wire [15:0] t2_r11_c4_rr0;
  wire [15:0] t2_r11_c4_rr1;
  wire [15:0] t2_r11_c4_rr2;
  wire [15:0] t2_r11_c4_rr3;
  wire [15:0] t3_r11_c4_rr0;
  wire [15:0] t3_r11_c4_rr1;
  wire [15:0] t4_r11_c4_rr0;
  wire [15:0] t0_r11_c5_rr0;
  wire [15:0] t0_r11_c5_rr1;
  wire [15:0] t0_r11_c5_rr2;
  wire [15:0] t0_r11_c5_rr3;
  wire [15:0] t0_r11_c5_rr4;
  wire [15:0] t0_r11_c5_rr5;
  wire [15:0] t0_r11_c5_rr6;
  wire [15:0] t0_r11_c5_rr7;
  wire [15:0] t0_r11_c5_rr8;
  wire [15:0] t0_r11_c5_rr9;
  wire [15:0] t0_r11_c5_rr10;
  wire [15:0] t0_r11_c5_rr11;
  wire [15:0] t0_r11_c5_rr12;
  wire [15:0] t0_r11_c5_rr13;
  wire [15:0] t0_r11_c5_rr14;
  wire [15:0] t1_r11_c5_rr0;
  wire [15:0] t1_r11_c5_rr1;
  wire [15:0] t1_r11_c5_rr2;
  wire [15:0] t1_r11_c5_rr3;
  wire [15:0] t1_r11_c5_rr4;
  wire [15:0] t1_r11_c5_rr5;
  wire [15:0] t1_r11_c5_rr6;
  wire [15:0] t1_r11_c5_rr7;
  wire [15:0] t2_r11_c5_rr0;
  wire [15:0] t2_r11_c5_rr1;
  wire [15:0] t2_r11_c5_rr2;
  wire [15:0] t2_r11_c5_rr3;
  wire [15:0] t3_r11_c5_rr0;
  wire [15:0] t3_r11_c5_rr1;
  wire [15:0] t4_r11_c5_rr0;
  wire [15:0] t0_r11_c6_rr0;
  wire [15:0] t0_r11_c6_rr1;
  wire [15:0] t0_r11_c6_rr2;
  wire [15:0] t0_r11_c6_rr3;
  wire [15:0] t0_r11_c6_rr4;
  wire [15:0] t0_r11_c6_rr5;
  wire [15:0] t0_r11_c6_rr6;
  wire [15:0] t0_r11_c6_rr7;
  wire [15:0] t0_r11_c6_rr8;
  wire [15:0] t0_r11_c6_rr9;
  wire [15:0] t0_r11_c6_rr10;
  wire [15:0] t0_r11_c6_rr11;
  wire [15:0] t0_r11_c6_rr12;
  wire [15:0] t0_r11_c6_rr13;
  wire [15:0] t0_r11_c6_rr14;
  wire [15:0] t1_r11_c6_rr0;
  wire [15:0] t1_r11_c6_rr1;
  wire [15:0] t1_r11_c6_rr2;
  wire [15:0] t1_r11_c6_rr3;
  wire [15:0] t1_r11_c6_rr4;
  wire [15:0] t1_r11_c6_rr5;
  wire [15:0] t1_r11_c6_rr6;
  wire [15:0] t1_r11_c6_rr7;
  wire [15:0] t2_r11_c6_rr0;
  wire [15:0] t2_r11_c6_rr1;
  wire [15:0] t2_r11_c6_rr2;
  wire [15:0] t2_r11_c6_rr3;
  wire [15:0] t3_r11_c6_rr0;
  wire [15:0] t3_r11_c6_rr1;
  wire [15:0] t4_r11_c6_rr0;
  wire [15:0] t0_r11_c7_rr0;
  wire [15:0] t0_r11_c7_rr1;
  wire [15:0] t0_r11_c7_rr2;
  wire [15:0] t0_r11_c7_rr3;
  wire [15:0] t0_r11_c7_rr4;
  wire [15:0] t0_r11_c7_rr5;
  wire [15:0] t0_r11_c7_rr6;
  wire [15:0] t0_r11_c7_rr7;
  wire [15:0] t0_r11_c7_rr8;
  wire [15:0] t0_r11_c7_rr9;
  wire [15:0] t0_r11_c7_rr10;
  wire [15:0] t0_r11_c7_rr11;
  wire [15:0] t0_r11_c7_rr12;
  wire [15:0] t0_r11_c7_rr13;
  wire [15:0] t0_r11_c7_rr14;
  wire [15:0] t1_r11_c7_rr0;
  wire [15:0] t1_r11_c7_rr1;
  wire [15:0] t1_r11_c7_rr2;
  wire [15:0] t1_r11_c7_rr3;
  wire [15:0] t1_r11_c7_rr4;
  wire [15:0] t1_r11_c7_rr5;
  wire [15:0] t1_r11_c7_rr6;
  wire [15:0] t1_r11_c7_rr7;
  wire [15:0] t2_r11_c7_rr0;
  wire [15:0] t2_r11_c7_rr1;
  wire [15:0] t2_r11_c7_rr2;
  wire [15:0] t2_r11_c7_rr3;
  wire [15:0] t3_r11_c7_rr0;
  wire [15:0] t3_r11_c7_rr1;
  wire [15:0] t4_r11_c7_rr0;
  wire [15:0] t0_r11_c8_rr0;
  wire [15:0] t0_r11_c8_rr1;
  wire [15:0] t0_r11_c8_rr2;
  wire [15:0] t0_r11_c8_rr3;
  wire [15:0] t0_r11_c8_rr4;
  wire [15:0] t0_r11_c8_rr5;
  wire [15:0] t0_r11_c8_rr6;
  wire [15:0] t0_r11_c8_rr7;
  wire [15:0] t0_r11_c8_rr8;
  wire [15:0] t0_r11_c8_rr9;
  wire [15:0] t0_r11_c8_rr10;
  wire [15:0] t0_r11_c8_rr11;
  wire [15:0] t0_r11_c8_rr12;
  wire [15:0] t0_r11_c8_rr13;
  wire [15:0] t0_r11_c8_rr14;
  wire [15:0] t1_r11_c8_rr0;
  wire [15:0] t1_r11_c8_rr1;
  wire [15:0] t1_r11_c8_rr2;
  wire [15:0] t1_r11_c8_rr3;
  wire [15:0] t1_r11_c8_rr4;
  wire [15:0] t1_r11_c8_rr5;
  wire [15:0] t1_r11_c8_rr6;
  wire [15:0] t1_r11_c8_rr7;
  wire [15:0] t2_r11_c8_rr0;
  wire [15:0] t2_r11_c8_rr1;
  wire [15:0] t2_r11_c8_rr2;
  wire [15:0] t2_r11_c8_rr3;
  wire [15:0] t3_r11_c8_rr0;
  wire [15:0] t3_r11_c8_rr1;
  wire [15:0] t4_r11_c8_rr0;
  wire [15:0] t0_r11_c9_rr0;
  wire [15:0] t0_r11_c9_rr1;
  wire [15:0] t0_r11_c9_rr2;
  wire [15:0] t0_r11_c9_rr3;
  wire [15:0] t0_r11_c9_rr4;
  wire [15:0] t0_r11_c9_rr5;
  wire [15:0] t0_r11_c9_rr6;
  wire [15:0] t0_r11_c9_rr7;
  wire [15:0] t0_r11_c9_rr8;
  wire [15:0] t0_r11_c9_rr9;
  wire [15:0] t0_r11_c9_rr10;
  wire [15:0] t0_r11_c9_rr11;
  wire [15:0] t0_r11_c9_rr12;
  wire [15:0] t0_r11_c9_rr13;
  wire [15:0] t0_r11_c9_rr14;
  wire [15:0] t1_r11_c9_rr0;
  wire [15:0] t1_r11_c9_rr1;
  wire [15:0] t1_r11_c9_rr2;
  wire [15:0] t1_r11_c9_rr3;
  wire [15:0] t1_r11_c9_rr4;
  wire [15:0] t1_r11_c9_rr5;
  wire [15:0] t1_r11_c9_rr6;
  wire [15:0] t1_r11_c9_rr7;
  wire [15:0] t2_r11_c9_rr0;
  wire [15:0] t2_r11_c9_rr1;
  wire [15:0] t2_r11_c9_rr2;
  wire [15:0] t2_r11_c9_rr3;
  wire [15:0] t3_r11_c9_rr0;
  wire [15:0] t3_r11_c9_rr1;
  wire [15:0] t4_r11_c9_rr0;
  wire [15:0] t0_r11_c10_rr0;
  wire [15:0] t0_r11_c10_rr1;
  wire [15:0] t0_r11_c10_rr2;
  wire [15:0] t0_r11_c10_rr3;
  wire [15:0] t0_r11_c10_rr4;
  wire [15:0] t0_r11_c10_rr5;
  wire [15:0] t0_r11_c10_rr6;
  wire [15:0] t0_r11_c10_rr7;
  wire [15:0] t0_r11_c10_rr8;
  wire [15:0] t0_r11_c10_rr9;
  wire [15:0] t0_r11_c10_rr10;
  wire [15:0] t0_r11_c10_rr11;
  wire [15:0] t0_r11_c10_rr12;
  wire [15:0] t0_r11_c10_rr13;
  wire [15:0] t0_r11_c10_rr14;
  wire [15:0] t1_r11_c10_rr0;
  wire [15:0] t1_r11_c10_rr1;
  wire [15:0] t1_r11_c10_rr2;
  wire [15:0] t1_r11_c10_rr3;
  wire [15:0] t1_r11_c10_rr4;
  wire [15:0] t1_r11_c10_rr5;
  wire [15:0] t1_r11_c10_rr6;
  wire [15:0] t1_r11_c10_rr7;
  wire [15:0] t2_r11_c10_rr0;
  wire [15:0] t2_r11_c10_rr1;
  wire [15:0] t2_r11_c10_rr2;
  wire [15:0] t2_r11_c10_rr3;
  wire [15:0] t3_r11_c10_rr0;
  wire [15:0] t3_r11_c10_rr1;
  wire [15:0] t4_r11_c10_rr0;
  wire [15:0] t0_r11_c11_rr0;
  wire [15:0] t0_r11_c11_rr1;
  wire [15:0] t0_r11_c11_rr2;
  wire [15:0] t0_r11_c11_rr3;
  wire [15:0] t0_r11_c11_rr4;
  wire [15:0] t0_r11_c11_rr5;
  wire [15:0] t0_r11_c11_rr6;
  wire [15:0] t0_r11_c11_rr7;
  wire [15:0] t0_r11_c11_rr8;
  wire [15:0] t0_r11_c11_rr9;
  wire [15:0] t0_r11_c11_rr10;
  wire [15:0] t0_r11_c11_rr11;
  wire [15:0] t0_r11_c11_rr12;
  wire [15:0] t0_r11_c11_rr13;
  wire [15:0] t0_r11_c11_rr14;
  wire [15:0] t1_r11_c11_rr0;
  wire [15:0] t1_r11_c11_rr1;
  wire [15:0] t1_r11_c11_rr2;
  wire [15:0] t1_r11_c11_rr3;
  wire [15:0] t1_r11_c11_rr4;
  wire [15:0] t1_r11_c11_rr5;
  wire [15:0] t1_r11_c11_rr6;
  wire [15:0] t1_r11_c11_rr7;
  wire [15:0] t2_r11_c11_rr0;
  wire [15:0] t2_r11_c11_rr1;
  wire [15:0] t2_r11_c11_rr2;
  wire [15:0] t2_r11_c11_rr3;
  wire [15:0] t3_r11_c11_rr0;
  wire [15:0] t3_r11_c11_rr1;
  wire [15:0] t4_r11_c11_rr0;
  wire [15:0] t0_r11_c12_rr0;
  wire [15:0] t0_r11_c12_rr1;
  wire [15:0] t0_r11_c12_rr2;
  wire [15:0] t0_r11_c12_rr3;
  wire [15:0] t0_r11_c12_rr4;
  wire [15:0] t0_r11_c12_rr5;
  wire [15:0] t0_r11_c12_rr6;
  wire [15:0] t0_r11_c12_rr7;
  wire [15:0] t0_r11_c12_rr8;
  wire [15:0] t0_r11_c12_rr9;
  wire [15:0] t0_r11_c12_rr10;
  wire [15:0] t0_r11_c12_rr11;
  wire [15:0] t0_r11_c12_rr12;
  wire [15:0] t0_r11_c12_rr13;
  wire [15:0] t0_r11_c12_rr14;
  wire [15:0] t1_r11_c12_rr0;
  wire [15:0] t1_r11_c12_rr1;
  wire [15:0] t1_r11_c12_rr2;
  wire [15:0] t1_r11_c12_rr3;
  wire [15:0] t1_r11_c12_rr4;
  wire [15:0] t1_r11_c12_rr5;
  wire [15:0] t1_r11_c12_rr6;
  wire [15:0] t1_r11_c12_rr7;
  wire [15:0] t2_r11_c12_rr0;
  wire [15:0] t2_r11_c12_rr1;
  wire [15:0] t2_r11_c12_rr2;
  wire [15:0] t2_r11_c12_rr3;
  wire [15:0] t3_r11_c12_rr0;
  wire [15:0] t3_r11_c12_rr1;
  wire [15:0] t4_r11_c12_rr0;
  wire [15:0] t0_r11_c13_rr0;
  wire [15:0] t0_r11_c13_rr1;
  wire [15:0] t0_r11_c13_rr2;
  wire [15:0] t0_r11_c13_rr3;
  wire [15:0] t0_r11_c13_rr4;
  wire [15:0] t0_r11_c13_rr5;
  wire [15:0] t0_r11_c13_rr6;
  wire [15:0] t0_r11_c13_rr7;
  wire [15:0] t0_r11_c13_rr8;
  wire [15:0] t0_r11_c13_rr9;
  wire [15:0] t0_r11_c13_rr10;
  wire [15:0] t0_r11_c13_rr11;
  wire [15:0] t0_r11_c13_rr12;
  wire [15:0] t0_r11_c13_rr13;
  wire [15:0] t0_r11_c13_rr14;
  wire [15:0] t1_r11_c13_rr0;
  wire [15:0] t1_r11_c13_rr1;
  wire [15:0] t1_r11_c13_rr2;
  wire [15:0] t1_r11_c13_rr3;
  wire [15:0] t1_r11_c13_rr4;
  wire [15:0] t1_r11_c13_rr5;
  wire [15:0] t1_r11_c13_rr6;
  wire [15:0] t1_r11_c13_rr7;
  wire [15:0] t2_r11_c13_rr0;
  wire [15:0] t2_r11_c13_rr1;
  wire [15:0] t2_r11_c13_rr2;
  wire [15:0] t2_r11_c13_rr3;
  wire [15:0] t3_r11_c13_rr0;
  wire [15:0] t3_r11_c13_rr1;
  wire [15:0] t4_r11_c13_rr0;
  wire [15:0] t0_r11_c14_rr0;
  wire [15:0] t0_r11_c14_rr1;
  wire [15:0] t0_r11_c14_rr2;
  wire [15:0] t0_r11_c14_rr3;
  wire [15:0] t0_r11_c14_rr4;
  wire [15:0] t0_r11_c14_rr5;
  wire [15:0] t0_r11_c14_rr6;
  wire [15:0] t0_r11_c14_rr7;
  wire [15:0] t0_r11_c14_rr8;
  wire [15:0] t0_r11_c14_rr9;
  wire [15:0] t0_r11_c14_rr10;
  wire [15:0] t0_r11_c14_rr11;
  wire [15:0] t0_r11_c14_rr12;
  wire [15:0] t0_r11_c14_rr13;
  wire [15:0] t0_r11_c14_rr14;
  wire [15:0] t1_r11_c14_rr0;
  wire [15:0] t1_r11_c14_rr1;
  wire [15:0] t1_r11_c14_rr2;
  wire [15:0] t1_r11_c14_rr3;
  wire [15:0] t1_r11_c14_rr4;
  wire [15:0] t1_r11_c14_rr5;
  wire [15:0] t1_r11_c14_rr6;
  wire [15:0] t1_r11_c14_rr7;
  wire [15:0] t2_r11_c14_rr0;
  wire [15:0] t2_r11_c14_rr1;
  wire [15:0] t2_r11_c14_rr2;
  wire [15:0] t2_r11_c14_rr3;
  wire [15:0] t3_r11_c14_rr0;
  wire [15:0] t3_r11_c14_rr1;
  wire [15:0] t4_r11_c14_rr0;
  wire [15:0] t0_r12_c0_rr0;
  wire [15:0] t0_r12_c0_rr1;
  wire [15:0] t0_r12_c0_rr2;
  wire [15:0] t0_r12_c0_rr3;
  wire [15:0] t0_r12_c0_rr4;
  wire [15:0] t0_r12_c0_rr5;
  wire [15:0] t0_r12_c0_rr6;
  wire [15:0] t0_r12_c0_rr7;
  wire [15:0] t0_r12_c0_rr8;
  wire [15:0] t0_r12_c0_rr9;
  wire [15:0] t0_r12_c0_rr10;
  wire [15:0] t0_r12_c0_rr11;
  wire [15:0] t0_r12_c0_rr12;
  wire [15:0] t0_r12_c0_rr13;
  wire [15:0] t0_r12_c0_rr14;
  wire [15:0] t1_r12_c0_rr0;
  wire [15:0] t1_r12_c0_rr1;
  wire [15:0] t1_r12_c0_rr2;
  wire [15:0] t1_r12_c0_rr3;
  wire [15:0] t1_r12_c0_rr4;
  wire [15:0] t1_r12_c0_rr5;
  wire [15:0] t1_r12_c0_rr6;
  wire [15:0] t1_r12_c0_rr7;
  wire [15:0] t2_r12_c0_rr0;
  wire [15:0] t2_r12_c0_rr1;
  wire [15:0] t2_r12_c0_rr2;
  wire [15:0] t2_r12_c0_rr3;
  wire [15:0] t3_r12_c0_rr0;
  wire [15:0] t3_r12_c0_rr1;
  wire [15:0] t4_r12_c0_rr0;
  wire [15:0] t0_r12_c1_rr0;
  wire [15:0] t0_r12_c1_rr1;
  wire [15:0] t0_r12_c1_rr2;
  wire [15:0] t0_r12_c1_rr3;
  wire [15:0] t0_r12_c1_rr4;
  wire [15:0] t0_r12_c1_rr5;
  wire [15:0] t0_r12_c1_rr6;
  wire [15:0] t0_r12_c1_rr7;
  wire [15:0] t0_r12_c1_rr8;
  wire [15:0] t0_r12_c1_rr9;
  wire [15:0] t0_r12_c1_rr10;
  wire [15:0] t0_r12_c1_rr11;
  wire [15:0] t0_r12_c1_rr12;
  wire [15:0] t0_r12_c1_rr13;
  wire [15:0] t0_r12_c1_rr14;
  wire [15:0] t1_r12_c1_rr0;
  wire [15:0] t1_r12_c1_rr1;
  wire [15:0] t1_r12_c1_rr2;
  wire [15:0] t1_r12_c1_rr3;
  wire [15:0] t1_r12_c1_rr4;
  wire [15:0] t1_r12_c1_rr5;
  wire [15:0] t1_r12_c1_rr6;
  wire [15:0] t1_r12_c1_rr7;
  wire [15:0] t2_r12_c1_rr0;
  wire [15:0] t2_r12_c1_rr1;
  wire [15:0] t2_r12_c1_rr2;
  wire [15:0] t2_r12_c1_rr3;
  wire [15:0] t3_r12_c1_rr0;
  wire [15:0] t3_r12_c1_rr1;
  wire [15:0] t4_r12_c1_rr0;
  wire [15:0] t0_r12_c2_rr0;
  wire [15:0] t0_r12_c2_rr1;
  wire [15:0] t0_r12_c2_rr2;
  wire [15:0] t0_r12_c2_rr3;
  wire [15:0] t0_r12_c2_rr4;
  wire [15:0] t0_r12_c2_rr5;
  wire [15:0] t0_r12_c2_rr6;
  wire [15:0] t0_r12_c2_rr7;
  wire [15:0] t0_r12_c2_rr8;
  wire [15:0] t0_r12_c2_rr9;
  wire [15:0] t0_r12_c2_rr10;
  wire [15:0] t0_r12_c2_rr11;
  wire [15:0] t0_r12_c2_rr12;
  wire [15:0] t0_r12_c2_rr13;
  wire [15:0] t0_r12_c2_rr14;
  wire [15:0] t1_r12_c2_rr0;
  wire [15:0] t1_r12_c2_rr1;
  wire [15:0] t1_r12_c2_rr2;
  wire [15:0] t1_r12_c2_rr3;
  wire [15:0] t1_r12_c2_rr4;
  wire [15:0] t1_r12_c2_rr5;
  wire [15:0] t1_r12_c2_rr6;
  wire [15:0] t1_r12_c2_rr7;
  wire [15:0] t2_r12_c2_rr0;
  wire [15:0] t2_r12_c2_rr1;
  wire [15:0] t2_r12_c2_rr2;
  wire [15:0] t2_r12_c2_rr3;
  wire [15:0] t3_r12_c2_rr0;
  wire [15:0] t3_r12_c2_rr1;
  wire [15:0] t4_r12_c2_rr0;
  wire [15:0] t0_r12_c3_rr0;
  wire [15:0] t0_r12_c3_rr1;
  wire [15:0] t0_r12_c3_rr2;
  wire [15:0] t0_r12_c3_rr3;
  wire [15:0] t0_r12_c3_rr4;
  wire [15:0] t0_r12_c3_rr5;
  wire [15:0] t0_r12_c3_rr6;
  wire [15:0] t0_r12_c3_rr7;
  wire [15:0] t0_r12_c3_rr8;
  wire [15:0] t0_r12_c3_rr9;
  wire [15:0] t0_r12_c3_rr10;
  wire [15:0] t0_r12_c3_rr11;
  wire [15:0] t0_r12_c3_rr12;
  wire [15:0] t0_r12_c3_rr13;
  wire [15:0] t0_r12_c3_rr14;
  wire [15:0] t1_r12_c3_rr0;
  wire [15:0] t1_r12_c3_rr1;
  wire [15:0] t1_r12_c3_rr2;
  wire [15:0] t1_r12_c3_rr3;
  wire [15:0] t1_r12_c3_rr4;
  wire [15:0] t1_r12_c3_rr5;
  wire [15:0] t1_r12_c3_rr6;
  wire [15:0] t1_r12_c3_rr7;
  wire [15:0] t2_r12_c3_rr0;
  wire [15:0] t2_r12_c3_rr1;
  wire [15:0] t2_r12_c3_rr2;
  wire [15:0] t2_r12_c3_rr3;
  wire [15:0] t3_r12_c3_rr0;
  wire [15:0] t3_r12_c3_rr1;
  wire [15:0] t4_r12_c3_rr0;
  wire [15:0] t0_r12_c4_rr0;
  wire [15:0] t0_r12_c4_rr1;
  wire [15:0] t0_r12_c4_rr2;
  wire [15:0] t0_r12_c4_rr3;
  wire [15:0] t0_r12_c4_rr4;
  wire [15:0] t0_r12_c4_rr5;
  wire [15:0] t0_r12_c4_rr6;
  wire [15:0] t0_r12_c4_rr7;
  wire [15:0] t0_r12_c4_rr8;
  wire [15:0] t0_r12_c4_rr9;
  wire [15:0] t0_r12_c4_rr10;
  wire [15:0] t0_r12_c4_rr11;
  wire [15:0] t0_r12_c4_rr12;
  wire [15:0] t0_r12_c4_rr13;
  wire [15:0] t0_r12_c4_rr14;
  wire [15:0] t1_r12_c4_rr0;
  wire [15:0] t1_r12_c4_rr1;
  wire [15:0] t1_r12_c4_rr2;
  wire [15:0] t1_r12_c4_rr3;
  wire [15:0] t1_r12_c4_rr4;
  wire [15:0] t1_r12_c4_rr5;
  wire [15:0] t1_r12_c4_rr6;
  wire [15:0] t1_r12_c4_rr7;
  wire [15:0] t2_r12_c4_rr0;
  wire [15:0] t2_r12_c4_rr1;
  wire [15:0] t2_r12_c4_rr2;
  wire [15:0] t2_r12_c4_rr3;
  wire [15:0] t3_r12_c4_rr0;
  wire [15:0] t3_r12_c4_rr1;
  wire [15:0] t4_r12_c4_rr0;
  wire [15:0] t0_r12_c5_rr0;
  wire [15:0] t0_r12_c5_rr1;
  wire [15:0] t0_r12_c5_rr2;
  wire [15:0] t0_r12_c5_rr3;
  wire [15:0] t0_r12_c5_rr4;
  wire [15:0] t0_r12_c5_rr5;
  wire [15:0] t0_r12_c5_rr6;
  wire [15:0] t0_r12_c5_rr7;
  wire [15:0] t0_r12_c5_rr8;
  wire [15:0] t0_r12_c5_rr9;
  wire [15:0] t0_r12_c5_rr10;
  wire [15:0] t0_r12_c5_rr11;
  wire [15:0] t0_r12_c5_rr12;
  wire [15:0] t0_r12_c5_rr13;
  wire [15:0] t0_r12_c5_rr14;
  wire [15:0] t1_r12_c5_rr0;
  wire [15:0] t1_r12_c5_rr1;
  wire [15:0] t1_r12_c5_rr2;
  wire [15:0] t1_r12_c5_rr3;
  wire [15:0] t1_r12_c5_rr4;
  wire [15:0] t1_r12_c5_rr5;
  wire [15:0] t1_r12_c5_rr6;
  wire [15:0] t1_r12_c5_rr7;
  wire [15:0] t2_r12_c5_rr0;
  wire [15:0] t2_r12_c5_rr1;
  wire [15:0] t2_r12_c5_rr2;
  wire [15:0] t2_r12_c5_rr3;
  wire [15:0] t3_r12_c5_rr0;
  wire [15:0] t3_r12_c5_rr1;
  wire [15:0] t4_r12_c5_rr0;
  wire [15:0] t0_r12_c6_rr0;
  wire [15:0] t0_r12_c6_rr1;
  wire [15:0] t0_r12_c6_rr2;
  wire [15:0] t0_r12_c6_rr3;
  wire [15:0] t0_r12_c6_rr4;
  wire [15:0] t0_r12_c6_rr5;
  wire [15:0] t0_r12_c6_rr6;
  wire [15:0] t0_r12_c6_rr7;
  wire [15:0] t0_r12_c6_rr8;
  wire [15:0] t0_r12_c6_rr9;
  wire [15:0] t0_r12_c6_rr10;
  wire [15:0] t0_r12_c6_rr11;
  wire [15:0] t0_r12_c6_rr12;
  wire [15:0] t0_r12_c6_rr13;
  wire [15:0] t0_r12_c6_rr14;
  wire [15:0] t1_r12_c6_rr0;
  wire [15:0] t1_r12_c6_rr1;
  wire [15:0] t1_r12_c6_rr2;
  wire [15:0] t1_r12_c6_rr3;
  wire [15:0] t1_r12_c6_rr4;
  wire [15:0] t1_r12_c6_rr5;
  wire [15:0] t1_r12_c6_rr6;
  wire [15:0] t1_r12_c6_rr7;
  wire [15:0] t2_r12_c6_rr0;
  wire [15:0] t2_r12_c6_rr1;
  wire [15:0] t2_r12_c6_rr2;
  wire [15:0] t2_r12_c6_rr3;
  wire [15:0] t3_r12_c6_rr0;
  wire [15:0] t3_r12_c6_rr1;
  wire [15:0] t4_r12_c6_rr0;
  wire [15:0] t0_r12_c7_rr0;
  wire [15:0] t0_r12_c7_rr1;
  wire [15:0] t0_r12_c7_rr2;
  wire [15:0] t0_r12_c7_rr3;
  wire [15:0] t0_r12_c7_rr4;
  wire [15:0] t0_r12_c7_rr5;
  wire [15:0] t0_r12_c7_rr6;
  wire [15:0] t0_r12_c7_rr7;
  wire [15:0] t0_r12_c7_rr8;
  wire [15:0] t0_r12_c7_rr9;
  wire [15:0] t0_r12_c7_rr10;
  wire [15:0] t0_r12_c7_rr11;
  wire [15:0] t0_r12_c7_rr12;
  wire [15:0] t0_r12_c7_rr13;
  wire [15:0] t0_r12_c7_rr14;
  wire [15:0] t1_r12_c7_rr0;
  wire [15:0] t1_r12_c7_rr1;
  wire [15:0] t1_r12_c7_rr2;
  wire [15:0] t1_r12_c7_rr3;
  wire [15:0] t1_r12_c7_rr4;
  wire [15:0] t1_r12_c7_rr5;
  wire [15:0] t1_r12_c7_rr6;
  wire [15:0] t1_r12_c7_rr7;
  wire [15:0] t2_r12_c7_rr0;
  wire [15:0] t2_r12_c7_rr1;
  wire [15:0] t2_r12_c7_rr2;
  wire [15:0] t2_r12_c7_rr3;
  wire [15:0] t3_r12_c7_rr0;
  wire [15:0] t3_r12_c7_rr1;
  wire [15:0] t4_r12_c7_rr0;
  wire [15:0] t0_r12_c8_rr0;
  wire [15:0] t0_r12_c8_rr1;
  wire [15:0] t0_r12_c8_rr2;
  wire [15:0] t0_r12_c8_rr3;
  wire [15:0] t0_r12_c8_rr4;
  wire [15:0] t0_r12_c8_rr5;
  wire [15:0] t0_r12_c8_rr6;
  wire [15:0] t0_r12_c8_rr7;
  wire [15:0] t0_r12_c8_rr8;
  wire [15:0] t0_r12_c8_rr9;
  wire [15:0] t0_r12_c8_rr10;
  wire [15:0] t0_r12_c8_rr11;
  wire [15:0] t0_r12_c8_rr12;
  wire [15:0] t0_r12_c8_rr13;
  wire [15:0] t0_r12_c8_rr14;
  wire [15:0] t1_r12_c8_rr0;
  wire [15:0] t1_r12_c8_rr1;
  wire [15:0] t1_r12_c8_rr2;
  wire [15:0] t1_r12_c8_rr3;
  wire [15:0] t1_r12_c8_rr4;
  wire [15:0] t1_r12_c8_rr5;
  wire [15:0] t1_r12_c8_rr6;
  wire [15:0] t1_r12_c8_rr7;
  wire [15:0] t2_r12_c8_rr0;
  wire [15:0] t2_r12_c8_rr1;
  wire [15:0] t2_r12_c8_rr2;
  wire [15:0] t2_r12_c8_rr3;
  wire [15:0] t3_r12_c8_rr0;
  wire [15:0] t3_r12_c8_rr1;
  wire [15:0] t4_r12_c8_rr0;
  wire [15:0] t0_r12_c9_rr0;
  wire [15:0] t0_r12_c9_rr1;
  wire [15:0] t0_r12_c9_rr2;
  wire [15:0] t0_r12_c9_rr3;
  wire [15:0] t0_r12_c9_rr4;
  wire [15:0] t0_r12_c9_rr5;
  wire [15:0] t0_r12_c9_rr6;
  wire [15:0] t0_r12_c9_rr7;
  wire [15:0] t0_r12_c9_rr8;
  wire [15:0] t0_r12_c9_rr9;
  wire [15:0] t0_r12_c9_rr10;
  wire [15:0] t0_r12_c9_rr11;
  wire [15:0] t0_r12_c9_rr12;
  wire [15:0] t0_r12_c9_rr13;
  wire [15:0] t0_r12_c9_rr14;
  wire [15:0] t1_r12_c9_rr0;
  wire [15:0] t1_r12_c9_rr1;
  wire [15:0] t1_r12_c9_rr2;
  wire [15:0] t1_r12_c9_rr3;
  wire [15:0] t1_r12_c9_rr4;
  wire [15:0] t1_r12_c9_rr5;
  wire [15:0] t1_r12_c9_rr6;
  wire [15:0] t1_r12_c9_rr7;
  wire [15:0] t2_r12_c9_rr0;
  wire [15:0] t2_r12_c9_rr1;
  wire [15:0] t2_r12_c9_rr2;
  wire [15:0] t2_r12_c9_rr3;
  wire [15:0] t3_r12_c9_rr0;
  wire [15:0] t3_r12_c9_rr1;
  wire [15:0] t4_r12_c9_rr0;
  wire [15:0] t0_r12_c10_rr0;
  wire [15:0] t0_r12_c10_rr1;
  wire [15:0] t0_r12_c10_rr2;
  wire [15:0] t0_r12_c10_rr3;
  wire [15:0] t0_r12_c10_rr4;
  wire [15:0] t0_r12_c10_rr5;
  wire [15:0] t0_r12_c10_rr6;
  wire [15:0] t0_r12_c10_rr7;
  wire [15:0] t0_r12_c10_rr8;
  wire [15:0] t0_r12_c10_rr9;
  wire [15:0] t0_r12_c10_rr10;
  wire [15:0] t0_r12_c10_rr11;
  wire [15:0] t0_r12_c10_rr12;
  wire [15:0] t0_r12_c10_rr13;
  wire [15:0] t0_r12_c10_rr14;
  wire [15:0] t1_r12_c10_rr0;
  wire [15:0] t1_r12_c10_rr1;
  wire [15:0] t1_r12_c10_rr2;
  wire [15:0] t1_r12_c10_rr3;
  wire [15:0] t1_r12_c10_rr4;
  wire [15:0] t1_r12_c10_rr5;
  wire [15:0] t1_r12_c10_rr6;
  wire [15:0] t1_r12_c10_rr7;
  wire [15:0] t2_r12_c10_rr0;
  wire [15:0] t2_r12_c10_rr1;
  wire [15:0] t2_r12_c10_rr2;
  wire [15:0] t2_r12_c10_rr3;
  wire [15:0] t3_r12_c10_rr0;
  wire [15:0] t3_r12_c10_rr1;
  wire [15:0] t4_r12_c10_rr0;
  wire [15:0] t0_r12_c11_rr0;
  wire [15:0] t0_r12_c11_rr1;
  wire [15:0] t0_r12_c11_rr2;
  wire [15:0] t0_r12_c11_rr3;
  wire [15:0] t0_r12_c11_rr4;
  wire [15:0] t0_r12_c11_rr5;
  wire [15:0] t0_r12_c11_rr6;
  wire [15:0] t0_r12_c11_rr7;
  wire [15:0] t0_r12_c11_rr8;
  wire [15:0] t0_r12_c11_rr9;
  wire [15:0] t0_r12_c11_rr10;
  wire [15:0] t0_r12_c11_rr11;
  wire [15:0] t0_r12_c11_rr12;
  wire [15:0] t0_r12_c11_rr13;
  wire [15:0] t0_r12_c11_rr14;
  wire [15:0] t1_r12_c11_rr0;
  wire [15:0] t1_r12_c11_rr1;
  wire [15:0] t1_r12_c11_rr2;
  wire [15:0] t1_r12_c11_rr3;
  wire [15:0] t1_r12_c11_rr4;
  wire [15:0] t1_r12_c11_rr5;
  wire [15:0] t1_r12_c11_rr6;
  wire [15:0] t1_r12_c11_rr7;
  wire [15:0] t2_r12_c11_rr0;
  wire [15:0] t2_r12_c11_rr1;
  wire [15:0] t2_r12_c11_rr2;
  wire [15:0] t2_r12_c11_rr3;
  wire [15:0] t3_r12_c11_rr0;
  wire [15:0] t3_r12_c11_rr1;
  wire [15:0] t4_r12_c11_rr0;
  wire [15:0] t0_r12_c12_rr0;
  wire [15:0] t0_r12_c12_rr1;
  wire [15:0] t0_r12_c12_rr2;
  wire [15:0] t0_r12_c12_rr3;
  wire [15:0] t0_r12_c12_rr4;
  wire [15:0] t0_r12_c12_rr5;
  wire [15:0] t0_r12_c12_rr6;
  wire [15:0] t0_r12_c12_rr7;
  wire [15:0] t0_r12_c12_rr8;
  wire [15:0] t0_r12_c12_rr9;
  wire [15:0] t0_r12_c12_rr10;
  wire [15:0] t0_r12_c12_rr11;
  wire [15:0] t0_r12_c12_rr12;
  wire [15:0] t0_r12_c12_rr13;
  wire [15:0] t0_r12_c12_rr14;
  wire [15:0] t1_r12_c12_rr0;
  wire [15:0] t1_r12_c12_rr1;
  wire [15:0] t1_r12_c12_rr2;
  wire [15:0] t1_r12_c12_rr3;
  wire [15:0] t1_r12_c12_rr4;
  wire [15:0] t1_r12_c12_rr5;
  wire [15:0] t1_r12_c12_rr6;
  wire [15:0] t1_r12_c12_rr7;
  wire [15:0] t2_r12_c12_rr0;
  wire [15:0] t2_r12_c12_rr1;
  wire [15:0] t2_r12_c12_rr2;
  wire [15:0] t2_r12_c12_rr3;
  wire [15:0] t3_r12_c12_rr0;
  wire [15:0] t3_r12_c12_rr1;
  wire [15:0] t4_r12_c12_rr0;
  wire [15:0] t0_r12_c13_rr0;
  wire [15:0] t0_r12_c13_rr1;
  wire [15:0] t0_r12_c13_rr2;
  wire [15:0] t0_r12_c13_rr3;
  wire [15:0] t0_r12_c13_rr4;
  wire [15:0] t0_r12_c13_rr5;
  wire [15:0] t0_r12_c13_rr6;
  wire [15:0] t0_r12_c13_rr7;
  wire [15:0] t0_r12_c13_rr8;
  wire [15:0] t0_r12_c13_rr9;
  wire [15:0] t0_r12_c13_rr10;
  wire [15:0] t0_r12_c13_rr11;
  wire [15:0] t0_r12_c13_rr12;
  wire [15:0] t0_r12_c13_rr13;
  wire [15:0] t0_r12_c13_rr14;
  wire [15:0] t1_r12_c13_rr0;
  wire [15:0] t1_r12_c13_rr1;
  wire [15:0] t1_r12_c13_rr2;
  wire [15:0] t1_r12_c13_rr3;
  wire [15:0] t1_r12_c13_rr4;
  wire [15:0] t1_r12_c13_rr5;
  wire [15:0] t1_r12_c13_rr6;
  wire [15:0] t1_r12_c13_rr7;
  wire [15:0] t2_r12_c13_rr0;
  wire [15:0] t2_r12_c13_rr1;
  wire [15:0] t2_r12_c13_rr2;
  wire [15:0] t2_r12_c13_rr3;
  wire [15:0] t3_r12_c13_rr0;
  wire [15:0] t3_r12_c13_rr1;
  wire [15:0] t4_r12_c13_rr0;
  wire [15:0] t0_r12_c14_rr0;
  wire [15:0] t0_r12_c14_rr1;
  wire [15:0] t0_r12_c14_rr2;
  wire [15:0] t0_r12_c14_rr3;
  wire [15:0] t0_r12_c14_rr4;
  wire [15:0] t0_r12_c14_rr5;
  wire [15:0] t0_r12_c14_rr6;
  wire [15:0] t0_r12_c14_rr7;
  wire [15:0] t0_r12_c14_rr8;
  wire [15:0] t0_r12_c14_rr9;
  wire [15:0] t0_r12_c14_rr10;
  wire [15:0] t0_r12_c14_rr11;
  wire [15:0] t0_r12_c14_rr12;
  wire [15:0] t0_r12_c14_rr13;
  wire [15:0] t0_r12_c14_rr14;
  wire [15:0] t1_r12_c14_rr0;
  wire [15:0] t1_r12_c14_rr1;
  wire [15:0] t1_r12_c14_rr2;
  wire [15:0] t1_r12_c14_rr3;
  wire [15:0] t1_r12_c14_rr4;
  wire [15:0] t1_r12_c14_rr5;
  wire [15:0] t1_r12_c14_rr6;
  wire [15:0] t1_r12_c14_rr7;
  wire [15:0] t2_r12_c14_rr0;
  wire [15:0] t2_r12_c14_rr1;
  wire [15:0] t2_r12_c14_rr2;
  wire [15:0] t2_r12_c14_rr3;
  wire [15:0] t3_r12_c14_rr0;
  wire [15:0] t3_r12_c14_rr1;
  wire [15:0] t4_r12_c14_rr0;
  wire [15:0] t0_r13_c0_rr0;
  wire [15:0] t0_r13_c0_rr1;
  wire [15:0] t0_r13_c0_rr2;
  wire [15:0] t0_r13_c0_rr3;
  wire [15:0] t0_r13_c0_rr4;
  wire [15:0] t0_r13_c0_rr5;
  wire [15:0] t0_r13_c0_rr6;
  wire [15:0] t0_r13_c0_rr7;
  wire [15:0] t0_r13_c0_rr8;
  wire [15:0] t0_r13_c0_rr9;
  wire [15:0] t0_r13_c0_rr10;
  wire [15:0] t0_r13_c0_rr11;
  wire [15:0] t0_r13_c0_rr12;
  wire [15:0] t0_r13_c0_rr13;
  wire [15:0] t0_r13_c0_rr14;
  wire [15:0] t1_r13_c0_rr0;
  wire [15:0] t1_r13_c0_rr1;
  wire [15:0] t1_r13_c0_rr2;
  wire [15:0] t1_r13_c0_rr3;
  wire [15:0] t1_r13_c0_rr4;
  wire [15:0] t1_r13_c0_rr5;
  wire [15:0] t1_r13_c0_rr6;
  wire [15:0] t1_r13_c0_rr7;
  wire [15:0] t2_r13_c0_rr0;
  wire [15:0] t2_r13_c0_rr1;
  wire [15:0] t2_r13_c0_rr2;
  wire [15:0] t2_r13_c0_rr3;
  wire [15:0] t3_r13_c0_rr0;
  wire [15:0] t3_r13_c0_rr1;
  wire [15:0] t4_r13_c0_rr0;
  wire [15:0] t0_r13_c1_rr0;
  wire [15:0] t0_r13_c1_rr1;
  wire [15:0] t0_r13_c1_rr2;
  wire [15:0] t0_r13_c1_rr3;
  wire [15:0] t0_r13_c1_rr4;
  wire [15:0] t0_r13_c1_rr5;
  wire [15:0] t0_r13_c1_rr6;
  wire [15:0] t0_r13_c1_rr7;
  wire [15:0] t0_r13_c1_rr8;
  wire [15:0] t0_r13_c1_rr9;
  wire [15:0] t0_r13_c1_rr10;
  wire [15:0] t0_r13_c1_rr11;
  wire [15:0] t0_r13_c1_rr12;
  wire [15:0] t0_r13_c1_rr13;
  wire [15:0] t0_r13_c1_rr14;
  wire [15:0] t1_r13_c1_rr0;
  wire [15:0] t1_r13_c1_rr1;
  wire [15:0] t1_r13_c1_rr2;
  wire [15:0] t1_r13_c1_rr3;
  wire [15:0] t1_r13_c1_rr4;
  wire [15:0] t1_r13_c1_rr5;
  wire [15:0] t1_r13_c1_rr6;
  wire [15:0] t1_r13_c1_rr7;
  wire [15:0] t2_r13_c1_rr0;
  wire [15:0] t2_r13_c1_rr1;
  wire [15:0] t2_r13_c1_rr2;
  wire [15:0] t2_r13_c1_rr3;
  wire [15:0] t3_r13_c1_rr0;
  wire [15:0] t3_r13_c1_rr1;
  wire [15:0] t4_r13_c1_rr0;
  wire [15:0] t0_r13_c2_rr0;
  wire [15:0] t0_r13_c2_rr1;
  wire [15:0] t0_r13_c2_rr2;
  wire [15:0] t0_r13_c2_rr3;
  wire [15:0] t0_r13_c2_rr4;
  wire [15:0] t0_r13_c2_rr5;
  wire [15:0] t0_r13_c2_rr6;
  wire [15:0] t0_r13_c2_rr7;
  wire [15:0] t0_r13_c2_rr8;
  wire [15:0] t0_r13_c2_rr9;
  wire [15:0] t0_r13_c2_rr10;
  wire [15:0] t0_r13_c2_rr11;
  wire [15:0] t0_r13_c2_rr12;
  wire [15:0] t0_r13_c2_rr13;
  wire [15:0] t0_r13_c2_rr14;
  wire [15:0] t1_r13_c2_rr0;
  wire [15:0] t1_r13_c2_rr1;
  wire [15:0] t1_r13_c2_rr2;
  wire [15:0] t1_r13_c2_rr3;
  wire [15:0] t1_r13_c2_rr4;
  wire [15:0] t1_r13_c2_rr5;
  wire [15:0] t1_r13_c2_rr6;
  wire [15:0] t1_r13_c2_rr7;
  wire [15:0] t2_r13_c2_rr0;
  wire [15:0] t2_r13_c2_rr1;
  wire [15:0] t2_r13_c2_rr2;
  wire [15:0] t2_r13_c2_rr3;
  wire [15:0] t3_r13_c2_rr0;
  wire [15:0] t3_r13_c2_rr1;
  wire [15:0] t4_r13_c2_rr0;
  wire [15:0] t0_r13_c3_rr0;
  wire [15:0] t0_r13_c3_rr1;
  wire [15:0] t0_r13_c3_rr2;
  wire [15:0] t0_r13_c3_rr3;
  wire [15:0] t0_r13_c3_rr4;
  wire [15:0] t0_r13_c3_rr5;
  wire [15:0] t0_r13_c3_rr6;
  wire [15:0] t0_r13_c3_rr7;
  wire [15:0] t0_r13_c3_rr8;
  wire [15:0] t0_r13_c3_rr9;
  wire [15:0] t0_r13_c3_rr10;
  wire [15:0] t0_r13_c3_rr11;
  wire [15:0] t0_r13_c3_rr12;
  wire [15:0] t0_r13_c3_rr13;
  wire [15:0] t0_r13_c3_rr14;
  wire [15:0] t1_r13_c3_rr0;
  wire [15:0] t1_r13_c3_rr1;
  wire [15:0] t1_r13_c3_rr2;
  wire [15:0] t1_r13_c3_rr3;
  wire [15:0] t1_r13_c3_rr4;
  wire [15:0] t1_r13_c3_rr5;
  wire [15:0] t1_r13_c3_rr6;
  wire [15:0] t1_r13_c3_rr7;
  wire [15:0] t2_r13_c3_rr0;
  wire [15:0] t2_r13_c3_rr1;
  wire [15:0] t2_r13_c3_rr2;
  wire [15:0] t2_r13_c3_rr3;
  wire [15:0] t3_r13_c3_rr0;
  wire [15:0] t3_r13_c3_rr1;
  wire [15:0] t4_r13_c3_rr0;
  wire [15:0] t0_r13_c4_rr0;
  wire [15:0] t0_r13_c4_rr1;
  wire [15:0] t0_r13_c4_rr2;
  wire [15:0] t0_r13_c4_rr3;
  wire [15:0] t0_r13_c4_rr4;
  wire [15:0] t0_r13_c4_rr5;
  wire [15:0] t0_r13_c4_rr6;
  wire [15:0] t0_r13_c4_rr7;
  wire [15:0] t0_r13_c4_rr8;
  wire [15:0] t0_r13_c4_rr9;
  wire [15:0] t0_r13_c4_rr10;
  wire [15:0] t0_r13_c4_rr11;
  wire [15:0] t0_r13_c4_rr12;
  wire [15:0] t0_r13_c4_rr13;
  wire [15:0] t0_r13_c4_rr14;
  wire [15:0] t1_r13_c4_rr0;
  wire [15:0] t1_r13_c4_rr1;
  wire [15:0] t1_r13_c4_rr2;
  wire [15:0] t1_r13_c4_rr3;
  wire [15:0] t1_r13_c4_rr4;
  wire [15:0] t1_r13_c4_rr5;
  wire [15:0] t1_r13_c4_rr6;
  wire [15:0] t1_r13_c4_rr7;
  wire [15:0] t2_r13_c4_rr0;
  wire [15:0] t2_r13_c4_rr1;
  wire [15:0] t2_r13_c4_rr2;
  wire [15:0] t2_r13_c4_rr3;
  wire [15:0] t3_r13_c4_rr0;
  wire [15:0] t3_r13_c4_rr1;
  wire [15:0] t4_r13_c4_rr0;
  wire [15:0] t0_r13_c5_rr0;
  wire [15:0] t0_r13_c5_rr1;
  wire [15:0] t0_r13_c5_rr2;
  wire [15:0] t0_r13_c5_rr3;
  wire [15:0] t0_r13_c5_rr4;
  wire [15:0] t0_r13_c5_rr5;
  wire [15:0] t0_r13_c5_rr6;
  wire [15:0] t0_r13_c5_rr7;
  wire [15:0] t0_r13_c5_rr8;
  wire [15:0] t0_r13_c5_rr9;
  wire [15:0] t0_r13_c5_rr10;
  wire [15:0] t0_r13_c5_rr11;
  wire [15:0] t0_r13_c5_rr12;
  wire [15:0] t0_r13_c5_rr13;
  wire [15:0] t0_r13_c5_rr14;
  wire [15:0] t1_r13_c5_rr0;
  wire [15:0] t1_r13_c5_rr1;
  wire [15:0] t1_r13_c5_rr2;
  wire [15:0] t1_r13_c5_rr3;
  wire [15:0] t1_r13_c5_rr4;
  wire [15:0] t1_r13_c5_rr5;
  wire [15:0] t1_r13_c5_rr6;
  wire [15:0] t1_r13_c5_rr7;
  wire [15:0] t2_r13_c5_rr0;
  wire [15:0] t2_r13_c5_rr1;
  wire [15:0] t2_r13_c5_rr2;
  wire [15:0] t2_r13_c5_rr3;
  wire [15:0] t3_r13_c5_rr0;
  wire [15:0] t3_r13_c5_rr1;
  wire [15:0] t4_r13_c5_rr0;
  wire [15:0] t0_r13_c6_rr0;
  wire [15:0] t0_r13_c6_rr1;
  wire [15:0] t0_r13_c6_rr2;
  wire [15:0] t0_r13_c6_rr3;
  wire [15:0] t0_r13_c6_rr4;
  wire [15:0] t0_r13_c6_rr5;
  wire [15:0] t0_r13_c6_rr6;
  wire [15:0] t0_r13_c6_rr7;
  wire [15:0] t0_r13_c6_rr8;
  wire [15:0] t0_r13_c6_rr9;
  wire [15:0] t0_r13_c6_rr10;
  wire [15:0] t0_r13_c6_rr11;
  wire [15:0] t0_r13_c6_rr12;
  wire [15:0] t0_r13_c6_rr13;
  wire [15:0] t0_r13_c6_rr14;
  wire [15:0] t1_r13_c6_rr0;
  wire [15:0] t1_r13_c6_rr1;
  wire [15:0] t1_r13_c6_rr2;
  wire [15:0] t1_r13_c6_rr3;
  wire [15:0] t1_r13_c6_rr4;
  wire [15:0] t1_r13_c6_rr5;
  wire [15:0] t1_r13_c6_rr6;
  wire [15:0] t1_r13_c6_rr7;
  wire [15:0] t2_r13_c6_rr0;
  wire [15:0] t2_r13_c6_rr1;
  wire [15:0] t2_r13_c6_rr2;
  wire [15:0] t2_r13_c6_rr3;
  wire [15:0] t3_r13_c6_rr0;
  wire [15:0] t3_r13_c6_rr1;
  wire [15:0] t4_r13_c6_rr0;
  wire [15:0] t0_r13_c7_rr0;
  wire [15:0] t0_r13_c7_rr1;
  wire [15:0] t0_r13_c7_rr2;
  wire [15:0] t0_r13_c7_rr3;
  wire [15:0] t0_r13_c7_rr4;
  wire [15:0] t0_r13_c7_rr5;
  wire [15:0] t0_r13_c7_rr6;
  wire [15:0] t0_r13_c7_rr7;
  wire [15:0] t0_r13_c7_rr8;
  wire [15:0] t0_r13_c7_rr9;
  wire [15:0] t0_r13_c7_rr10;
  wire [15:0] t0_r13_c7_rr11;
  wire [15:0] t0_r13_c7_rr12;
  wire [15:0] t0_r13_c7_rr13;
  wire [15:0] t0_r13_c7_rr14;
  wire [15:0] t1_r13_c7_rr0;
  wire [15:0] t1_r13_c7_rr1;
  wire [15:0] t1_r13_c7_rr2;
  wire [15:0] t1_r13_c7_rr3;
  wire [15:0] t1_r13_c7_rr4;
  wire [15:0] t1_r13_c7_rr5;
  wire [15:0] t1_r13_c7_rr6;
  wire [15:0] t1_r13_c7_rr7;
  wire [15:0] t2_r13_c7_rr0;
  wire [15:0] t2_r13_c7_rr1;
  wire [15:0] t2_r13_c7_rr2;
  wire [15:0] t2_r13_c7_rr3;
  wire [15:0] t3_r13_c7_rr0;
  wire [15:0] t3_r13_c7_rr1;
  wire [15:0] t4_r13_c7_rr0;
  wire [15:0] t0_r13_c8_rr0;
  wire [15:0] t0_r13_c8_rr1;
  wire [15:0] t0_r13_c8_rr2;
  wire [15:0] t0_r13_c8_rr3;
  wire [15:0] t0_r13_c8_rr4;
  wire [15:0] t0_r13_c8_rr5;
  wire [15:0] t0_r13_c8_rr6;
  wire [15:0] t0_r13_c8_rr7;
  wire [15:0] t0_r13_c8_rr8;
  wire [15:0] t0_r13_c8_rr9;
  wire [15:0] t0_r13_c8_rr10;
  wire [15:0] t0_r13_c8_rr11;
  wire [15:0] t0_r13_c8_rr12;
  wire [15:0] t0_r13_c8_rr13;
  wire [15:0] t0_r13_c8_rr14;
  wire [15:0] t1_r13_c8_rr0;
  wire [15:0] t1_r13_c8_rr1;
  wire [15:0] t1_r13_c8_rr2;
  wire [15:0] t1_r13_c8_rr3;
  wire [15:0] t1_r13_c8_rr4;
  wire [15:0] t1_r13_c8_rr5;
  wire [15:0] t1_r13_c8_rr6;
  wire [15:0] t1_r13_c8_rr7;
  wire [15:0] t2_r13_c8_rr0;
  wire [15:0] t2_r13_c8_rr1;
  wire [15:0] t2_r13_c8_rr2;
  wire [15:0] t2_r13_c8_rr3;
  wire [15:0] t3_r13_c8_rr0;
  wire [15:0] t3_r13_c8_rr1;
  wire [15:0] t4_r13_c8_rr0;
  wire [15:0] t0_r13_c9_rr0;
  wire [15:0] t0_r13_c9_rr1;
  wire [15:0] t0_r13_c9_rr2;
  wire [15:0] t0_r13_c9_rr3;
  wire [15:0] t0_r13_c9_rr4;
  wire [15:0] t0_r13_c9_rr5;
  wire [15:0] t0_r13_c9_rr6;
  wire [15:0] t0_r13_c9_rr7;
  wire [15:0] t0_r13_c9_rr8;
  wire [15:0] t0_r13_c9_rr9;
  wire [15:0] t0_r13_c9_rr10;
  wire [15:0] t0_r13_c9_rr11;
  wire [15:0] t0_r13_c9_rr12;
  wire [15:0] t0_r13_c9_rr13;
  wire [15:0] t0_r13_c9_rr14;
  wire [15:0] t1_r13_c9_rr0;
  wire [15:0] t1_r13_c9_rr1;
  wire [15:0] t1_r13_c9_rr2;
  wire [15:0] t1_r13_c9_rr3;
  wire [15:0] t1_r13_c9_rr4;
  wire [15:0] t1_r13_c9_rr5;
  wire [15:0] t1_r13_c9_rr6;
  wire [15:0] t1_r13_c9_rr7;
  wire [15:0] t2_r13_c9_rr0;
  wire [15:0] t2_r13_c9_rr1;
  wire [15:0] t2_r13_c9_rr2;
  wire [15:0] t2_r13_c9_rr3;
  wire [15:0] t3_r13_c9_rr0;
  wire [15:0] t3_r13_c9_rr1;
  wire [15:0] t4_r13_c9_rr0;
  wire [15:0] t0_r13_c10_rr0;
  wire [15:0] t0_r13_c10_rr1;
  wire [15:0] t0_r13_c10_rr2;
  wire [15:0] t0_r13_c10_rr3;
  wire [15:0] t0_r13_c10_rr4;
  wire [15:0] t0_r13_c10_rr5;
  wire [15:0] t0_r13_c10_rr6;
  wire [15:0] t0_r13_c10_rr7;
  wire [15:0] t0_r13_c10_rr8;
  wire [15:0] t0_r13_c10_rr9;
  wire [15:0] t0_r13_c10_rr10;
  wire [15:0] t0_r13_c10_rr11;
  wire [15:0] t0_r13_c10_rr12;
  wire [15:0] t0_r13_c10_rr13;
  wire [15:0] t0_r13_c10_rr14;
  wire [15:0] t1_r13_c10_rr0;
  wire [15:0] t1_r13_c10_rr1;
  wire [15:0] t1_r13_c10_rr2;
  wire [15:0] t1_r13_c10_rr3;
  wire [15:0] t1_r13_c10_rr4;
  wire [15:0] t1_r13_c10_rr5;
  wire [15:0] t1_r13_c10_rr6;
  wire [15:0] t1_r13_c10_rr7;
  wire [15:0] t2_r13_c10_rr0;
  wire [15:0] t2_r13_c10_rr1;
  wire [15:0] t2_r13_c10_rr2;
  wire [15:0] t2_r13_c10_rr3;
  wire [15:0] t3_r13_c10_rr0;
  wire [15:0] t3_r13_c10_rr1;
  wire [15:0] t4_r13_c10_rr0;
  wire [15:0] t0_r13_c11_rr0;
  wire [15:0] t0_r13_c11_rr1;
  wire [15:0] t0_r13_c11_rr2;
  wire [15:0] t0_r13_c11_rr3;
  wire [15:0] t0_r13_c11_rr4;
  wire [15:0] t0_r13_c11_rr5;
  wire [15:0] t0_r13_c11_rr6;
  wire [15:0] t0_r13_c11_rr7;
  wire [15:0] t0_r13_c11_rr8;
  wire [15:0] t0_r13_c11_rr9;
  wire [15:0] t0_r13_c11_rr10;
  wire [15:0] t0_r13_c11_rr11;
  wire [15:0] t0_r13_c11_rr12;
  wire [15:0] t0_r13_c11_rr13;
  wire [15:0] t0_r13_c11_rr14;
  wire [15:0] t1_r13_c11_rr0;
  wire [15:0] t1_r13_c11_rr1;
  wire [15:0] t1_r13_c11_rr2;
  wire [15:0] t1_r13_c11_rr3;
  wire [15:0] t1_r13_c11_rr4;
  wire [15:0] t1_r13_c11_rr5;
  wire [15:0] t1_r13_c11_rr6;
  wire [15:0] t1_r13_c11_rr7;
  wire [15:0] t2_r13_c11_rr0;
  wire [15:0] t2_r13_c11_rr1;
  wire [15:0] t2_r13_c11_rr2;
  wire [15:0] t2_r13_c11_rr3;
  wire [15:0] t3_r13_c11_rr0;
  wire [15:0] t3_r13_c11_rr1;
  wire [15:0] t4_r13_c11_rr0;
  wire [15:0] t0_r13_c12_rr0;
  wire [15:0] t0_r13_c12_rr1;
  wire [15:0] t0_r13_c12_rr2;
  wire [15:0] t0_r13_c12_rr3;
  wire [15:0] t0_r13_c12_rr4;
  wire [15:0] t0_r13_c12_rr5;
  wire [15:0] t0_r13_c12_rr6;
  wire [15:0] t0_r13_c12_rr7;
  wire [15:0] t0_r13_c12_rr8;
  wire [15:0] t0_r13_c12_rr9;
  wire [15:0] t0_r13_c12_rr10;
  wire [15:0] t0_r13_c12_rr11;
  wire [15:0] t0_r13_c12_rr12;
  wire [15:0] t0_r13_c12_rr13;
  wire [15:0] t0_r13_c12_rr14;
  wire [15:0] t1_r13_c12_rr0;
  wire [15:0] t1_r13_c12_rr1;
  wire [15:0] t1_r13_c12_rr2;
  wire [15:0] t1_r13_c12_rr3;
  wire [15:0] t1_r13_c12_rr4;
  wire [15:0] t1_r13_c12_rr5;
  wire [15:0] t1_r13_c12_rr6;
  wire [15:0] t1_r13_c12_rr7;
  wire [15:0] t2_r13_c12_rr0;
  wire [15:0] t2_r13_c12_rr1;
  wire [15:0] t2_r13_c12_rr2;
  wire [15:0] t2_r13_c12_rr3;
  wire [15:0] t3_r13_c12_rr0;
  wire [15:0] t3_r13_c12_rr1;
  wire [15:0] t4_r13_c12_rr0;
  wire [15:0] t0_r13_c13_rr0;
  wire [15:0] t0_r13_c13_rr1;
  wire [15:0] t0_r13_c13_rr2;
  wire [15:0] t0_r13_c13_rr3;
  wire [15:0] t0_r13_c13_rr4;
  wire [15:0] t0_r13_c13_rr5;
  wire [15:0] t0_r13_c13_rr6;
  wire [15:0] t0_r13_c13_rr7;
  wire [15:0] t0_r13_c13_rr8;
  wire [15:0] t0_r13_c13_rr9;
  wire [15:0] t0_r13_c13_rr10;
  wire [15:0] t0_r13_c13_rr11;
  wire [15:0] t0_r13_c13_rr12;
  wire [15:0] t0_r13_c13_rr13;
  wire [15:0] t0_r13_c13_rr14;
  wire [15:0] t1_r13_c13_rr0;
  wire [15:0] t1_r13_c13_rr1;
  wire [15:0] t1_r13_c13_rr2;
  wire [15:0] t1_r13_c13_rr3;
  wire [15:0] t1_r13_c13_rr4;
  wire [15:0] t1_r13_c13_rr5;
  wire [15:0] t1_r13_c13_rr6;
  wire [15:0] t1_r13_c13_rr7;
  wire [15:0] t2_r13_c13_rr0;
  wire [15:0] t2_r13_c13_rr1;
  wire [15:0] t2_r13_c13_rr2;
  wire [15:0] t2_r13_c13_rr3;
  wire [15:0] t3_r13_c13_rr0;
  wire [15:0] t3_r13_c13_rr1;
  wire [15:0] t4_r13_c13_rr0;
  wire [15:0] t0_r13_c14_rr0;
  wire [15:0] t0_r13_c14_rr1;
  wire [15:0] t0_r13_c14_rr2;
  wire [15:0] t0_r13_c14_rr3;
  wire [15:0] t0_r13_c14_rr4;
  wire [15:0] t0_r13_c14_rr5;
  wire [15:0] t0_r13_c14_rr6;
  wire [15:0] t0_r13_c14_rr7;
  wire [15:0] t0_r13_c14_rr8;
  wire [15:0] t0_r13_c14_rr9;
  wire [15:0] t0_r13_c14_rr10;
  wire [15:0] t0_r13_c14_rr11;
  wire [15:0] t0_r13_c14_rr12;
  wire [15:0] t0_r13_c14_rr13;
  wire [15:0] t0_r13_c14_rr14;
  wire [15:0] t1_r13_c14_rr0;
  wire [15:0] t1_r13_c14_rr1;
  wire [15:0] t1_r13_c14_rr2;
  wire [15:0] t1_r13_c14_rr3;
  wire [15:0] t1_r13_c14_rr4;
  wire [15:0] t1_r13_c14_rr5;
  wire [15:0] t1_r13_c14_rr6;
  wire [15:0] t1_r13_c14_rr7;
  wire [15:0] t2_r13_c14_rr0;
  wire [15:0] t2_r13_c14_rr1;
  wire [15:0] t2_r13_c14_rr2;
  wire [15:0] t2_r13_c14_rr3;
  wire [15:0] t3_r13_c14_rr0;
  wire [15:0] t3_r13_c14_rr1;
  wire [15:0] t4_r13_c14_rr0;
  wire [15:0] t0_r14_c0_rr0;
  wire [15:0] t0_r14_c0_rr1;
  wire [15:0] t0_r14_c0_rr2;
  wire [15:0] t0_r14_c0_rr3;
  wire [15:0] t0_r14_c0_rr4;
  wire [15:0] t0_r14_c0_rr5;
  wire [15:0] t0_r14_c0_rr6;
  wire [15:0] t0_r14_c0_rr7;
  wire [15:0] t0_r14_c0_rr8;
  wire [15:0] t0_r14_c0_rr9;
  wire [15:0] t0_r14_c0_rr10;
  wire [15:0] t0_r14_c0_rr11;
  wire [15:0] t0_r14_c0_rr12;
  wire [15:0] t0_r14_c0_rr13;
  wire [15:0] t0_r14_c0_rr14;
  wire [15:0] t1_r14_c0_rr0;
  wire [15:0] t1_r14_c0_rr1;
  wire [15:0] t1_r14_c0_rr2;
  wire [15:0] t1_r14_c0_rr3;
  wire [15:0] t1_r14_c0_rr4;
  wire [15:0] t1_r14_c0_rr5;
  wire [15:0] t1_r14_c0_rr6;
  wire [15:0] t1_r14_c0_rr7;
  wire [15:0] t2_r14_c0_rr0;
  wire [15:0] t2_r14_c0_rr1;
  wire [15:0] t2_r14_c0_rr2;
  wire [15:0] t2_r14_c0_rr3;
  wire [15:0] t3_r14_c0_rr0;
  wire [15:0] t3_r14_c0_rr1;
  wire [15:0] t4_r14_c0_rr0;
  wire [15:0] t0_r14_c1_rr0;
  wire [15:0] t0_r14_c1_rr1;
  wire [15:0] t0_r14_c1_rr2;
  wire [15:0] t0_r14_c1_rr3;
  wire [15:0] t0_r14_c1_rr4;
  wire [15:0] t0_r14_c1_rr5;
  wire [15:0] t0_r14_c1_rr6;
  wire [15:0] t0_r14_c1_rr7;
  wire [15:0] t0_r14_c1_rr8;
  wire [15:0] t0_r14_c1_rr9;
  wire [15:0] t0_r14_c1_rr10;
  wire [15:0] t0_r14_c1_rr11;
  wire [15:0] t0_r14_c1_rr12;
  wire [15:0] t0_r14_c1_rr13;
  wire [15:0] t0_r14_c1_rr14;
  wire [15:0] t1_r14_c1_rr0;
  wire [15:0] t1_r14_c1_rr1;
  wire [15:0] t1_r14_c1_rr2;
  wire [15:0] t1_r14_c1_rr3;
  wire [15:0] t1_r14_c1_rr4;
  wire [15:0] t1_r14_c1_rr5;
  wire [15:0] t1_r14_c1_rr6;
  wire [15:0] t1_r14_c1_rr7;
  wire [15:0] t2_r14_c1_rr0;
  wire [15:0] t2_r14_c1_rr1;
  wire [15:0] t2_r14_c1_rr2;
  wire [15:0] t2_r14_c1_rr3;
  wire [15:0] t3_r14_c1_rr0;
  wire [15:0] t3_r14_c1_rr1;
  wire [15:0] t4_r14_c1_rr0;
  wire [15:0] t0_r14_c2_rr0;
  wire [15:0] t0_r14_c2_rr1;
  wire [15:0] t0_r14_c2_rr2;
  wire [15:0] t0_r14_c2_rr3;
  wire [15:0] t0_r14_c2_rr4;
  wire [15:0] t0_r14_c2_rr5;
  wire [15:0] t0_r14_c2_rr6;
  wire [15:0] t0_r14_c2_rr7;
  wire [15:0] t0_r14_c2_rr8;
  wire [15:0] t0_r14_c2_rr9;
  wire [15:0] t0_r14_c2_rr10;
  wire [15:0] t0_r14_c2_rr11;
  wire [15:0] t0_r14_c2_rr12;
  wire [15:0] t0_r14_c2_rr13;
  wire [15:0] t0_r14_c2_rr14;
  wire [15:0] t1_r14_c2_rr0;
  wire [15:0] t1_r14_c2_rr1;
  wire [15:0] t1_r14_c2_rr2;
  wire [15:0] t1_r14_c2_rr3;
  wire [15:0] t1_r14_c2_rr4;
  wire [15:0] t1_r14_c2_rr5;
  wire [15:0] t1_r14_c2_rr6;
  wire [15:0] t1_r14_c2_rr7;
  wire [15:0] t2_r14_c2_rr0;
  wire [15:0] t2_r14_c2_rr1;
  wire [15:0] t2_r14_c2_rr2;
  wire [15:0] t2_r14_c2_rr3;
  wire [15:0] t3_r14_c2_rr0;
  wire [15:0] t3_r14_c2_rr1;
  wire [15:0] t4_r14_c2_rr0;
  wire [15:0] t0_r14_c3_rr0;
  wire [15:0] t0_r14_c3_rr1;
  wire [15:0] t0_r14_c3_rr2;
  wire [15:0] t0_r14_c3_rr3;
  wire [15:0] t0_r14_c3_rr4;
  wire [15:0] t0_r14_c3_rr5;
  wire [15:0] t0_r14_c3_rr6;
  wire [15:0] t0_r14_c3_rr7;
  wire [15:0] t0_r14_c3_rr8;
  wire [15:0] t0_r14_c3_rr9;
  wire [15:0] t0_r14_c3_rr10;
  wire [15:0] t0_r14_c3_rr11;
  wire [15:0] t0_r14_c3_rr12;
  wire [15:0] t0_r14_c3_rr13;
  wire [15:0] t0_r14_c3_rr14;
  wire [15:0] t1_r14_c3_rr0;
  wire [15:0] t1_r14_c3_rr1;
  wire [15:0] t1_r14_c3_rr2;
  wire [15:0] t1_r14_c3_rr3;
  wire [15:0] t1_r14_c3_rr4;
  wire [15:0] t1_r14_c3_rr5;
  wire [15:0] t1_r14_c3_rr6;
  wire [15:0] t1_r14_c3_rr7;
  wire [15:0] t2_r14_c3_rr0;
  wire [15:0] t2_r14_c3_rr1;
  wire [15:0] t2_r14_c3_rr2;
  wire [15:0] t2_r14_c3_rr3;
  wire [15:0] t3_r14_c3_rr0;
  wire [15:0] t3_r14_c3_rr1;
  wire [15:0] t4_r14_c3_rr0;
  wire [15:0] t0_r14_c4_rr0;
  wire [15:0] t0_r14_c4_rr1;
  wire [15:0] t0_r14_c4_rr2;
  wire [15:0] t0_r14_c4_rr3;
  wire [15:0] t0_r14_c4_rr4;
  wire [15:0] t0_r14_c4_rr5;
  wire [15:0] t0_r14_c4_rr6;
  wire [15:0] t0_r14_c4_rr7;
  wire [15:0] t0_r14_c4_rr8;
  wire [15:0] t0_r14_c4_rr9;
  wire [15:0] t0_r14_c4_rr10;
  wire [15:0] t0_r14_c4_rr11;
  wire [15:0] t0_r14_c4_rr12;
  wire [15:0] t0_r14_c4_rr13;
  wire [15:0] t0_r14_c4_rr14;
  wire [15:0] t1_r14_c4_rr0;
  wire [15:0] t1_r14_c4_rr1;
  wire [15:0] t1_r14_c4_rr2;
  wire [15:0] t1_r14_c4_rr3;
  wire [15:0] t1_r14_c4_rr4;
  wire [15:0] t1_r14_c4_rr5;
  wire [15:0] t1_r14_c4_rr6;
  wire [15:0] t1_r14_c4_rr7;
  wire [15:0] t2_r14_c4_rr0;
  wire [15:0] t2_r14_c4_rr1;
  wire [15:0] t2_r14_c4_rr2;
  wire [15:0] t2_r14_c4_rr3;
  wire [15:0] t3_r14_c4_rr0;
  wire [15:0] t3_r14_c4_rr1;
  wire [15:0] t4_r14_c4_rr0;
  wire [15:0] t0_r14_c5_rr0;
  wire [15:0] t0_r14_c5_rr1;
  wire [15:0] t0_r14_c5_rr2;
  wire [15:0] t0_r14_c5_rr3;
  wire [15:0] t0_r14_c5_rr4;
  wire [15:0] t0_r14_c5_rr5;
  wire [15:0] t0_r14_c5_rr6;
  wire [15:0] t0_r14_c5_rr7;
  wire [15:0] t0_r14_c5_rr8;
  wire [15:0] t0_r14_c5_rr9;
  wire [15:0] t0_r14_c5_rr10;
  wire [15:0] t0_r14_c5_rr11;
  wire [15:0] t0_r14_c5_rr12;
  wire [15:0] t0_r14_c5_rr13;
  wire [15:0] t0_r14_c5_rr14;
  wire [15:0] t1_r14_c5_rr0;
  wire [15:0] t1_r14_c5_rr1;
  wire [15:0] t1_r14_c5_rr2;
  wire [15:0] t1_r14_c5_rr3;
  wire [15:0] t1_r14_c5_rr4;
  wire [15:0] t1_r14_c5_rr5;
  wire [15:0] t1_r14_c5_rr6;
  wire [15:0] t1_r14_c5_rr7;
  wire [15:0] t2_r14_c5_rr0;
  wire [15:0] t2_r14_c5_rr1;
  wire [15:0] t2_r14_c5_rr2;
  wire [15:0] t2_r14_c5_rr3;
  wire [15:0] t3_r14_c5_rr0;
  wire [15:0] t3_r14_c5_rr1;
  wire [15:0] t4_r14_c5_rr0;
  wire [15:0] t0_r14_c6_rr0;
  wire [15:0] t0_r14_c6_rr1;
  wire [15:0] t0_r14_c6_rr2;
  wire [15:0] t0_r14_c6_rr3;
  wire [15:0] t0_r14_c6_rr4;
  wire [15:0] t0_r14_c6_rr5;
  wire [15:0] t0_r14_c6_rr6;
  wire [15:0] t0_r14_c6_rr7;
  wire [15:0] t0_r14_c6_rr8;
  wire [15:0] t0_r14_c6_rr9;
  wire [15:0] t0_r14_c6_rr10;
  wire [15:0] t0_r14_c6_rr11;
  wire [15:0] t0_r14_c6_rr12;
  wire [15:0] t0_r14_c6_rr13;
  wire [15:0] t0_r14_c6_rr14;
  wire [15:0] t1_r14_c6_rr0;
  wire [15:0] t1_r14_c6_rr1;
  wire [15:0] t1_r14_c6_rr2;
  wire [15:0] t1_r14_c6_rr3;
  wire [15:0] t1_r14_c6_rr4;
  wire [15:0] t1_r14_c6_rr5;
  wire [15:0] t1_r14_c6_rr6;
  wire [15:0] t1_r14_c6_rr7;
  wire [15:0] t2_r14_c6_rr0;
  wire [15:0] t2_r14_c6_rr1;
  wire [15:0] t2_r14_c6_rr2;
  wire [15:0] t2_r14_c6_rr3;
  wire [15:0] t3_r14_c6_rr0;
  wire [15:0] t3_r14_c6_rr1;
  wire [15:0] t4_r14_c6_rr0;
  wire [15:0] t0_r14_c7_rr0;
  wire [15:0] t0_r14_c7_rr1;
  wire [15:0] t0_r14_c7_rr2;
  wire [15:0] t0_r14_c7_rr3;
  wire [15:0] t0_r14_c7_rr4;
  wire [15:0] t0_r14_c7_rr5;
  wire [15:0] t0_r14_c7_rr6;
  wire [15:0] t0_r14_c7_rr7;
  wire [15:0] t0_r14_c7_rr8;
  wire [15:0] t0_r14_c7_rr9;
  wire [15:0] t0_r14_c7_rr10;
  wire [15:0] t0_r14_c7_rr11;
  wire [15:0] t0_r14_c7_rr12;
  wire [15:0] t0_r14_c7_rr13;
  wire [15:0] t0_r14_c7_rr14;
  wire [15:0] t1_r14_c7_rr0;
  wire [15:0] t1_r14_c7_rr1;
  wire [15:0] t1_r14_c7_rr2;
  wire [15:0] t1_r14_c7_rr3;
  wire [15:0] t1_r14_c7_rr4;
  wire [15:0] t1_r14_c7_rr5;
  wire [15:0] t1_r14_c7_rr6;
  wire [15:0] t1_r14_c7_rr7;
  wire [15:0] t2_r14_c7_rr0;
  wire [15:0] t2_r14_c7_rr1;
  wire [15:0] t2_r14_c7_rr2;
  wire [15:0] t2_r14_c7_rr3;
  wire [15:0] t3_r14_c7_rr0;
  wire [15:0] t3_r14_c7_rr1;
  wire [15:0] t4_r14_c7_rr0;
  wire [15:0] t0_r14_c8_rr0;
  wire [15:0] t0_r14_c8_rr1;
  wire [15:0] t0_r14_c8_rr2;
  wire [15:0] t0_r14_c8_rr3;
  wire [15:0] t0_r14_c8_rr4;
  wire [15:0] t0_r14_c8_rr5;
  wire [15:0] t0_r14_c8_rr6;
  wire [15:0] t0_r14_c8_rr7;
  wire [15:0] t0_r14_c8_rr8;
  wire [15:0] t0_r14_c8_rr9;
  wire [15:0] t0_r14_c8_rr10;
  wire [15:0] t0_r14_c8_rr11;
  wire [15:0] t0_r14_c8_rr12;
  wire [15:0] t0_r14_c8_rr13;
  wire [15:0] t0_r14_c8_rr14;
  wire [15:0] t1_r14_c8_rr0;
  wire [15:0] t1_r14_c8_rr1;
  wire [15:0] t1_r14_c8_rr2;
  wire [15:0] t1_r14_c8_rr3;
  wire [15:0] t1_r14_c8_rr4;
  wire [15:0] t1_r14_c8_rr5;
  wire [15:0] t1_r14_c8_rr6;
  wire [15:0] t1_r14_c8_rr7;
  wire [15:0] t2_r14_c8_rr0;
  wire [15:0] t2_r14_c8_rr1;
  wire [15:0] t2_r14_c8_rr2;
  wire [15:0] t2_r14_c8_rr3;
  wire [15:0] t3_r14_c8_rr0;
  wire [15:0] t3_r14_c8_rr1;
  wire [15:0] t4_r14_c8_rr0;
  wire [15:0] t0_r14_c9_rr0;
  wire [15:0] t0_r14_c9_rr1;
  wire [15:0] t0_r14_c9_rr2;
  wire [15:0] t0_r14_c9_rr3;
  wire [15:0] t0_r14_c9_rr4;
  wire [15:0] t0_r14_c9_rr5;
  wire [15:0] t0_r14_c9_rr6;
  wire [15:0] t0_r14_c9_rr7;
  wire [15:0] t0_r14_c9_rr8;
  wire [15:0] t0_r14_c9_rr9;
  wire [15:0] t0_r14_c9_rr10;
  wire [15:0] t0_r14_c9_rr11;
  wire [15:0] t0_r14_c9_rr12;
  wire [15:0] t0_r14_c9_rr13;
  wire [15:0] t0_r14_c9_rr14;
  wire [15:0] t1_r14_c9_rr0;
  wire [15:0] t1_r14_c9_rr1;
  wire [15:0] t1_r14_c9_rr2;
  wire [15:0] t1_r14_c9_rr3;
  wire [15:0] t1_r14_c9_rr4;
  wire [15:0] t1_r14_c9_rr5;
  wire [15:0] t1_r14_c9_rr6;
  wire [15:0] t1_r14_c9_rr7;
  wire [15:0] t2_r14_c9_rr0;
  wire [15:0] t2_r14_c9_rr1;
  wire [15:0] t2_r14_c9_rr2;
  wire [15:0] t2_r14_c9_rr3;
  wire [15:0] t3_r14_c9_rr0;
  wire [15:0] t3_r14_c9_rr1;
  wire [15:0] t4_r14_c9_rr0;
  wire [15:0] t0_r14_c10_rr0;
  wire [15:0] t0_r14_c10_rr1;
  wire [15:0] t0_r14_c10_rr2;
  wire [15:0] t0_r14_c10_rr3;
  wire [15:0] t0_r14_c10_rr4;
  wire [15:0] t0_r14_c10_rr5;
  wire [15:0] t0_r14_c10_rr6;
  wire [15:0] t0_r14_c10_rr7;
  wire [15:0] t0_r14_c10_rr8;
  wire [15:0] t0_r14_c10_rr9;
  wire [15:0] t0_r14_c10_rr10;
  wire [15:0] t0_r14_c10_rr11;
  wire [15:0] t0_r14_c10_rr12;
  wire [15:0] t0_r14_c10_rr13;
  wire [15:0] t0_r14_c10_rr14;
  wire [15:0] t1_r14_c10_rr0;
  wire [15:0] t1_r14_c10_rr1;
  wire [15:0] t1_r14_c10_rr2;
  wire [15:0] t1_r14_c10_rr3;
  wire [15:0] t1_r14_c10_rr4;
  wire [15:0] t1_r14_c10_rr5;
  wire [15:0] t1_r14_c10_rr6;
  wire [15:0] t1_r14_c10_rr7;
  wire [15:0] t2_r14_c10_rr0;
  wire [15:0] t2_r14_c10_rr1;
  wire [15:0] t2_r14_c10_rr2;
  wire [15:0] t2_r14_c10_rr3;
  wire [15:0] t3_r14_c10_rr0;
  wire [15:0] t3_r14_c10_rr1;
  wire [15:0] t4_r14_c10_rr0;
  wire [15:0] t0_r14_c11_rr0;
  wire [15:0] t0_r14_c11_rr1;
  wire [15:0] t0_r14_c11_rr2;
  wire [15:0] t0_r14_c11_rr3;
  wire [15:0] t0_r14_c11_rr4;
  wire [15:0] t0_r14_c11_rr5;
  wire [15:0] t0_r14_c11_rr6;
  wire [15:0] t0_r14_c11_rr7;
  wire [15:0] t0_r14_c11_rr8;
  wire [15:0] t0_r14_c11_rr9;
  wire [15:0] t0_r14_c11_rr10;
  wire [15:0] t0_r14_c11_rr11;
  wire [15:0] t0_r14_c11_rr12;
  wire [15:0] t0_r14_c11_rr13;
  wire [15:0] t0_r14_c11_rr14;
  wire [15:0] t1_r14_c11_rr0;
  wire [15:0] t1_r14_c11_rr1;
  wire [15:0] t1_r14_c11_rr2;
  wire [15:0] t1_r14_c11_rr3;
  wire [15:0] t1_r14_c11_rr4;
  wire [15:0] t1_r14_c11_rr5;
  wire [15:0] t1_r14_c11_rr6;
  wire [15:0] t1_r14_c11_rr7;
  wire [15:0] t2_r14_c11_rr0;
  wire [15:0] t2_r14_c11_rr1;
  wire [15:0] t2_r14_c11_rr2;
  wire [15:0] t2_r14_c11_rr3;
  wire [15:0] t3_r14_c11_rr0;
  wire [15:0] t3_r14_c11_rr1;
  wire [15:0] t4_r14_c11_rr0;
  wire [15:0] t0_r14_c12_rr0;
  wire [15:0] t0_r14_c12_rr1;
  wire [15:0] t0_r14_c12_rr2;
  wire [15:0] t0_r14_c12_rr3;
  wire [15:0] t0_r14_c12_rr4;
  wire [15:0] t0_r14_c12_rr5;
  wire [15:0] t0_r14_c12_rr6;
  wire [15:0] t0_r14_c12_rr7;
  wire [15:0] t0_r14_c12_rr8;
  wire [15:0] t0_r14_c12_rr9;
  wire [15:0] t0_r14_c12_rr10;
  wire [15:0] t0_r14_c12_rr11;
  wire [15:0] t0_r14_c12_rr12;
  wire [15:0] t0_r14_c12_rr13;
  wire [15:0] t0_r14_c12_rr14;
  wire [15:0] t1_r14_c12_rr0;
  wire [15:0] t1_r14_c12_rr1;
  wire [15:0] t1_r14_c12_rr2;
  wire [15:0] t1_r14_c12_rr3;
  wire [15:0] t1_r14_c12_rr4;
  wire [15:0] t1_r14_c12_rr5;
  wire [15:0] t1_r14_c12_rr6;
  wire [15:0] t1_r14_c12_rr7;
  wire [15:0] t2_r14_c12_rr0;
  wire [15:0] t2_r14_c12_rr1;
  wire [15:0] t2_r14_c12_rr2;
  wire [15:0] t2_r14_c12_rr3;
  wire [15:0] t3_r14_c12_rr0;
  wire [15:0] t3_r14_c12_rr1;
  wire [15:0] t4_r14_c12_rr0;
  wire [15:0] t0_r14_c13_rr0;
  wire [15:0] t0_r14_c13_rr1;
  wire [15:0] t0_r14_c13_rr2;
  wire [15:0] t0_r14_c13_rr3;
  wire [15:0] t0_r14_c13_rr4;
  wire [15:0] t0_r14_c13_rr5;
  wire [15:0] t0_r14_c13_rr6;
  wire [15:0] t0_r14_c13_rr7;
  wire [15:0] t0_r14_c13_rr8;
  wire [15:0] t0_r14_c13_rr9;
  wire [15:0] t0_r14_c13_rr10;
  wire [15:0] t0_r14_c13_rr11;
  wire [15:0] t0_r14_c13_rr12;
  wire [15:0] t0_r14_c13_rr13;
  wire [15:0] t0_r14_c13_rr14;
  wire [15:0] t1_r14_c13_rr0;
  wire [15:0] t1_r14_c13_rr1;
  wire [15:0] t1_r14_c13_rr2;
  wire [15:0] t1_r14_c13_rr3;
  wire [15:0] t1_r14_c13_rr4;
  wire [15:0] t1_r14_c13_rr5;
  wire [15:0] t1_r14_c13_rr6;
  wire [15:0] t1_r14_c13_rr7;
  wire [15:0] t2_r14_c13_rr0;
  wire [15:0] t2_r14_c13_rr1;
  wire [15:0] t2_r14_c13_rr2;
  wire [15:0] t2_r14_c13_rr3;
  wire [15:0] t3_r14_c13_rr0;
  wire [15:0] t3_r14_c13_rr1;
  wire [15:0] t4_r14_c13_rr0;
  wire [15:0] t0_r14_c14_rr0;
  wire [15:0] t0_r14_c14_rr1;
  wire [15:0] t0_r14_c14_rr2;
  wire [15:0] t0_r14_c14_rr3;
  wire [15:0] t0_r14_c14_rr4;
  wire [15:0] t0_r14_c14_rr5;
  wire [15:0] t0_r14_c14_rr6;
  wire [15:0] t0_r14_c14_rr7;
  wire [15:0] t0_r14_c14_rr8;
  wire [15:0] t0_r14_c14_rr9;
  wire [15:0] t0_r14_c14_rr10;
  wire [15:0] t0_r14_c14_rr11;
  wire [15:0] t0_r14_c14_rr12;
  wire [15:0] t0_r14_c14_rr13;
  wire [15:0] t0_r14_c14_rr14;
  wire [15:0] t1_r14_c14_rr0;
  wire [15:0] t1_r14_c14_rr1;
  wire [15:0] t1_r14_c14_rr2;
  wire [15:0] t1_r14_c14_rr3;
  wire [15:0] t1_r14_c14_rr4;
  wire [15:0] t1_r14_c14_rr5;
  wire [15:0] t1_r14_c14_rr6;
  wire [15:0] t1_r14_c14_rr7;
  wire [15:0] t2_r14_c14_rr0;
  wire [15:0] t2_r14_c14_rr1;
  wire [15:0] t2_r14_c14_rr2;
  wire [15:0] t2_r14_c14_rr3;
  wire [15:0] t3_r14_c14_rr0;
  wire [15:0] t3_r14_c14_rr1;
  wire [15:0] t4_r14_c14_rr0;

  assign t0_r0_c0_rr0 = a_0_0 * b_0_0;
  assign t0_r0_c0_rr1 = a_0_1 * b_1_0;
  assign t0_r0_c0_rr2 = a_0_2 * b_2_0;
  assign t0_r0_c0_rr3 = a_0_3 * b_3_0;
  assign t0_r0_c0_rr4 = a_0_4 * b_4_0;
  assign t0_r0_c0_rr5 = a_0_5 * b_5_0;
  assign t0_r0_c0_rr6 = a_0_6 * b_6_0;
  assign t0_r0_c0_rr7 = a_0_7 * b_7_0;
  assign t0_r0_c0_rr8 = a_0_8 * b_8_0;
  assign t0_r0_c0_rr9 = a_0_9 * b_9_0;
  assign t0_r0_c0_rr10 = a_0_10 * b_10_0;
  assign t0_r0_c0_rr11 = a_0_11 * b_11_0;
  assign t0_r0_c0_rr12 = a_0_12 * b_12_0;
  assign t0_r0_c0_rr13 = a_0_13 * b_13_0;
  assign t0_r0_c0_rr14 = a_0_14 * b_14_0;
  assign t1_r0_c0_rr0 = t0_r0_c0_rr0 + t0_r0_c0_rr1;
  assign t1_r0_c0_rr1 = t0_r0_c0_rr2 + t0_r0_c0_rr3;
  assign t1_r0_c0_rr2 = t0_r0_c0_rr4 + t0_r0_c0_rr5;
  assign t1_r0_c0_rr3 = t0_r0_c0_rr6 + t0_r0_c0_rr7;
  assign t1_r0_c0_rr4 = t0_r0_c0_rr8 + t0_r0_c0_rr9;
  assign t1_r0_c0_rr5 = t0_r0_c0_rr10 + t0_r0_c0_rr11;
  assign t1_r0_c0_rr6 = t0_r0_c0_rr12 + t0_r0_c0_rr13;
  assign t1_r0_c0_rr7 = t0_r0_c0_rr14;

  assign t2_r0_c0_rr0 = t1_r0_c0_rr0 + t1_r0_c0_rr1;
  assign t2_r0_c0_rr1 = t1_r0_c0_rr2 + t1_r0_c0_rr3;
  assign t2_r0_c0_rr2 = t1_r0_c0_rr4 + t1_r0_c0_rr5;
  assign t2_r0_c0_rr3 = t1_r0_c0_rr6 + t1_r0_c0_rr7;

  assign t3_r0_c0_rr0 = t2_r0_c0_rr0 + t2_r0_c0_rr1;
  assign t3_r0_c0_rr1 = t2_r0_c0_rr2 + t2_r0_c0_rr3;

  assign t4_r0_c0_rr0 = t3_r0_c0_rr0 + t3_r0_c0_rr1;

  assign c_0_0 = t4_r0_c0_rr0;
  assign t0_r0_c1_rr0 = a_0_0 * b_0_1;
  assign t0_r0_c1_rr1 = a_0_1 * b_1_1;
  assign t0_r0_c1_rr2 = a_0_2 * b_2_1;
  assign t0_r0_c1_rr3 = a_0_3 * b_3_1;
  assign t0_r0_c1_rr4 = a_0_4 * b_4_1;
  assign t0_r0_c1_rr5 = a_0_5 * b_5_1;
  assign t0_r0_c1_rr6 = a_0_6 * b_6_1;
  assign t0_r0_c1_rr7 = a_0_7 * b_7_1;
  assign t0_r0_c1_rr8 = a_0_8 * b_8_1;
  assign t0_r0_c1_rr9 = a_0_9 * b_9_1;
  assign t0_r0_c1_rr10 = a_0_10 * b_10_1;
  assign t0_r0_c1_rr11 = a_0_11 * b_11_1;
  assign t0_r0_c1_rr12 = a_0_12 * b_12_1;
  assign t0_r0_c1_rr13 = a_0_13 * b_13_1;
  assign t0_r0_c1_rr14 = a_0_14 * b_14_1;
  assign t1_r0_c1_rr0 = t0_r0_c1_rr0 + t0_r0_c1_rr1;
  assign t1_r0_c1_rr1 = t0_r0_c1_rr2 + t0_r0_c1_rr3;
  assign t1_r0_c1_rr2 = t0_r0_c1_rr4 + t0_r0_c1_rr5;
  assign t1_r0_c1_rr3 = t0_r0_c1_rr6 + t0_r0_c1_rr7;
  assign t1_r0_c1_rr4 = t0_r0_c1_rr8 + t0_r0_c1_rr9;
  assign t1_r0_c1_rr5 = t0_r0_c1_rr10 + t0_r0_c1_rr11;
  assign t1_r0_c1_rr6 = t0_r0_c1_rr12 + t0_r0_c1_rr13;
  assign t1_r0_c1_rr7 = t0_r0_c1_rr14;

  assign t2_r0_c1_rr0 = t1_r0_c1_rr0 + t1_r0_c1_rr1;
  assign t2_r0_c1_rr1 = t1_r0_c1_rr2 + t1_r0_c1_rr3;
  assign t2_r0_c1_rr2 = t1_r0_c1_rr4 + t1_r0_c1_rr5;
  assign t2_r0_c1_rr3 = t1_r0_c1_rr6 + t1_r0_c1_rr7;

  assign t3_r0_c1_rr0 = t2_r0_c1_rr0 + t2_r0_c1_rr1;
  assign t3_r0_c1_rr1 = t2_r0_c1_rr2 + t2_r0_c1_rr3;

  assign t4_r0_c1_rr0 = t3_r0_c1_rr0 + t3_r0_c1_rr1;

  assign c_0_1 = t4_r0_c1_rr0;
  assign t0_r0_c2_rr0 = a_0_0 * b_0_2;
  assign t0_r0_c2_rr1 = a_0_1 * b_1_2;
  assign t0_r0_c2_rr2 = a_0_2 * b_2_2;
  assign t0_r0_c2_rr3 = a_0_3 * b_3_2;
  assign t0_r0_c2_rr4 = a_0_4 * b_4_2;
  assign t0_r0_c2_rr5 = a_0_5 * b_5_2;
  assign t0_r0_c2_rr6 = a_0_6 * b_6_2;
  assign t0_r0_c2_rr7 = a_0_7 * b_7_2;
  assign t0_r0_c2_rr8 = a_0_8 * b_8_2;
  assign t0_r0_c2_rr9 = a_0_9 * b_9_2;
  assign t0_r0_c2_rr10 = a_0_10 * b_10_2;
  assign t0_r0_c2_rr11 = a_0_11 * b_11_2;
  assign t0_r0_c2_rr12 = a_0_12 * b_12_2;
  assign t0_r0_c2_rr13 = a_0_13 * b_13_2;
  assign t0_r0_c2_rr14 = a_0_14 * b_14_2;
  assign t1_r0_c2_rr0 = t0_r0_c2_rr0 + t0_r0_c2_rr1;
  assign t1_r0_c2_rr1 = t0_r0_c2_rr2 + t0_r0_c2_rr3;
  assign t1_r0_c2_rr2 = t0_r0_c2_rr4 + t0_r0_c2_rr5;
  assign t1_r0_c2_rr3 = t0_r0_c2_rr6 + t0_r0_c2_rr7;
  assign t1_r0_c2_rr4 = t0_r0_c2_rr8 + t0_r0_c2_rr9;
  assign t1_r0_c2_rr5 = t0_r0_c2_rr10 + t0_r0_c2_rr11;
  assign t1_r0_c2_rr6 = t0_r0_c2_rr12 + t0_r0_c2_rr13;
  assign t1_r0_c2_rr7 = t0_r0_c2_rr14;

  assign t2_r0_c2_rr0 = t1_r0_c2_rr0 + t1_r0_c2_rr1;
  assign t2_r0_c2_rr1 = t1_r0_c2_rr2 + t1_r0_c2_rr3;
  assign t2_r0_c2_rr2 = t1_r0_c2_rr4 + t1_r0_c2_rr5;
  assign t2_r0_c2_rr3 = t1_r0_c2_rr6 + t1_r0_c2_rr7;

  assign t3_r0_c2_rr0 = t2_r0_c2_rr0 + t2_r0_c2_rr1;
  assign t3_r0_c2_rr1 = t2_r0_c2_rr2 + t2_r0_c2_rr3;

  assign t4_r0_c2_rr0 = t3_r0_c2_rr0 + t3_r0_c2_rr1;

  assign c_0_2 = t4_r0_c2_rr0;
  assign t0_r0_c3_rr0 = a_0_0 * b_0_3;
  assign t0_r0_c3_rr1 = a_0_1 * b_1_3;
  assign t0_r0_c3_rr2 = a_0_2 * b_2_3;
  assign t0_r0_c3_rr3 = a_0_3 * b_3_3;
  assign t0_r0_c3_rr4 = a_0_4 * b_4_3;
  assign t0_r0_c3_rr5 = a_0_5 * b_5_3;
  assign t0_r0_c3_rr6 = a_0_6 * b_6_3;
  assign t0_r0_c3_rr7 = a_0_7 * b_7_3;
  assign t0_r0_c3_rr8 = a_0_8 * b_8_3;
  assign t0_r0_c3_rr9 = a_0_9 * b_9_3;
  assign t0_r0_c3_rr10 = a_0_10 * b_10_3;
  assign t0_r0_c3_rr11 = a_0_11 * b_11_3;
  assign t0_r0_c3_rr12 = a_0_12 * b_12_3;
  assign t0_r0_c3_rr13 = a_0_13 * b_13_3;
  assign t0_r0_c3_rr14 = a_0_14 * b_14_3;
  assign t1_r0_c3_rr0 = t0_r0_c3_rr0 + t0_r0_c3_rr1;
  assign t1_r0_c3_rr1 = t0_r0_c3_rr2 + t0_r0_c3_rr3;
  assign t1_r0_c3_rr2 = t0_r0_c3_rr4 + t0_r0_c3_rr5;
  assign t1_r0_c3_rr3 = t0_r0_c3_rr6 + t0_r0_c3_rr7;
  assign t1_r0_c3_rr4 = t0_r0_c3_rr8 + t0_r0_c3_rr9;
  assign t1_r0_c3_rr5 = t0_r0_c3_rr10 + t0_r0_c3_rr11;
  assign t1_r0_c3_rr6 = t0_r0_c3_rr12 + t0_r0_c3_rr13;
  assign t1_r0_c3_rr7 = t0_r0_c3_rr14;

  assign t2_r0_c3_rr0 = t1_r0_c3_rr0 + t1_r0_c3_rr1;
  assign t2_r0_c3_rr1 = t1_r0_c3_rr2 + t1_r0_c3_rr3;
  assign t2_r0_c3_rr2 = t1_r0_c3_rr4 + t1_r0_c3_rr5;
  assign t2_r0_c3_rr3 = t1_r0_c3_rr6 + t1_r0_c3_rr7;

  assign t3_r0_c3_rr0 = t2_r0_c3_rr0 + t2_r0_c3_rr1;
  assign t3_r0_c3_rr1 = t2_r0_c3_rr2 + t2_r0_c3_rr3;

  assign t4_r0_c3_rr0 = t3_r0_c3_rr0 + t3_r0_c3_rr1;

  assign c_0_3 = t4_r0_c3_rr0;
  assign t0_r0_c4_rr0 = a_0_0 * b_0_4;
  assign t0_r0_c4_rr1 = a_0_1 * b_1_4;
  assign t0_r0_c4_rr2 = a_0_2 * b_2_4;
  assign t0_r0_c4_rr3 = a_0_3 * b_3_4;
  assign t0_r0_c4_rr4 = a_0_4 * b_4_4;
  assign t0_r0_c4_rr5 = a_0_5 * b_5_4;
  assign t0_r0_c4_rr6 = a_0_6 * b_6_4;
  assign t0_r0_c4_rr7 = a_0_7 * b_7_4;
  assign t0_r0_c4_rr8 = a_0_8 * b_8_4;
  assign t0_r0_c4_rr9 = a_0_9 * b_9_4;
  assign t0_r0_c4_rr10 = a_0_10 * b_10_4;
  assign t0_r0_c4_rr11 = a_0_11 * b_11_4;
  assign t0_r0_c4_rr12 = a_0_12 * b_12_4;
  assign t0_r0_c4_rr13 = a_0_13 * b_13_4;
  assign t0_r0_c4_rr14 = a_0_14 * b_14_4;
  assign t1_r0_c4_rr0 = t0_r0_c4_rr0 + t0_r0_c4_rr1;
  assign t1_r0_c4_rr1 = t0_r0_c4_rr2 + t0_r0_c4_rr3;
  assign t1_r0_c4_rr2 = t0_r0_c4_rr4 + t0_r0_c4_rr5;
  assign t1_r0_c4_rr3 = t0_r0_c4_rr6 + t0_r0_c4_rr7;
  assign t1_r0_c4_rr4 = t0_r0_c4_rr8 + t0_r0_c4_rr9;
  assign t1_r0_c4_rr5 = t0_r0_c4_rr10 + t0_r0_c4_rr11;
  assign t1_r0_c4_rr6 = t0_r0_c4_rr12 + t0_r0_c4_rr13;
  assign t1_r0_c4_rr7 = t0_r0_c4_rr14;

  assign t2_r0_c4_rr0 = t1_r0_c4_rr0 + t1_r0_c4_rr1;
  assign t2_r0_c4_rr1 = t1_r0_c4_rr2 + t1_r0_c4_rr3;
  assign t2_r0_c4_rr2 = t1_r0_c4_rr4 + t1_r0_c4_rr5;
  assign t2_r0_c4_rr3 = t1_r0_c4_rr6 + t1_r0_c4_rr7;

  assign t3_r0_c4_rr0 = t2_r0_c4_rr0 + t2_r0_c4_rr1;
  assign t3_r0_c4_rr1 = t2_r0_c4_rr2 + t2_r0_c4_rr3;

  assign t4_r0_c4_rr0 = t3_r0_c4_rr0 + t3_r0_c4_rr1;

  assign c_0_4 = t4_r0_c4_rr0;
  assign t0_r0_c5_rr0 = a_0_0 * b_0_5;
  assign t0_r0_c5_rr1 = a_0_1 * b_1_5;
  assign t0_r0_c5_rr2 = a_0_2 * b_2_5;
  assign t0_r0_c5_rr3 = a_0_3 * b_3_5;
  assign t0_r0_c5_rr4 = a_0_4 * b_4_5;
  assign t0_r0_c5_rr5 = a_0_5 * b_5_5;
  assign t0_r0_c5_rr6 = a_0_6 * b_6_5;
  assign t0_r0_c5_rr7 = a_0_7 * b_7_5;
  assign t0_r0_c5_rr8 = a_0_8 * b_8_5;
  assign t0_r0_c5_rr9 = a_0_9 * b_9_5;
  assign t0_r0_c5_rr10 = a_0_10 * b_10_5;
  assign t0_r0_c5_rr11 = a_0_11 * b_11_5;
  assign t0_r0_c5_rr12 = a_0_12 * b_12_5;
  assign t0_r0_c5_rr13 = a_0_13 * b_13_5;
  assign t0_r0_c5_rr14 = a_0_14 * b_14_5;
  assign t1_r0_c5_rr0 = t0_r0_c5_rr0 + t0_r0_c5_rr1;
  assign t1_r0_c5_rr1 = t0_r0_c5_rr2 + t0_r0_c5_rr3;
  assign t1_r0_c5_rr2 = t0_r0_c5_rr4 + t0_r0_c5_rr5;
  assign t1_r0_c5_rr3 = t0_r0_c5_rr6 + t0_r0_c5_rr7;
  assign t1_r0_c5_rr4 = t0_r0_c5_rr8 + t0_r0_c5_rr9;
  assign t1_r0_c5_rr5 = t0_r0_c5_rr10 + t0_r0_c5_rr11;
  assign t1_r0_c5_rr6 = t0_r0_c5_rr12 + t0_r0_c5_rr13;
  assign t1_r0_c5_rr7 = t0_r0_c5_rr14;

  assign t2_r0_c5_rr0 = t1_r0_c5_rr0 + t1_r0_c5_rr1;
  assign t2_r0_c5_rr1 = t1_r0_c5_rr2 + t1_r0_c5_rr3;
  assign t2_r0_c5_rr2 = t1_r0_c5_rr4 + t1_r0_c5_rr5;
  assign t2_r0_c5_rr3 = t1_r0_c5_rr6 + t1_r0_c5_rr7;

  assign t3_r0_c5_rr0 = t2_r0_c5_rr0 + t2_r0_c5_rr1;
  assign t3_r0_c5_rr1 = t2_r0_c5_rr2 + t2_r0_c5_rr3;

  assign t4_r0_c5_rr0 = t3_r0_c5_rr0 + t3_r0_c5_rr1;

  assign c_0_5 = t4_r0_c5_rr0;
  assign t0_r0_c6_rr0 = a_0_0 * b_0_6;
  assign t0_r0_c6_rr1 = a_0_1 * b_1_6;
  assign t0_r0_c6_rr2 = a_0_2 * b_2_6;
  assign t0_r0_c6_rr3 = a_0_3 * b_3_6;
  assign t0_r0_c6_rr4 = a_0_4 * b_4_6;
  assign t0_r0_c6_rr5 = a_0_5 * b_5_6;
  assign t0_r0_c6_rr6 = a_0_6 * b_6_6;
  assign t0_r0_c6_rr7 = a_0_7 * b_7_6;
  assign t0_r0_c6_rr8 = a_0_8 * b_8_6;
  assign t0_r0_c6_rr9 = a_0_9 * b_9_6;
  assign t0_r0_c6_rr10 = a_0_10 * b_10_6;
  assign t0_r0_c6_rr11 = a_0_11 * b_11_6;
  assign t0_r0_c6_rr12 = a_0_12 * b_12_6;
  assign t0_r0_c6_rr13 = a_0_13 * b_13_6;
  assign t0_r0_c6_rr14 = a_0_14 * b_14_6;
  assign t1_r0_c6_rr0 = t0_r0_c6_rr0 + t0_r0_c6_rr1;
  assign t1_r0_c6_rr1 = t0_r0_c6_rr2 + t0_r0_c6_rr3;
  assign t1_r0_c6_rr2 = t0_r0_c6_rr4 + t0_r0_c6_rr5;
  assign t1_r0_c6_rr3 = t0_r0_c6_rr6 + t0_r0_c6_rr7;
  assign t1_r0_c6_rr4 = t0_r0_c6_rr8 + t0_r0_c6_rr9;
  assign t1_r0_c6_rr5 = t0_r0_c6_rr10 + t0_r0_c6_rr11;
  assign t1_r0_c6_rr6 = t0_r0_c6_rr12 + t0_r0_c6_rr13;
  assign t1_r0_c6_rr7 = t0_r0_c6_rr14;

  assign t2_r0_c6_rr0 = t1_r0_c6_rr0 + t1_r0_c6_rr1;
  assign t2_r0_c6_rr1 = t1_r0_c6_rr2 + t1_r0_c6_rr3;
  assign t2_r0_c6_rr2 = t1_r0_c6_rr4 + t1_r0_c6_rr5;
  assign t2_r0_c6_rr3 = t1_r0_c6_rr6 + t1_r0_c6_rr7;

  assign t3_r0_c6_rr0 = t2_r0_c6_rr0 + t2_r0_c6_rr1;
  assign t3_r0_c6_rr1 = t2_r0_c6_rr2 + t2_r0_c6_rr3;

  assign t4_r0_c6_rr0 = t3_r0_c6_rr0 + t3_r0_c6_rr1;

  assign c_0_6 = t4_r0_c6_rr0;
  assign t0_r0_c7_rr0 = a_0_0 * b_0_7;
  assign t0_r0_c7_rr1 = a_0_1 * b_1_7;
  assign t0_r0_c7_rr2 = a_0_2 * b_2_7;
  assign t0_r0_c7_rr3 = a_0_3 * b_3_7;
  assign t0_r0_c7_rr4 = a_0_4 * b_4_7;
  assign t0_r0_c7_rr5 = a_0_5 * b_5_7;
  assign t0_r0_c7_rr6 = a_0_6 * b_6_7;
  assign t0_r0_c7_rr7 = a_0_7 * b_7_7;
  assign t0_r0_c7_rr8 = a_0_8 * b_8_7;
  assign t0_r0_c7_rr9 = a_0_9 * b_9_7;
  assign t0_r0_c7_rr10 = a_0_10 * b_10_7;
  assign t0_r0_c7_rr11 = a_0_11 * b_11_7;
  assign t0_r0_c7_rr12 = a_0_12 * b_12_7;
  assign t0_r0_c7_rr13 = a_0_13 * b_13_7;
  assign t0_r0_c7_rr14 = a_0_14 * b_14_7;
  assign t1_r0_c7_rr0 = t0_r0_c7_rr0 + t0_r0_c7_rr1;
  assign t1_r0_c7_rr1 = t0_r0_c7_rr2 + t0_r0_c7_rr3;
  assign t1_r0_c7_rr2 = t0_r0_c7_rr4 + t0_r0_c7_rr5;
  assign t1_r0_c7_rr3 = t0_r0_c7_rr6 + t0_r0_c7_rr7;
  assign t1_r0_c7_rr4 = t0_r0_c7_rr8 + t0_r0_c7_rr9;
  assign t1_r0_c7_rr5 = t0_r0_c7_rr10 + t0_r0_c7_rr11;
  assign t1_r0_c7_rr6 = t0_r0_c7_rr12 + t0_r0_c7_rr13;
  assign t1_r0_c7_rr7 = t0_r0_c7_rr14;

  assign t2_r0_c7_rr0 = t1_r0_c7_rr0 + t1_r0_c7_rr1;
  assign t2_r0_c7_rr1 = t1_r0_c7_rr2 + t1_r0_c7_rr3;
  assign t2_r0_c7_rr2 = t1_r0_c7_rr4 + t1_r0_c7_rr5;
  assign t2_r0_c7_rr3 = t1_r0_c7_rr6 + t1_r0_c7_rr7;

  assign t3_r0_c7_rr0 = t2_r0_c7_rr0 + t2_r0_c7_rr1;
  assign t3_r0_c7_rr1 = t2_r0_c7_rr2 + t2_r0_c7_rr3;

  assign t4_r0_c7_rr0 = t3_r0_c7_rr0 + t3_r0_c7_rr1;

  assign c_0_7 = t4_r0_c7_rr0;
  assign t0_r0_c8_rr0 = a_0_0 * b_0_8;
  assign t0_r0_c8_rr1 = a_0_1 * b_1_8;
  assign t0_r0_c8_rr2 = a_0_2 * b_2_8;
  assign t0_r0_c8_rr3 = a_0_3 * b_3_8;
  assign t0_r0_c8_rr4 = a_0_4 * b_4_8;
  assign t0_r0_c8_rr5 = a_0_5 * b_5_8;
  assign t0_r0_c8_rr6 = a_0_6 * b_6_8;
  assign t0_r0_c8_rr7 = a_0_7 * b_7_8;
  assign t0_r0_c8_rr8 = a_0_8 * b_8_8;
  assign t0_r0_c8_rr9 = a_0_9 * b_9_8;
  assign t0_r0_c8_rr10 = a_0_10 * b_10_8;
  assign t0_r0_c8_rr11 = a_0_11 * b_11_8;
  assign t0_r0_c8_rr12 = a_0_12 * b_12_8;
  assign t0_r0_c8_rr13 = a_0_13 * b_13_8;
  assign t0_r0_c8_rr14 = a_0_14 * b_14_8;
  assign t1_r0_c8_rr0 = t0_r0_c8_rr0 + t0_r0_c8_rr1;
  assign t1_r0_c8_rr1 = t0_r0_c8_rr2 + t0_r0_c8_rr3;
  assign t1_r0_c8_rr2 = t0_r0_c8_rr4 + t0_r0_c8_rr5;
  assign t1_r0_c8_rr3 = t0_r0_c8_rr6 + t0_r0_c8_rr7;
  assign t1_r0_c8_rr4 = t0_r0_c8_rr8 + t0_r0_c8_rr9;
  assign t1_r0_c8_rr5 = t0_r0_c8_rr10 + t0_r0_c8_rr11;
  assign t1_r0_c8_rr6 = t0_r0_c8_rr12 + t0_r0_c8_rr13;
  assign t1_r0_c8_rr7 = t0_r0_c8_rr14;

  assign t2_r0_c8_rr0 = t1_r0_c8_rr0 + t1_r0_c8_rr1;
  assign t2_r0_c8_rr1 = t1_r0_c8_rr2 + t1_r0_c8_rr3;
  assign t2_r0_c8_rr2 = t1_r0_c8_rr4 + t1_r0_c8_rr5;
  assign t2_r0_c8_rr3 = t1_r0_c8_rr6 + t1_r0_c8_rr7;

  assign t3_r0_c8_rr0 = t2_r0_c8_rr0 + t2_r0_c8_rr1;
  assign t3_r0_c8_rr1 = t2_r0_c8_rr2 + t2_r0_c8_rr3;

  assign t4_r0_c8_rr0 = t3_r0_c8_rr0 + t3_r0_c8_rr1;

  assign c_0_8 = t4_r0_c8_rr0;
  assign t0_r0_c9_rr0 = a_0_0 * b_0_9;
  assign t0_r0_c9_rr1 = a_0_1 * b_1_9;
  assign t0_r0_c9_rr2 = a_0_2 * b_2_9;
  assign t0_r0_c9_rr3 = a_0_3 * b_3_9;
  assign t0_r0_c9_rr4 = a_0_4 * b_4_9;
  assign t0_r0_c9_rr5 = a_0_5 * b_5_9;
  assign t0_r0_c9_rr6 = a_0_6 * b_6_9;
  assign t0_r0_c9_rr7 = a_0_7 * b_7_9;
  assign t0_r0_c9_rr8 = a_0_8 * b_8_9;
  assign t0_r0_c9_rr9 = a_0_9 * b_9_9;
  assign t0_r0_c9_rr10 = a_0_10 * b_10_9;
  assign t0_r0_c9_rr11 = a_0_11 * b_11_9;
  assign t0_r0_c9_rr12 = a_0_12 * b_12_9;
  assign t0_r0_c9_rr13 = a_0_13 * b_13_9;
  assign t0_r0_c9_rr14 = a_0_14 * b_14_9;
  assign t1_r0_c9_rr0 = t0_r0_c9_rr0 + t0_r0_c9_rr1;
  assign t1_r0_c9_rr1 = t0_r0_c9_rr2 + t0_r0_c9_rr3;
  assign t1_r0_c9_rr2 = t0_r0_c9_rr4 + t0_r0_c9_rr5;
  assign t1_r0_c9_rr3 = t0_r0_c9_rr6 + t0_r0_c9_rr7;
  assign t1_r0_c9_rr4 = t0_r0_c9_rr8 + t0_r0_c9_rr9;
  assign t1_r0_c9_rr5 = t0_r0_c9_rr10 + t0_r0_c9_rr11;
  assign t1_r0_c9_rr6 = t0_r0_c9_rr12 + t0_r0_c9_rr13;
  assign t1_r0_c9_rr7 = t0_r0_c9_rr14;

  assign t2_r0_c9_rr0 = t1_r0_c9_rr0 + t1_r0_c9_rr1;
  assign t2_r0_c9_rr1 = t1_r0_c9_rr2 + t1_r0_c9_rr3;
  assign t2_r0_c9_rr2 = t1_r0_c9_rr4 + t1_r0_c9_rr5;
  assign t2_r0_c9_rr3 = t1_r0_c9_rr6 + t1_r0_c9_rr7;

  assign t3_r0_c9_rr0 = t2_r0_c9_rr0 + t2_r0_c9_rr1;
  assign t3_r0_c9_rr1 = t2_r0_c9_rr2 + t2_r0_c9_rr3;

  assign t4_r0_c9_rr0 = t3_r0_c9_rr0 + t3_r0_c9_rr1;

  assign c_0_9 = t4_r0_c9_rr0;
  assign t0_r0_c10_rr0 = a_0_0 * b_0_10;
  assign t0_r0_c10_rr1 = a_0_1 * b_1_10;
  assign t0_r0_c10_rr2 = a_0_2 * b_2_10;
  assign t0_r0_c10_rr3 = a_0_3 * b_3_10;
  assign t0_r0_c10_rr4 = a_0_4 * b_4_10;
  assign t0_r0_c10_rr5 = a_0_5 * b_5_10;
  assign t0_r0_c10_rr6 = a_0_6 * b_6_10;
  assign t0_r0_c10_rr7 = a_0_7 * b_7_10;
  assign t0_r0_c10_rr8 = a_0_8 * b_8_10;
  assign t0_r0_c10_rr9 = a_0_9 * b_9_10;
  assign t0_r0_c10_rr10 = a_0_10 * b_10_10;
  assign t0_r0_c10_rr11 = a_0_11 * b_11_10;
  assign t0_r0_c10_rr12 = a_0_12 * b_12_10;
  assign t0_r0_c10_rr13 = a_0_13 * b_13_10;
  assign t0_r0_c10_rr14 = a_0_14 * b_14_10;
  assign t1_r0_c10_rr0 = t0_r0_c10_rr0 + t0_r0_c10_rr1;
  assign t1_r0_c10_rr1 = t0_r0_c10_rr2 + t0_r0_c10_rr3;
  assign t1_r0_c10_rr2 = t0_r0_c10_rr4 + t0_r0_c10_rr5;
  assign t1_r0_c10_rr3 = t0_r0_c10_rr6 + t0_r0_c10_rr7;
  assign t1_r0_c10_rr4 = t0_r0_c10_rr8 + t0_r0_c10_rr9;
  assign t1_r0_c10_rr5 = t0_r0_c10_rr10 + t0_r0_c10_rr11;
  assign t1_r0_c10_rr6 = t0_r0_c10_rr12 + t0_r0_c10_rr13;
  assign t1_r0_c10_rr7 = t0_r0_c10_rr14;

  assign t2_r0_c10_rr0 = t1_r0_c10_rr0 + t1_r0_c10_rr1;
  assign t2_r0_c10_rr1 = t1_r0_c10_rr2 + t1_r0_c10_rr3;
  assign t2_r0_c10_rr2 = t1_r0_c10_rr4 + t1_r0_c10_rr5;
  assign t2_r0_c10_rr3 = t1_r0_c10_rr6 + t1_r0_c10_rr7;

  assign t3_r0_c10_rr0 = t2_r0_c10_rr0 + t2_r0_c10_rr1;
  assign t3_r0_c10_rr1 = t2_r0_c10_rr2 + t2_r0_c10_rr3;

  assign t4_r0_c10_rr0 = t3_r0_c10_rr0 + t3_r0_c10_rr1;

  assign c_0_10 = t4_r0_c10_rr0;
  assign t0_r0_c11_rr0 = a_0_0 * b_0_11;
  assign t0_r0_c11_rr1 = a_0_1 * b_1_11;
  assign t0_r0_c11_rr2 = a_0_2 * b_2_11;
  assign t0_r0_c11_rr3 = a_0_3 * b_3_11;
  assign t0_r0_c11_rr4 = a_0_4 * b_4_11;
  assign t0_r0_c11_rr5 = a_0_5 * b_5_11;
  assign t0_r0_c11_rr6 = a_0_6 * b_6_11;
  assign t0_r0_c11_rr7 = a_0_7 * b_7_11;
  assign t0_r0_c11_rr8 = a_0_8 * b_8_11;
  assign t0_r0_c11_rr9 = a_0_9 * b_9_11;
  assign t0_r0_c11_rr10 = a_0_10 * b_10_11;
  assign t0_r0_c11_rr11 = a_0_11 * b_11_11;
  assign t0_r0_c11_rr12 = a_0_12 * b_12_11;
  assign t0_r0_c11_rr13 = a_0_13 * b_13_11;
  assign t0_r0_c11_rr14 = a_0_14 * b_14_11;
  assign t1_r0_c11_rr0 = t0_r0_c11_rr0 + t0_r0_c11_rr1;
  assign t1_r0_c11_rr1 = t0_r0_c11_rr2 + t0_r0_c11_rr3;
  assign t1_r0_c11_rr2 = t0_r0_c11_rr4 + t0_r0_c11_rr5;
  assign t1_r0_c11_rr3 = t0_r0_c11_rr6 + t0_r0_c11_rr7;
  assign t1_r0_c11_rr4 = t0_r0_c11_rr8 + t0_r0_c11_rr9;
  assign t1_r0_c11_rr5 = t0_r0_c11_rr10 + t0_r0_c11_rr11;
  assign t1_r0_c11_rr6 = t0_r0_c11_rr12 + t0_r0_c11_rr13;
  assign t1_r0_c11_rr7 = t0_r0_c11_rr14;

  assign t2_r0_c11_rr0 = t1_r0_c11_rr0 + t1_r0_c11_rr1;
  assign t2_r0_c11_rr1 = t1_r0_c11_rr2 + t1_r0_c11_rr3;
  assign t2_r0_c11_rr2 = t1_r0_c11_rr4 + t1_r0_c11_rr5;
  assign t2_r0_c11_rr3 = t1_r0_c11_rr6 + t1_r0_c11_rr7;

  assign t3_r0_c11_rr0 = t2_r0_c11_rr0 + t2_r0_c11_rr1;
  assign t3_r0_c11_rr1 = t2_r0_c11_rr2 + t2_r0_c11_rr3;

  assign t4_r0_c11_rr0 = t3_r0_c11_rr0 + t3_r0_c11_rr1;

  assign c_0_11 = t4_r0_c11_rr0;
  assign t0_r0_c12_rr0 = a_0_0 * b_0_12;
  assign t0_r0_c12_rr1 = a_0_1 * b_1_12;
  assign t0_r0_c12_rr2 = a_0_2 * b_2_12;
  assign t0_r0_c12_rr3 = a_0_3 * b_3_12;
  assign t0_r0_c12_rr4 = a_0_4 * b_4_12;
  assign t0_r0_c12_rr5 = a_0_5 * b_5_12;
  assign t0_r0_c12_rr6 = a_0_6 * b_6_12;
  assign t0_r0_c12_rr7 = a_0_7 * b_7_12;
  assign t0_r0_c12_rr8 = a_0_8 * b_8_12;
  assign t0_r0_c12_rr9 = a_0_9 * b_9_12;
  assign t0_r0_c12_rr10 = a_0_10 * b_10_12;
  assign t0_r0_c12_rr11 = a_0_11 * b_11_12;
  assign t0_r0_c12_rr12 = a_0_12 * b_12_12;
  assign t0_r0_c12_rr13 = a_0_13 * b_13_12;
  assign t0_r0_c12_rr14 = a_0_14 * b_14_12;
  assign t1_r0_c12_rr0 = t0_r0_c12_rr0 + t0_r0_c12_rr1;
  assign t1_r0_c12_rr1 = t0_r0_c12_rr2 + t0_r0_c12_rr3;
  assign t1_r0_c12_rr2 = t0_r0_c12_rr4 + t0_r0_c12_rr5;
  assign t1_r0_c12_rr3 = t0_r0_c12_rr6 + t0_r0_c12_rr7;
  assign t1_r0_c12_rr4 = t0_r0_c12_rr8 + t0_r0_c12_rr9;
  assign t1_r0_c12_rr5 = t0_r0_c12_rr10 + t0_r0_c12_rr11;
  assign t1_r0_c12_rr6 = t0_r0_c12_rr12 + t0_r0_c12_rr13;
  assign t1_r0_c12_rr7 = t0_r0_c12_rr14;

  assign t2_r0_c12_rr0 = t1_r0_c12_rr0 + t1_r0_c12_rr1;
  assign t2_r0_c12_rr1 = t1_r0_c12_rr2 + t1_r0_c12_rr3;
  assign t2_r0_c12_rr2 = t1_r0_c12_rr4 + t1_r0_c12_rr5;
  assign t2_r0_c12_rr3 = t1_r0_c12_rr6 + t1_r0_c12_rr7;

  assign t3_r0_c12_rr0 = t2_r0_c12_rr0 + t2_r0_c12_rr1;
  assign t3_r0_c12_rr1 = t2_r0_c12_rr2 + t2_r0_c12_rr3;

  assign t4_r0_c12_rr0 = t3_r0_c12_rr0 + t3_r0_c12_rr1;

  assign c_0_12 = t4_r0_c12_rr0;
  assign t0_r0_c13_rr0 = a_0_0 * b_0_13;
  assign t0_r0_c13_rr1 = a_0_1 * b_1_13;
  assign t0_r0_c13_rr2 = a_0_2 * b_2_13;
  assign t0_r0_c13_rr3 = a_0_3 * b_3_13;
  assign t0_r0_c13_rr4 = a_0_4 * b_4_13;
  assign t0_r0_c13_rr5 = a_0_5 * b_5_13;
  assign t0_r0_c13_rr6 = a_0_6 * b_6_13;
  assign t0_r0_c13_rr7 = a_0_7 * b_7_13;
  assign t0_r0_c13_rr8 = a_0_8 * b_8_13;
  assign t0_r0_c13_rr9 = a_0_9 * b_9_13;
  assign t0_r0_c13_rr10 = a_0_10 * b_10_13;
  assign t0_r0_c13_rr11 = a_0_11 * b_11_13;
  assign t0_r0_c13_rr12 = a_0_12 * b_12_13;
  assign t0_r0_c13_rr13 = a_0_13 * b_13_13;
  assign t0_r0_c13_rr14 = a_0_14 * b_14_13;
  assign t1_r0_c13_rr0 = t0_r0_c13_rr0 + t0_r0_c13_rr1;
  assign t1_r0_c13_rr1 = t0_r0_c13_rr2 + t0_r0_c13_rr3;
  assign t1_r0_c13_rr2 = t0_r0_c13_rr4 + t0_r0_c13_rr5;
  assign t1_r0_c13_rr3 = t0_r0_c13_rr6 + t0_r0_c13_rr7;
  assign t1_r0_c13_rr4 = t0_r0_c13_rr8 + t0_r0_c13_rr9;
  assign t1_r0_c13_rr5 = t0_r0_c13_rr10 + t0_r0_c13_rr11;
  assign t1_r0_c13_rr6 = t0_r0_c13_rr12 + t0_r0_c13_rr13;
  assign t1_r0_c13_rr7 = t0_r0_c13_rr14;

  assign t2_r0_c13_rr0 = t1_r0_c13_rr0 + t1_r0_c13_rr1;
  assign t2_r0_c13_rr1 = t1_r0_c13_rr2 + t1_r0_c13_rr3;
  assign t2_r0_c13_rr2 = t1_r0_c13_rr4 + t1_r0_c13_rr5;
  assign t2_r0_c13_rr3 = t1_r0_c13_rr6 + t1_r0_c13_rr7;

  assign t3_r0_c13_rr0 = t2_r0_c13_rr0 + t2_r0_c13_rr1;
  assign t3_r0_c13_rr1 = t2_r0_c13_rr2 + t2_r0_c13_rr3;

  assign t4_r0_c13_rr0 = t3_r0_c13_rr0 + t3_r0_c13_rr1;

  assign c_0_13 = t4_r0_c13_rr0;
  assign t0_r0_c14_rr0 = a_0_0 * b_0_14;
  assign t0_r0_c14_rr1 = a_0_1 * b_1_14;
  assign t0_r0_c14_rr2 = a_0_2 * b_2_14;
  assign t0_r0_c14_rr3 = a_0_3 * b_3_14;
  assign t0_r0_c14_rr4 = a_0_4 * b_4_14;
  assign t0_r0_c14_rr5 = a_0_5 * b_5_14;
  assign t0_r0_c14_rr6 = a_0_6 * b_6_14;
  assign t0_r0_c14_rr7 = a_0_7 * b_7_14;
  assign t0_r0_c14_rr8 = a_0_8 * b_8_14;
  assign t0_r0_c14_rr9 = a_0_9 * b_9_14;
  assign t0_r0_c14_rr10 = a_0_10 * b_10_14;
  assign t0_r0_c14_rr11 = a_0_11 * b_11_14;
  assign t0_r0_c14_rr12 = a_0_12 * b_12_14;
  assign t0_r0_c14_rr13 = a_0_13 * b_13_14;
  assign t0_r0_c14_rr14 = a_0_14 * b_14_14;
  assign t1_r0_c14_rr0 = t0_r0_c14_rr0 + t0_r0_c14_rr1;
  assign t1_r0_c14_rr1 = t0_r0_c14_rr2 + t0_r0_c14_rr3;
  assign t1_r0_c14_rr2 = t0_r0_c14_rr4 + t0_r0_c14_rr5;
  assign t1_r0_c14_rr3 = t0_r0_c14_rr6 + t0_r0_c14_rr7;
  assign t1_r0_c14_rr4 = t0_r0_c14_rr8 + t0_r0_c14_rr9;
  assign t1_r0_c14_rr5 = t0_r0_c14_rr10 + t0_r0_c14_rr11;
  assign t1_r0_c14_rr6 = t0_r0_c14_rr12 + t0_r0_c14_rr13;
  assign t1_r0_c14_rr7 = t0_r0_c14_rr14;

  assign t2_r0_c14_rr0 = t1_r0_c14_rr0 + t1_r0_c14_rr1;
  assign t2_r0_c14_rr1 = t1_r0_c14_rr2 + t1_r0_c14_rr3;
  assign t2_r0_c14_rr2 = t1_r0_c14_rr4 + t1_r0_c14_rr5;
  assign t2_r0_c14_rr3 = t1_r0_c14_rr6 + t1_r0_c14_rr7;

  assign t3_r0_c14_rr0 = t2_r0_c14_rr0 + t2_r0_c14_rr1;
  assign t3_r0_c14_rr1 = t2_r0_c14_rr2 + t2_r0_c14_rr3;

  assign t4_r0_c14_rr0 = t3_r0_c14_rr0 + t3_r0_c14_rr1;

  assign c_0_14 = t4_r0_c14_rr0;
  assign t0_r1_c0_rr0 = a_1_0 * b_0_0;
  assign t0_r1_c0_rr1 = a_1_1 * b_1_0;
  assign t0_r1_c0_rr2 = a_1_2 * b_2_0;
  assign t0_r1_c0_rr3 = a_1_3 * b_3_0;
  assign t0_r1_c0_rr4 = a_1_4 * b_4_0;
  assign t0_r1_c0_rr5 = a_1_5 * b_5_0;
  assign t0_r1_c0_rr6 = a_1_6 * b_6_0;
  assign t0_r1_c0_rr7 = a_1_7 * b_7_0;
  assign t0_r1_c0_rr8 = a_1_8 * b_8_0;
  assign t0_r1_c0_rr9 = a_1_9 * b_9_0;
  assign t0_r1_c0_rr10 = a_1_10 * b_10_0;
  assign t0_r1_c0_rr11 = a_1_11 * b_11_0;
  assign t0_r1_c0_rr12 = a_1_12 * b_12_0;
  assign t0_r1_c0_rr13 = a_1_13 * b_13_0;
  assign t0_r1_c0_rr14 = a_1_14 * b_14_0;
  assign t1_r1_c0_rr0 = t0_r1_c0_rr0 + t0_r1_c0_rr1;
  assign t1_r1_c0_rr1 = t0_r1_c0_rr2 + t0_r1_c0_rr3;
  assign t1_r1_c0_rr2 = t0_r1_c0_rr4 + t0_r1_c0_rr5;
  assign t1_r1_c0_rr3 = t0_r1_c0_rr6 + t0_r1_c0_rr7;
  assign t1_r1_c0_rr4 = t0_r1_c0_rr8 + t0_r1_c0_rr9;
  assign t1_r1_c0_rr5 = t0_r1_c0_rr10 + t0_r1_c0_rr11;
  assign t1_r1_c0_rr6 = t0_r1_c0_rr12 + t0_r1_c0_rr13;
  assign t1_r1_c0_rr7 = t0_r1_c0_rr14;

  assign t2_r1_c0_rr0 = t1_r1_c0_rr0 + t1_r1_c0_rr1;
  assign t2_r1_c0_rr1 = t1_r1_c0_rr2 + t1_r1_c0_rr3;
  assign t2_r1_c0_rr2 = t1_r1_c0_rr4 + t1_r1_c0_rr5;
  assign t2_r1_c0_rr3 = t1_r1_c0_rr6 + t1_r1_c0_rr7;

  assign t3_r1_c0_rr0 = t2_r1_c0_rr0 + t2_r1_c0_rr1;
  assign t3_r1_c0_rr1 = t2_r1_c0_rr2 + t2_r1_c0_rr3;

  assign t4_r1_c0_rr0 = t3_r1_c0_rr0 + t3_r1_c0_rr1;

  assign c_1_0 = t4_r1_c0_rr0;
  assign t0_r1_c1_rr0 = a_1_0 * b_0_1;
  assign t0_r1_c1_rr1 = a_1_1 * b_1_1;
  assign t0_r1_c1_rr2 = a_1_2 * b_2_1;
  assign t0_r1_c1_rr3 = a_1_3 * b_3_1;
  assign t0_r1_c1_rr4 = a_1_4 * b_4_1;
  assign t0_r1_c1_rr5 = a_1_5 * b_5_1;
  assign t0_r1_c1_rr6 = a_1_6 * b_6_1;
  assign t0_r1_c1_rr7 = a_1_7 * b_7_1;
  assign t0_r1_c1_rr8 = a_1_8 * b_8_1;
  assign t0_r1_c1_rr9 = a_1_9 * b_9_1;
  assign t0_r1_c1_rr10 = a_1_10 * b_10_1;
  assign t0_r1_c1_rr11 = a_1_11 * b_11_1;
  assign t0_r1_c1_rr12 = a_1_12 * b_12_1;
  assign t0_r1_c1_rr13 = a_1_13 * b_13_1;
  assign t0_r1_c1_rr14 = a_1_14 * b_14_1;
  assign t1_r1_c1_rr0 = t0_r1_c1_rr0 + t0_r1_c1_rr1;
  assign t1_r1_c1_rr1 = t0_r1_c1_rr2 + t0_r1_c1_rr3;
  assign t1_r1_c1_rr2 = t0_r1_c1_rr4 + t0_r1_c1_rr5;
  assign t1_r1_c1_rr3 = t0_r1_c1_rr6 + t0_r1_c1_rr7;
  assign t1_r1_c1_rr4 = t0_r1_c1_rr8 + t0_r1_c1_rr9;
  assign t1_r1_c1_rr5 = t0_r1_c1_rr10 + t0_r1_c1_rr11;
  assign t1_r1_c1_rr6 = t0_r1_c1_rr12 + t0_r1_c1_rr13;
  assign t1_r1_c1_rr7 = t0_r1_c1_rr14;

  assign t2_r1_c1_rr0 = t1_r1_c1_rr0 + t1_r1_c1_rr1;
  assign t2_r1_c1_rr1 = t1_r1_c1_rr2 + t1_r1_c1_rr3;
  assign t2_r1_c1_rr2 = t1_r1_c1_rr4 + t1_r1_c1_rr5;
  assign t2_r1_c1_rr3 = t1_r1_c1_rr6 + t1_r1_c1_rr7;

  assign t3_r1_c1_rr0 = t2_r1_c1_rr0 + t2_r1_c1_rr1;
  assign t3_r1_c1_rr1 = t2_r1_c1_rr2 + t2_r1_c1_rr3;

  assign t4_r1_c1_rr0 = t3_r1_c1_rr0 + t3_r1_c1_rr1;

  assign c_1_1 = t4_r1_c1_rr0;
  assign t0_r1_c2_rr0 = a_1_0 * b_0_2;
  assign t0_r1_c2_rr1 = a_1_1 * b_1_2;
  assign t0_r1_c2_rr2 = a_1_2 * b_2_2;
  assign t0_r1_c2_rr3 = a_1_3 * b_3_2;
  assign t0_r1_c2_rr4 = a_1_4 * b_4_2;
  assign t0_r1_c2_rr5 = a_1_5 * b_5_2;
  assign t0_r1_c2_rr6 = a_1_6 * b_6_2;
  assign t0_r1_c2_rr7 = a_1_7 * b_7_2;
  assign t0_r1_c2_rr8 = a_1_8 * b_8_2;
  assign t0_r1_c2_rr9 = a_1_9 * b_9_2;
  assign t0_r1_c2_rr10 = a_1_10 * b_10_2;
  assign t0_r1_c2_rr11 = a_1_11 * b_11_2;
  assign t0_r1_c2_rr12 = a_1_12 * b_12_2;
  assign t0_r1_c2_rr13 = a_1_13 * b_13_2;
  assign t0_r1_c2_rr14 = a_1_14 * b_14_2;
  assign t1_r1_c2_rr0 = t0_r1_c2_rr0 + t0_r1_c2_rr1;
  assign t1_r1_c2_rr1 = t0_r1_c2_rr2 + t0_r1_c2_rr3;
  assign t1_r1_c2_rr2 = t0_r1_c2_rr4 + t0_r1_c2_rr5;
  assign t1_r1_c2_rr3 = t0_r1_c2_rr6 + t0_r1_c2_rr7;
  assign t1_r1_c2_rr4 = t0_r1_c2_rr8 + t0_r1_c2_rr9;
  assign t1_r1_c2_rr5 = t0_r1_c2_rr10 + t0_r1_c2_rr11;
  assign t1_r1_c2_rr6 = t0_r1_c2_rr12 + t0_r1_c2_rr13;
  assign t1_r1_c2_rr7 = t0_r1_c2_rr14;

  assign t2_r1_c2_rr0 = t1_r1_c2_rr0 + t1_r1_c2_rr1;
  assign t2_r1_c2_rr1 = t1_r1_c2_rr2 + t1_r1_c2_rr3;
  assign t2_r1_c2_rr2 = t1_r1_c2_rr4 + t1_r1_c2_rr5;
  assign t2_r1_c2_rr3 = t1_r1_c2_rr6 + t1_r1_c2_rr7;

  assign t3_r1_c2_rr0 = t2_r1_c2_rr0 + t2_r1_c2_rr1;
  assign t3_r1_c2_rr1 = t2_r1_c2_rr2 + t2_r1_c2_rr3;

  assign t4_r1_c2_rr0 = t3_r1_c2_rr0 + t3_r1_c2_rr1;

  assign c_1_2 = t4_r1_c2_rr0;
  assign t0_r1_c3_rr0 = a_1_0 * b_0_3;
  assign t0_r1_c3_rr1 = a_1_1 * b_1_3;
  assign t0_r1_c3_rr2 = a_1_2 * b_2_3;
  assign t0_r1_c3_rr3 = a_1_3 * b_3_3;
  assign t0_r1_c3_rr4 = a_1_4 * b_4_3;
  assign t0_r1_c3_rr5 = a_1_5 * b_5_3;
  assign t0_r1_c3_rr6 = a_1_6 * b_6_3;
  assign t0_r1_c3_rr7 = a_1_7 * b_7_3;
  assign t0_r1_c3_rr8 = a_1_8 * b_8_3;
  assign t0_r1_c3_rr9 = a_1_9 * b_9_3;
  assign t0_r1_c3_rr10 = a_1_10 * b_10_3;
  assign t0_r1_c3_rr11 = a_1_11 * b_11_3;
  assign t0_r1_c3_rr12 = a_1_12 * b_12_3;
  assign t0_r1_c3_rr13 = a_1_13 * b_13_3;
  assign t0_r1_c3_rr14 = a_1_14 * b_14_3;
  assign t1_r1_c3_rr0 = t0_r1_c3_rr0 + t0_r1_c3_rr1;
  assign t1_r1_c3_rr1 = t0_r1_c3_rr2 + t0_r1_c3_rr3;
  assign t1_r1_c3_rr2 = t0_r1_c3_rr4 + t0_r1_c3_rr5;
  assign t1_r1_c3_rr3 = t0_r1_c3_rr6 + t0_r1_c3_rr7;
  assign t1_r1_c3_rr4 = t0_r1_c3_rr8 + t0_r1_c3_rr9;
  assign t1_r1_c3_rr5 = t0_r1_c3_rr10 + t0_r1_c3_rr11;
  assign t1_r1_c3_rr6 = t0_r1_c3_rr12 + t0_r1_c3_rr13;
  assign t1_r1_c3_rr7 = t0_r1_c3_rr14;

  assign t2_r1_c3_rr0 = t1_r1_c3_rr0 + t1_r1_c3_rr1;
  assign t2_r1_c3_rr1 = t1_r1_c3_rr2 + t1_r1_c3_rr3;
  assign t2_r1_c3_rr2 = t1_r1_c3_rr4 + t1_r1_c3_rr5;
  assign t2_r1_c3_rr3 = t1_r1_c3_rr6 + t1_r1_c3_rr7;

  assign t3_r1_c3_rr0 = t2_r1_c3_rr0 + t2_r1_c3_rr1;
  assign t3_r1_c3_rr1 = t2_r1_c3_rr2 + t2_r1_c3_rr3;

  assign t4_r1_c3_rr0 = t3_r1_c3_rr0 + t3_r1_c3_rr1;

  assign c_1_3 = t4_r1_c3_rr0;
  assign t0_r1_c4_rr0 = a_1_0 * b_0_4;
  assign t0_r1_c4_rr1 = a_1_1 * b_1_4;
  assign t0_r1_c4_rr2 = a_1_2 * b_2_4;
  assign t0_r1_c4_rr3 = a_1_3 * b_3_4;
  assign t0_r1_c4_rr4 = a_1_4 * b_4_4;
  assign t0_r1_c4_rr5 = a_1_5 * b_5_4;
  assign t0_r1_c4_rr6 = a_1_6 * b_6_4;
  assign t0_r1_c4_rr7 = a_1_7 * b_7_4;
  assign t0_r1_c4_rr8 = a_1_8 * b_8_4;
  assign t0_r1_c4_rr9 = a_1_9 * b_9_4;
  assign t0_r1_c4_rr10 = a_1_10 * b_10_4;
  assign t0_r1_c4_rr11 = a_1_11 * b_11_4;
  assign t0_r1_c4_rr12 = a_1_12 * b_12_4;
  assign t0_r1_c4_rr13 = a_1_13 * b_13_4;
  assign t0_r1_c4_rr14 = a_1_14 * b_14_4;
  assign t1_r1_c4_rr0 = t0_r1_c4_rr0 + t0_r1_c4_rr1;
  assign t1_r1_c4_rr1 = t0_r1_c4_rr2 + t0_r1_c4_rr3;
  assign t1_r1_c4_rr2 = t0_r1_c4_rr4 + t0_r1_c4_rr5;
  assign t1_r1_c4_rr3 = t0_r1_c4_rr6 + t0_r1_c4_rr7;
  assign t1_r1_c4_rr4 = t0_r1_c4_rr8 + t0_r1_c4_rr9;
  assign t1_r1_c4_rr5 = t0_r1_c4_rr10 + t0_r1_c4_rr11;
  assign t1_r1_c4_rr6 = t0_r1_c4_rr12 + t0_r1_c4_rr13;
  assign t1_r1_c4_rr7 = t0_r1_c4_rr14;

  assign t2_r1_c4_rr0 = t1_r1_c4_rr0 + t1_r1_c4_rr1;
  assign t2_r1_c4_rr1 = t1_r1_c4_rr2 + t1_r1_c4_rr3;
  assign t2_r1_c4_rr2 = t1_r1_c4_rr4 + t1_r1_c4_rr5;
  assign t2_r1_c4_rr3 = t1_r1_c4_rr6 + t1_r1_c4_rr7;

  assign t3_r1_c4_rr0 = t2_r1_c4_rr0 + t2_r1_c4_rr1;
  assign t3_r1_c4_rr1 = t2_r1_c4_rr2 + t2_r1_c4_rr3;

  assign t4_r1_c4_rr0 = t3_r1_c4_rr0 + t3_r1_c4_rr1;

  assign c_1_4 = t4_r1_c4_rr0;
  assign t0_r1_c5_rr0 = a_1_0 * b_0_5;
  assign t0_r1_c5_rr1 = a_1_1 * b_1_5;
  assign t0_r1_c5_rr2 = a_1_2 * b_2_5;
  assign t0_r1_c5_rr3 = a_1_3 * b_3_5;
  assign t0_r1_c5_rr4 = a_1_4 * b_4_5;
  assign t0_r1_c5_rr5 = a_1_5 * b_5_5;
  assign t0_r1_c5_rr6 = a_1_6 * b_6_5;
  assign t0_r1_c5_rr7 = a_1_7 * b_7_5;
  assign t0_r1_c5_rr8 = a_1_8 * b_8_5;
  assign t0_r1_c5_rr9 = a_1_9 * b_9_5;
  assign t0_r1_c5_rr10 = a_1_10 * b_10_5;
  assign t0_r1_c5_rr11 = a_1_11 * b_11_5;
  assign t0_r1_c5_rr12 = a_1_12 * b_12_5;
  assign t0_r1_c5_rr13 = a_1_13 * b_13_5;
  assign t0_r1_c5_rr14 = a_1_14 * b_14_5;
  assign t1_r1_c5_rr0 = t0_r1_c5_rr0 + t0_r1_c5_rr1;
  assign t1_r1_c5_rr1 = t0_r1_c5_rr2 + t0_r1_c5_rr3;
  assign t1_r1_c5_rr2 = t0_r1_c5_rr4 + t0_r1_c5_rr5;
  assign t1_r1_c5_rr3 = t0_r1_c5_rr6 + t0_r1_c5_rr7;
  assign t1_r1_c5_rr4 = t0_r1_c5_rr8 + t0_r1_c5_rr9;
  assign t1_r1_c5_rr5 = t0_r1_c5_rr10 + t0_r1_c5_rr11;
  assign t1_r1_c5_rr6 = t0_r1_c5_rr12 + t0_r1_c5_rr13;
  assign t1_r1_c5_rr7 = t0_r1_c5_rr14;

  assign t2_r1_c5_rr0 = t1_r1_c5_rr0 + t1_r1_c5_rr1;
  assign t2_r1_c5_rr1 = t1_r1_c5_rr2 + t1_r1_c5_rr3;
  assign t2_r1_c5_rr2 = t1_r1_c5_rr4 + t1_r1_c5_rr5;
  assign t2_r1_c5_rr3 = t1_r1_c5_rr6 + t1_r1_c5_rr7;

  assign t3_r1_c5_rr0 = t2_r1_c5_rr0 + t2_r1_c5_rr1;
  assign t3_r1_c5_rr1 = t2_r1_c5_rr2 + t2_r1_c5_rr3;

  assign t4_r1_c5_rr0 = t3_r1_c5_rr0 + t3_r1_c5_rr1;

  assign c_1_5 = t4_r1_c5_rr0;
  assign t0_r1_c6_rr0 = a_1_0 * b_0_6;
  assign t0_r1_c6_rr1 = a_1_1 * b_1_6;
  assign t0_r1_c6_rr2 = a_1_2 * b_2_6;
  assign t0_r1_c6_rr3 = a_1_3 * b_3_6;
  assign t0_r1_c6_rr4 = a_1_4 * b_4_6;
  assign t0_r1_c6_rr5 = a_1_5 * b_5_6;
  assign t0_r1_c6_rr6 = a_1_6 * b_6_6;
  assign t0_r1_c6_rr7 = a_1_7 * b_7_6;
  assign t0_r1_c6_rr8 = a_1_8 * b_8_6;
  assign t0_r1_c6_rr9 = a_1_9 * b_9_6;
  assign t0_r1_c6_rr10 = a_1_10 * b_10_6;
  assign t0_r1_c6_rr11 = a_1_11 * b_11_6;
  assign t0_r1_c6_rr12 = a_1_12 * b_12_6;
  assign t0_r1_c6_rr13 = a_1_13 * b_13_6;
  assign t0_r1_c6_rr14 = a_1_14 * b_14_6;
  assign t1_r1_c6_rr0 = t0_r1_c6_rr0 + t0_r1_c6_rr1;
  assign t1_r1_c6_rr1 = t0_r1_c6_rr2 + t0_r1_c6_rr3;
  assign t1_r1_c6_rr2 = t0_r1_c6_rr4 + t0_r1_c6_rr5;
  assign t1_r1_c6_rr3 = t0_r1_c6_rr6 + t0_r1_c6_rr7;
  assign t1_r1_c6_rr4 = t0_r1_c6_rr8 + t0_r1_c6_rr9;
  assign t1_r1_c6_rr5 = t0_r1_c6_rr10 + t0_r1_c6_rr11;
  assign t1_r1_c6_rr6 = t0_r1_c6_rr12 + t0_r1_c6_rr13;
  assign t1_r1_c6_rr7 = t0_r1_c6_rr14;

  assign t2_r1_c6_rr0 = t1_r1_c6_rr0 + t1_r1_c6_rr1;
  assign t2_r1_c6_rr1 = t1_r1_c6_rr2 + t1_r1_c6_rr3;
  assign t2_r1_c6_rr2 = t1_r1_c6_rr4 + t1_r1_c6_rr5;
  assign t2_r1_c6_rr3 = t1_r1_c6_rr6 + t1_r1_c6_rr7;

  assign t3_r1_c6_rr0 = t2_r1_c6_rr0 + t2_r1_c6_rr1;
  assign t3_r1_c6_rr1 = t2_r1_c6_rr2 + t2_r1_c6_rr3;

  assign t4_r1_c6_rr0 = t3_r1_c6_rr0 + t3_r1_c6_rr1;

  assign c_1_6 = t4_r1_c6_rr0;
  assign t0_r1_c7_rr0 = a_1_0 * b_0_7;
  assign t0_r1_c7_rr1 = a_1_1 * b_1_7;
  assign t0_r1_c7_rr2 = a_1_2 * b_2_7;
  assign t0_r1_c7_rr3 = a_1_3 * b_3_7;
  assign t0_r1_c7_rr4 = a_1_4 * b_4_7;
  assign t0_r1_c7_rr5 = a_1_5 * b_5_7;
  assign t0_r1_c7_rr6 = a_1_6 * b_6_7;
  assign t0_r1_c7_rr7 = a_1_7 * b_7_7;
  assign t0_r1_c7_rr8 = a_1_8 * b_8_7;
  assign t0_r1_c7_rr9 = a_1_9 * b_9_7;
  assign t0_r1_c7_rr10 = a_1_10 * b_10_7;
  assign t0_r1_c7_rr11 = a_1_11 * b_11_7;
  assign t0_r1_c7_rr12 = a_1_12 * b_12_7;
  assign t0_r1_c7_rr13 = a_1_13 * b_13_7;
  assign t0_r1_c7_rr14 = a_1_14 * b_14_7;
  assign t1_r1_c7_rr0 = t0_r1_c7_rr0 + t0_r1_c7_rr1;
  assign t1_r1_c7_rr1 = t0_r1_c7_rr2 + t0_r1_c7_rr3;
  assign t1_r1_c7_rr2 = t0_r1_c7_rr4 + t0_r1_c7_rr5;
  assign t1_r1_c7_rr3 = t0_r1_c7_rr6 + t0_r1_c7_rr7;
  assign t1_r1_c7_rr4 = t0_r1_c7_rr8 + t0_r1_c7_rr9;
  assign t1_r1_c7_rr5 = t0_r1_c7_rr10 + t0_r1_c7_rr11;
  assign t1_r1_c7_rr6 = t0_r1_c7_rr12 + t0_r1_c7_rr13;
  assign t1_r1_c7_rr7 = t0_r1_c7_rr14;

  assign t2_r1_c7_rr0 = t1_r1_c7_rr0 + t1_r1_c7_rr1;
  assign t2_r1_c7_rr1 = t1_r1_c7_rr2 + t1_r1_c7_rr3;
  assign t2_r1_c7_rr2 = t1_r1_c7_rr4 + t1_r1_c7_rr5;
  assign t2_r1_c7_rr3 = t1_r1_c7_rr6 + t1_r1_c7_rr7;

  assign t3_r1_c7_rr0 = t2_r1_c7_rr0 + t2_r1_c7_rr1;
  assign t3_r1_c7_rr1 = t2_r1_c7_rr2 + t2_r1_c7_rr3;

  assign t4_r1_c7_rr0 = t3_r1_c7_rr0 + t3_r1_c7_rr1;

  assign c_1_7 = t4_r1_c7_rr0;
  assign t0_r1_c8_rr0 = a_1_0 * b_0_8;
  assign t0_r1_c8_rr1 = a_1_1 * b_1_8;
  assign t0_r1_c8_rr2 = a_1_2 * b_2_8;
  assign t0_r1_c8_rr3 = a_1_3 * b_3_8;
  assign t0_r1_c8_rr4 = a_1_4 * b_4_8;
  assign t0_r1_c8_rr5 = a_1_5 * b_5_8;
  assign t0_r1_c8_rr6 = a_1_6 * b_6_8;
  assign t0_r1_c8_rr7 = a_1_7 * b_7_8;
  assign t0_r1_c8_rr8 = a_1_8 * b_8_8;
  assign t0_r1_c8_rr9 = a_1_9 * b_9_8;
  assign t0_r1_c8_rr10 = a_1_10 * b_10_8;
  assign t0_r1_c8_rr11 = a_1_11 * b_11_8;
  assign t0_r1_c8_rr12 = a_1_12 * b_12_8;
  assign t0_r1_c8_rr13 = a_1_13 * b_13_8;
  assign t0_r1_c8_rr14 = a_1_14 * b_14_8;
  assign t1_r1_c8_rr0 = t0_r1_c8_rr0 + t0_r1_c8_rr1;
  assign t1_r1_c8_rr1 = t0_r1_c8_rr2 + t0_r1_c8_rr3;
  assign t1_r1_c8_rr2 = t0_r1_c8_rr4 + t0_r1_c8_rr5;
  assign t1_r1_c8_rr3 = t0_r1_c8_rr6 + t0_r1_c8_rr7;
  assign t1_r1_c8_rr4 = t0_r1_c8_rr8 + t0_r1_c8_rr9;
  assign t1_r1_c8_rr5 = t0_r1_c8_rr10 + t0_r1_c8_rr11;
  assign t1_r1_c8_rr6 = t0_r1_c8_rr12 + t0_r1_c8_rr13;
  assign t1_r1_c8_rr7 = t0_r1_c8_rr14;

  assign t2_r1_c8_rr0 = t1_r1_c8_rr0 + t1_r1_c8_rr1;
  assign t2_r1_c8_rr1 = t1_r1_c8_rr2 + t1_r1_c8_rr3;
  assign t2_r1_c8_rr2 = t1_r1_c8_rr4 + t1_r1_c8_rr5;
  assign t2_r1_c8_rr3 = t1_r1_c8_rr6 + t1_r1_c8_rr7;

  assign t3_r1_c8_rr0 = t2_r1_c8_rr0 + t2_r1_c8_rr1;
  assign t3_r1_c8_rr1 = t2_r1_c8_rr2 + t2_r1_c8_rr3;

  assign t4_r1_c8_rr0 = t3_r1_c8_rr0 + t3_r1_c8_rr1;

  assign c_1_8 = t4_r1_c8_rr0;
  assign t0_r1_c9_rr0 = a_1_0 * b_0_9;
  assign t0_r1_c9_rr1 = a_1_1 * b_1_9;
  assign t0_r1_c9_rr2 = a_1_2 * b_2_9;
  assign t0_r1_c9_rr3 = a_1_3 * b_3_9;
  assign t0_r1_c9_rr4 = a_1_4 * b_4_9;
  assign t0_r1_c9_rr5 = a_1_5 * b_5_9;
  assign t0_r1_c9_rr6 = a_1_6 * b_6_9;
  assign t0_r1_c9_rr7 = a_1_7 * b_7_9;
  assign t0_r1_c9_rr8 = a_1_8 * b_8_9;
  assign t0_r1_c9_rr9 = a_1_9 * b_9_9;
  assign t0_r1_c9_rr10 = a_1_10 * b_10_9;
  assign t0_r1_c9_rr11 = a_1_11 * b_11_9;
  assign t0_r1_c9_rr12 = a_1_12 * b_12_9;
  assign t0_r1_c9_rr13 = a_1_13 * b_13_9;
  assign t0_r1_c9_rr14 = a_1_14 * b_14_9;
  assign t1_r1_c9_rr0 = t0_r1_c9_rr0 + t0_r1_c9_rr1;
  assign t1_r1_c9_rr1 = t0_r1_c9_rr2 + t0_r1_c9_rr3;
  assign t1_r1_c9_rr2 = t0_r1_c9_rr4 + t0_r1_c9_rr5;
  assign t1_r1_c9_rr3 = t0_r1_c9_rr6 + t0_r1_c9_rr7;
  assign t1_r1_c9_rr4 = t0_r1_c9_rr8 + t0_r1_c9_rr9;
  assign t1_r1_c9_rr5 = t0_r1_c9_rr10 + t0_r1_c9_rr11;
  assign t1_r1_c9_rr6 = t0_r1_c9_rr12 + t0_r1_c9_rr13;
  assign t1_r1_c9_rr7 = t0_r1_c9_rr14;

  assign t2_r1_c9_rr0 = t1_r1_c9_rr0 + t1_r1_c9_rr1;
  assign t2_r1_c9_rr1 = t1_r1_c9_rr2 + t1_r1_c9_rr3;
  assign t2_r1_c9_rr2 = t1_r1_c9_rr4 + t1_r1_c9_rr5;
  assign t2_r1_c9_rr3 = t1_r1_c9_rr6 + t1_r1_c9_rr7;

  assign t3_r1_c9_rr0 = t2_r1_c9_rr0 + t2_r1_c9_rr1;
  assign t3_r1_c9_rr1 = t2_r1_c9_rr2 + t2_r1_c9_rr3;

  assign t4_r1_c9_rr0 = t3_r1_c9_rr0 + t3_r1_c9_rr1;

  assign c_1_9 = t4_r1_c9_rr0;
  assign t0_r1_c10_rr0 = a_1_0 * b_0_10;
  assign t0_r1_c10_rr1 = a_1_1 * b_1_10;
  assign t0_r1_c10_rr2 = a_1_2 * b_2_10;
  assign t0_r1_c10_rr3 = a_1_3 * b_3_10;
  assign t0_r1_c10_rr4 = a_1_4 * b_4_10;
  assign t0_r1_c10_rr5 = a_1_5 * b_5_10;
  assign t0_r1_c10_rr6 = a_1_6 * b_6_10;
  assign t0_r1_c10_rr7 = a_1_7 * b_7_10;
  assign t0_r1_c10_rr8 = a_1_8 * b_8_10;
  assign t0_r1_c10_rr9 = a_1_9 * b_9_10;
  assign t0_r1_c10_rr10 = a_1_10 * b_10_10;
  assign t0_r1_c10_rr11 = a_1_11 * b_11_10;
  assign t0_r1_c10_rr12 = a_1_12 * b_12_10;
  assign t0_r1_c10_rr13 = a_1_13 * b_13_10;
  assign t0_r1_c10_rr14 = a_1_14 * b_14_10;
  assign t1_r1_c10_rr0 = t0_r1_c10_rr0 + t0_r1_c10_rr1;
  assign t1_r1_c10_rr1 = t0_r1_c10_rr2 + t0_r1_c10_rr3;
  assign t1_r1_c10_rr2 = t0_r1_c10_rr4 + t0_r1_c10_rr5;
  assign t1_r1_c10_rr3 = t0_r1_c10_rr6 + t0_r1_c10_rr7;
  assign t1_r1_c10_rr4 = t0_r1_c10_rr8 + t0_r1_c10_rr9;
  assign t1_r1_c10_rr5 = t0_r1_c10_rr10 + t0_r1_c10_rr11;
  assign t1_r1_c10_rr6 = t0_r1_c10_rr12 + t0_r1_c10_rr13;
  assign t1_r1_c10_rr7 = t0_r1_c10_rr14;

  assign t2_r1_c10_rr0 = t1_r1_c10_rr0 + t1_r1_c10_rr1;
  assign t2_r1_c10_rr1 = t1_r1_c10_rr2 + t1_r1_c10_rr3;
  assign t2_r1_c10_rr2 = t1_r1_c10_rr4 + t1_r1_c10_rr5;
  assign t2_r1_c10_rr3 = t1_r1_c10_rr6 + t1_r1_c10_rr7;

  assign t3_r1_c10_rr0 = t2_r1_c10_rr0 + t2_r1_c10_rr1;
  assign t3_r1_c10_rr1 = t2_r1_c10_rr2 + t2_r1_c10_rr3;

  assign t4_r1_c10_rr0 = t3_r1_c10_rr0 + t3_r1_c10_rr1;

  assign c_1_10 = t4_r1_c10_rr0;
  assign t0_r1_c11_rr0 = a_1_0 * b_0_11;
  assign t0_r1_c11_rr1 = a_1_1 * b_1_11;
  assign t0_r1_c11_rr2 = a_1_2 * b_2_11;
  assign t0_r1_c11_rr3 = a_1_3 * b_3_11;
  assign t0_r1_c11_rr4 = a_1_4 * b_4_11;
  assign t0_r1_c11_rr5 = a_1_5 * b_5_11;
  assign t0_r1_c11_rr6 = a_1_6 * b_6_11;
  assign t0_r1_c11_rr7 = a_1_7 * b_7_11;
  assign t0_r1_c11_rr8 = a_1_8 * b_8_11;
  assign t0_r1_c11_rr9 = a_1_9 * b_9_11;
  assign t0_r1_c11_rr10 = a_1_10 * b_10_11;
  assign t0_r1_c11_rr11 = a_1_11 * b_11_11;
  assign t0_r1_c11_rr12 = a_1_12 * b_12_11;
  assign t0_r1_c11_rr13 = a_1_13 * b_13_11;
  assign t0_r1_c11_rr14 = a_1_14 * b_14_11;
  assign t1_r1_c11_rr0 = t0_r1_c11_rr0 + t0_r1_c11_rr1;
  assign t1_r1_c11_rr1 = t0_r1_c11_rr2 + t0_r1_c11_rr3;
  assign t1_r1_c11_rr2 = t0_r1_c11_rr4 + t0_r1_c11_rr5;
  assign t1_r1_c11_rr3 = t0_r1_c11_rr6 + t0_r1_c11_rr7;
  assign t1_r1_c11_rr4 = t0_r1_c11_rr8 + t0_r1_c11_rr9;
  assign t1_r1_c11_rr5 = t0_r1_c11_rr10 + t0_r1_c11_rr11;
  assign t1_r1_c11_rr6 = t0_r1_c11_rr12 + t0_r1_c11_rr13;
  assign t1_r1_c11_rr7 = t0_r1_c11_rr14;

  assign t2_r1_c11_rr0 = t1_r1_c11_rr0 + t1_r1_c11_rr1;
  assign t2_r1_c11_rr1 = t1_r1_c11_rr2 + t1_r1_c11_rr3;
  assign t2_r1_c11_rr2 = t1_r1_c11_rr4 + t1_r1_c11_rr5;
  assign t2_r1_c11_rr3 = t1_r1_c11_rr6 + t1_r1_c11_rr7;

  assign t3_r1_c11_rr0 = t2_r1_c11_rr0 + t2_r1_c11_rr1;
  assign t3_r1_c11_rr1 = t2_r1_c11_rr2 + t2_r1_c11_rr3;

  assign t4_r1_c11_rr0 = t3_r1_c11_rr0 + t3_r1_c11_rr1;

  assign c_1_11 = t4_r1_c11_rr0;
  assign t0_r1_c12_rr0 = a_1_0 * b_0_12;
  assign t0_r1_c12_rr1 = a_1_1 * b_1_12;
  assign t0_r1_c12_rr2 = a_1_2 * b_2_12;
  assign t0_r1_c12_rr3 = a_1_3 * b_3_12;
  assign t0_r1_c12_rr4 = a_1_4 * b_4_12;
  assign t0_r1_c12_rr5 = a_1_5 * b_5_12;
  assign t0_r1_c12_rr6 = a_1_6 * b_6_12;
  assign t0_r1_c12_rr7 = a_1_7 * b_7_12;
  assign t0_r1_c12_rr8 = a_1_8 * b_8_12;
  assign t0_r1_c12_rr9 = a_1_9 * b_9_12;
  assign t0_r1_c12_rr10 = a_1_10 * b_10_12;
  assign t0_r1_c12_rr11 = a_1_11 * b_11_12;
  assign t0_r1_c12_rr12 = a_1_12 * b_12_12;
  assign t0_r1_c12_rr13 = a_1_13 * b_13_12;
  assign t0_r1_c12_rr14 = a_1_14 * b_14_12;
  assign t1_r1_c12_rr0 = t0_r1_c12_rr0 + t0_r1_c12_rr1;
  assign t1_r1_c12_rr1 = t0_r1_c12_rr2 + t0_r1_c12_rr3;
  assign t1_r1_c12_rr2 = t0_r1_c12_rr4 + t0_r1_c12_rr5;
  assign t1_r1_c12_rr3 = t0_r1_c12_rr6 + t0_r1_c12_rr7;
  assign t1_r1_c12_rr4 = t0_r1_c12_rr8 + t0_r1_c12_rr9;
  assign t1_r1_c12_rr5 = t0_r1_c12_rr10 + t0_r1_c12_rr11;
  assign t1_r1_c12_rr6 = t0_r1_c12_rr12 + t0_r1_c12_rr13;
  assign t1_r1_c12_rr7 = t0_r1_c12_rr14;

  assign t2_r1_c12_rr0 = t1_r1_c12_rr0 + t1_r1_c12_rr1;
  assign t2_r1_c12_rr1 = t1_r1_c12_rr2 + t1_r1_c12_rr3;
  assign t2_r1_c12_rr2 = t1_r1_c12_rr4 + t1_r1_c12_rr5;
  assign t2_r1_c12_rr3 = t1_r1_c12_rr6 + t1_r1_c12_rr7;

  assign t3_r1_c12_rr0 = t2_r1_c12_rr0 + t2_r1_c12_rr1;
  assign t3_r1_c12_rr1 = t2_r1_c12_rr2 + t2_r1_c12_rr3;

  assign t4_r1_c12_rr0 = t3_r1_c12_rr0 + t3_r1_c12_rr1;

  assign c_1_12 = t4_r1_c12_rr0;
  assign t0_r1_c13_rr0 = a_1_0 * b_0_13;
  assign t0_r1_c13_rr1 = a_1_1 * b_1_13;
  assign t0_r1_c13_rr2 = a_1_2 * b_2_13;
  assign t0_r1_c13_rr3 = a_1_3 * b_3_13;
  assign t0_r1_c13_rr4 = a_1_4 * b_4_13;
  assign t0_r1_c13_rr5 = a_1_5 * b_5_13;
  assign t0_r1_c13_rr6 = a_1_6 * b_6_13;
  assign t0_r1_c13_rr7 = a_1_7 * b_7_13;
  assign t0_r1_c13_rr8 = a_1_8 * b_8_13;
  assign t0_r1_c13_rr9 = a_1_9 * b_9_13;
  assign t0_r1_c13_rr10 = a_1_10 * b_10_13;
  assign t0_r1_c13_rr11 = a_1_11 * b_11_13;
  assign t0_r1_c13_rr12 = a_1_12 * b_12_13;
  assign t0_r1_c13_rr13 = a_1_13 * b_13_13;
  assign t0_r1_c13_rr14 = a_1_14 * b_14_13;
  assign t1_r1_c13_rr0 = t0_r1_c13_rr0 + t0_r1_c13_rr1;
  assign t1_r1_c13_rr1 = t0_r1_c13_rr2 + t0_r1_c13_rr3;
  assign t1_r1_c13_rr2 = t0_r1_c13_rr4 + t0_r1_c13_rr5;
  assign t1_r1_c13_rr3 = t0_r1_c13_rr6 + t0_r1_c13_rr7;
  assign t1_r1_c13_rr4 = t0_r1_c13_rr8 + t0_r1_c13_rr9;
  assign t1_r1_c13_rr5 = t0_r1_c13_rr10 + t0_r1_c13_rr11;
  assign t1_r1_c13_rr6 = t0_r1_c13_rr12 + t0_r1_c13_rr13;
  assign t1_r1_c13_rr7 = t0_r1_c13_rr14;

  assign t2_r1_c13_rr0 = t1_r1_c13_rr0 + t1_r1_c13_rr1;
  assign t2_r1_c13_rr1 = t1_r1_c13_rr2 + t1_r1_c13_rr3;
  assign t2_r1_c13_rr2 = t1_r1_c13_rr4 + t1_r1_c13_rr5;
  assign t2_r1_c13_rr3 = t1_r1_c13_rr6 + t1_r1_c13_rr7;

  assign t3_r1_c13_rr0 = t2_r1_c13_rr0 + t2_r1_c13_rr1;
  assign t3_r1_c13_rr1 = t2_r1_c13_rr2 + t2_r1_c13_rr3;

  assign t4_r1_c13_rr0 = t3_r1_c13_rr0 + t3_r1_c13_rr1;

  assign c_1_13 = t4_r1_c13_rr0;
  assign t0_r1_c14_rr0 = a_1_0 * b_0_14;
  assign t0_r1_c14_rr1 = a_1_1 * b_1_14;
  assign t0_r1_c14_rr2 = a_1_2 * b_2_14;
  assign t0_r1_c14_rr3 = a_1_3 * b_3_14;
  assign t0_r1_c14_rr4 = a_1_4 * b_4_14;
  assign t0_r1_c14_rr5 = a_1_5 * b_5_14;
  assign t0_r1_c14_rr6 = a_1_6 * b_6_14;
  assign t0_r1_c14_rr7 = a_1_7 * b_7_14;
  assign t0_r1_c14_rr8 = a_1_8 * b_8_14;
  assign t0_r1_c14_rr9 = a_1_9 * b_9_14;
  assign t0_r1_c14_rr10 = a_1_10 * b_10_14;
  assign t0_r1_c14_rr11 = a_1_11 * b_11_14;
  assign t0_r1_c14_rr12 = a_1_12 * b_12_14;
  assign t0_r1_c14_rr13 = a_1_13 * b_13_14;
  assign t0_r1_c14_rr14 = a_1_14 * b_14_14;
  assign t1_r1_c14_rr0 = t0_r1_c14_rr0 + t0_r1_c14_rr1;
  assign t1_r1_c14_rr1 = t0_r1_c14_rr2 + t0_r1_c14_rr3;
  assign t1_r1_c14_rr2 = t0_r1_c14_rr4 + t0_r1_c14_rr5;
  assign t1_r1_c14_rr3 = t0_r1_c14_rr6 + t0_r1_c14_rr7;
  assign t1_r1_c14_rr4 = t0_r1_c14_rr8 + t0_r1_c14_rr9;
  assign t1_r1_c14_rr5 = t0_r1_c14_rr10 + t0_r1_c14_rr11;
  assign t1_r1_c14_rr6 = t0_r1_c14_rr12 + t0_r1_c14_rr13;
  assign t1_r1_c14_rr7 = t0_r1_c14_rr14;

  assign t2_r1_c14_rr0 = t1_r1_c14_rr0 + t1_r1_c14_rr1;
  assign t2_r1_c14_rr1 = t1_r1_c14_rr2 + t1_r1_c14_rr3;
  assign t2_r1_c14_rr2 = t1_r1_c14_rr4 + t1_r1_c14_rr5;
  assign t2_r1_c14_rr3 = t1_r1_c14_rr6 + t1_r1_c14_rr7;

  assign t3_r1_c14_rr0 = t2_r1_c14_rr0 + t2_r1_c14_rr1;
  assign t3_r1_c14_rr1 = t2_r1_c14_rr2 + t2_r1_c14_rr3;

  assign t4_r1_c14_rr0 = t3_r1_c14_rr0 + t3_r1_c14_rr1;

  assign c_1_14 = t4_r1_c14_rr0;
  assign t0_r2_c0_rr0 = a_2_0 * b_0_0;
  assign t0_r2_c0_rr1 = a_2_1 * b_1_0;
  assign t0_r2_c0_rr2 = a_2_2 * b_2_0;
  assign t0_r2_c0_rr3 = a_2_3 * b_3_0;
  assign t0_r2_c0_rr4 = a_2_4 * b_4_0;
  assign t0_r2_c0_rr5 = a_2_5 * b_5_0;
  assign t0_r2_c0_rr6 = a_2_6 * b_6_0;
  assign t0_r2_c0_rr7 = a_2_7 * b_7_0;
  assign t0_r2_c0_rr8 = a_2_8 * b_8_0;
  assign t0_r2_c0_rr9 = a_2_9 * b_9_0;
  assign t0_r2_c0_rr10 = a_2_10 * b_10_0;
  assign t0_r2_c0_rr11 = a_2_11 * b_11_0;
  assign t0_r2_c0_rr12 = a_2_12 * b_12_0;
  assign t0_r2_c0_rr13 = a_2_13 * b_13_0;
  assign t0_r2_c0_rr14 = a_2_14 * b_14_0;
  assign t1_r2_c0_rr0 = t0_r2_c0_rr0 + t0_r2_c0_rr1;
  assign t1_r2_c0_rr1 = t0_r2_c0_rr2 + t0_r2_c0_rr3;
  assign t1_r2_c0_rr2 = t0_r2_c0_rr4 + t0_r2_c0_rr5;
  assign t1_r2_c0_rr3 = t0_r2_c0_rr6 + t0_r2_c0_rr7;
  assign t1_r2_c0_rr4 = t0_r2_c0_rr8 + t0_r2_c0_rr9;
  assign t1_r2_c0_rr5 = t0_r2_c0_rr10 + t0_r2_c0_rr11;
  assign t1_r2_c0_rr6 = t0_r2_c0_rr12 + t0_r2_c0_rr13;
  assign t1_r2_c0_rr7 = t0_r2_c0_rr14;

  assign t2_r2_c0_rr0 = t1_r2_c0_rr0 + t1_r2_c0_rr1;
  assign t2_r2_c0_rr1 = t1_r2_c0_rr2 + t1_r2_c0_rr3;
  assign t2_r2_c0_rr2 = t1_r2_c0_rr4 + t1_r2_c0_rr5;
  assign t2_r2_c0_rr3 = t1_r2_c0_rr6 + t1_r2_c0_rr7;

  assign t3_r2_c0_rr0 = t2_r2_c0_rr0 + t2_r2_c0_rr1;
  assign t3_r2_c0_rr1 = t2_r2_c0_rr2 + t2_r2_c0_rr3;

  assign t4_r2_c0_rr0 = t3_r2_c0_rr0 + t3_r2_c0_rr1;

  assign c_2_0 = t4_r2_c0_rr0;
  assign t0_r2_c1_rr0 = a_2_0 * b_0_1;
  assign t0_r2_c1_rr1 = a_2_1 * b_1_1;
  assign t0_r2_c1_rr2 = a_2_2 * b_2_1;
  assign t0_r2_c1_rr3 = a_2_3 * b_3_1;
  assign t0_r2_c1_rr4 = a_2_4 * b_4_1;
  assign t0_r2_c1_rr5 = a_2_5 * b_5_1;
  assign t0_r2_c1_rr6 = a_2_6 * b_6_1;
  assign t0_r2_c1_rr7 = a_2_7 * b_7_1;
  assign t0_r2_c1_rr8 = a_2_8 * b_8_1;
  assign t0_r2_c1_rr9 = a_2_9 * b_9_1;
  assign t0_r2_c1_rr10 = a_2_10 * b_10_1;
  assign t0_r2_c1_rr11 = a_2_11 * b_11_1;
  assign t0_r2_c1_rr12 = a_2_12 * b_12_1;
  assign t0_r2_c1_rr13 = a_2_13 * b_13_1;
  assign t0_r2_c1_rr14 = a_2_14 * b_14_1;
  assign t1_r2_c1_rr0 = t0_r2_c1_rr0 + t0_r2_c1_rr1;
  assign t1_r2_c1_rr1 = t0_r2_c1_rr2 + t0_r2_c1_rr3;
  assign t1_r2_c1_rr2 = t0_r2_c1_rr4 + t0_r2_c1_rr5;
  assign t1_r2_c1_rr3 = t0_r2_c1_rr6 + t0_r2_c1_rr7;
  assign t1_r2_c1_rr4 = t0_r2_c1_rr8 + t0_r2_c1_rr9;
  assign t1_r2_c1_rr5 = t0_r2_c1_rr10 + t0_r2_c1_rr11;
  assign t1_r2_c1_rr6 = t0_r2_c1_rr12 + t0_r2_c1_rr13;
  assign t1_r2_c1_rr7 = t0_r2_c1_rr14;

  assign t2_r2_c1_rr0 = t1_r2_c1_rr0 + t1_r2_c1_rr1;
  assign t2_r2_c1_rr1 = t1_r2_c1_rr2 + t1_r2_c1_rr3;
  assign t2_r2_c1_rr2 = t1_r2_c1_rr4 + t1_r2_c1_rr5;
  assign t2_r2_c1_rr3 = t1_r2_c1_rr6 + t1_r2_c1_rr7;

  assign t3_r2_c1_rr0 = t2_r2_c1_rr0 + t2_r2_c1_rr1;
  assign t3_r2_c1_rr1 = t2_r2_c1_rr2 + t2_r2_c1_rr3;

  assign t4_r2_c1_rr0 = t3_r2_c1_rr0 + t3_r2_c1_rr1;

  assign c_2_1 = t4_r2_c1_rr0;
  assign t0_r2_c2_rr0 = a_2_0 * b_0_2;
  assign t0_r2_c2_rr1 = a_2_1 * b_1_2;
  assign t0_r2_c2_rr2 = a_2_2 * b_2_2;
  assign t0_r2_c2_rr3 = a_2_3 * b_3_2;
  assign t0_r2_c2_rr4 = a_2_4 * b_4_2;
  assign t0_r2_c2_rr5 = a_2_5 * b_5_2;
  assign t0_r2_c2_rr6 = a_2_6 * b_6_2;
  assign t0_r2_c2_rr7 = a_2_7 * b_7_2;
  assign t0_r2_c2_rr8 = a_2_8 * b_8_2;
  assign t0_r2_c2_rr9 = a_2_9 * b_9_2;
  assign t0_r2_c2_rr10 = a_2_10 * b_10_2;
  assign t0_r2_c2_rr11 = a_2_11 * b_11_2;
  assign t0_r2_c2_rr12 = a_2_12 * b_12_2;
  assign t0_r2_c2_rr13 = a_2_13 * b_13_2;
  assign t0_r2_c2_rr14 = a_2_14 * b_14_2;
  assign t1_r2_c2_rr0 = t0_r2_c2_rr0 + t0_r2_c2_rr1;
  assign t1_r2_c2_rr1 = t0_r2_c2_rr2 + t0_r2_c2_rr3;
  assign t1_r2_c2_rr2 = t0_r2_c2_rr4 + t0_r2_c2_rr5;
  assign t1_r2_c2_rr3 = t0_r2_c2_rr6 + t0_r2_c2_rr7;
  assign t1_r2_c2_rr4 = t0_r2_c2_rr8 + t0_r2_c2_rr9;
  assign t1_r2_c2_rr5 = t0_r2_c2_rr10 + t0_r2_c2_rr11;
  assign t1_r2_c2_rr6 = t0_r2_c2_rr12 + t0_r2_c2_rr13;
  assign t1_r2_c2_rr7 = t0_r2_c2_rr14;

  assign t2_r2_c2_rr0 = t1_r2_c2_rr0 + t1_r2_c2_rr1;
  assign t2_r2_c2_rr1 = t1_r2_c2_rr2 + t1_r2_c2_rr3;
  assign t2_r2_c2_rr2 = t1_r2_c2_rr4 + t1_r2_c2_rr5;
  assign t2_r2_c2_rr3 = t1_r2_c2_rr6 + t1_r2_c2_rr7;

  assign t3_r2_c2_rr0 = t2_r2_c2_rr0 + t2_r2_c2_rr1;
  assign t3_r2_c2_rr1 = t2_r2_c2_rr2 + t2_r2_c2_rr3;

  assign t4_r2_c2_rr0 = t3_r2_c2_rr0 + t3_r2_c2_rr1;

  assign c_2_2 = t4_r2_c2_rr0;
  assign t0_r2_c3_rr0 = a_2_0 * b_0_3;
  assign t0_r2_c3_rr1 = a_2_1 * b_1_3;
  assign t0_r2_c3_rr2 = a_2_2 * b_2_3;
  assign t0_r2_c3_rr3 = a_2_3 * b_3_3;
  assign t0_r2_c3_rr4 = a_2_4 * b_4_3;
  assign t0_r2_c3_rr5 = a_2_5 * b_5_3;
  assign t0_r2_c3_rr6 = a_2_6 * b_6_3;
  assign t0_r2_c3_rr7 = a_2_7 * b_7_3;
  assign t0_r2_c3_rr8 = a_2_8 * b_8_3;
  assign t0_r2_c3_rr9 = a_2_9 * b_9_3;
  assign t0_r2_c3_rr10 = a_2_10 * b_10_3;
  assign t0_r2_c3_rr11 = a_2_11 * b_11_3;
  assign t0_r2_c3_rr12 = a_2_12 * b_12_3;
  assign t0_r2_c3_rr13 = a_2_13 * b_13_3;
  assign t0_r2_c3_rr14 = a_2_14 * b_14_3;
  assign t1_r2_c3_rr0 = t0_r2_c3_rr0 + t0_r2_c3_rr1;
  assign t1_r2_c3_rr1 = t0_r2_c3_rr2 + t0_r2_c3_rr3;
  assign t1_r2_c3_rr2 = t0_r2_c3_rr4 + t0_r2_c3_rr5;
  assign t1_r2_c3_rr3 = t0_r2_c3_rr6 + t0_r2_c3_rr7;
  assign t1_r2_c3_rr4 = t0_r2_c3_rr8 + t0_r2_c3_rr9;
  assign t1_r2_c3_rr5 = t0_r2_c3_rr10 + t0_r2_c3_rr11;
  assign t1_r2_c3_rr6 = t0_r2_c3_rr12 + t0_r2_c3_rr13;
  assign t1_r2_c3_rr7 = t0_r2_c3_rr14;

  assign t2_r2_c3_rr0 = t1_r2_c3_rr0 + t1_r2_c3_rr1;
  assign t2_r2_c3_rr1 = t1_r2_c3_rr2 + t1_r2_c3_rr3;
  assign t2_r2_c3_rr2 = t1_r2_c3_rr4 + t1_r2_c3_rr5;
  assign t2_r2_c3_rr3 = t1_r2_c3_rr6 + t1_r2_c3_rr7;

  assign t3_r2_c3_rr0 = t2_r2_c3_rr0 + t2_r2_c3_rr1;
  assign t3_r2_c3_rr1 = t2_r2_c3_rr2 + t2_r2_c3_rr3;

  assign t4_r2_c3_rr0 = t3_r2_c3_rr0 + t3_r2_c3_rr1;

  assign c_2_3 = t4_r2_c3_rr0;
  assign t0_r2_c4_rr0 = a_2_0 * b_0_4;
  assign t0_r2_c4_rr1 = a_2_1 * b_1_4;
  assign t0_r2_c4_rr2 = a_2_2 * b_2_4;
  assign t0_r2_c4_rr3 = a_2_3 * b_3_4;
  assign t0_r2_c4_rr4 = a_2_4 * b_4_4;
  assign t0_r2_c4_rr5 = a_2_5 * b_5_4;
  assign t0_r2_c4_rr6 = a_2_6 * b_6_4;
  assign t0_r2_c4_rr7 = a_2_7 * b_7_4;
  assign t0_r2_c4_rr8 = a_2_8 * b_8_4;
  assign t0_r2_c4_rr9 = a_2_9 * b_9_4;
  assign t0_r2_c4_rr10 = a_2_10 * b_10_4;
  assign t0_r2_c4_rr11 = a_2_11 * b_11_4;
  assign t0_r2_c4_rr12 = a_2_12 * b_12_4;
  assign t0_r2_c4_rr13 = a_2_13 * b_13_4;
  assign t0_r2_c4_rr14 = a_2_14 * b_14_4;
  assign t1_r2_c4_rr0 = t0_r2_c4_rr0 + t0_r2_c4_rr1;
  assign t1_r2_c4_rr1 = t0_r2_c4_rr2 + t0_r2_c4_rr3;
  assign t1_r2_c4_rr2 = t0_r2_c4_rr4 + t0_r2_c4_rr5;
  assign t1_r2_c4_rr3 = t0_r2_c4_rr6 + t0_r2_c4_rr7;
  assign t1_r2_c4_rr4 = t0_r2_c4_rr8 + t0_r2_c4_rr9;
  assign t1_r2_c4_rr5 = t0_r2_c4_rr10 + t0_r2_c4_rr11;
  assign t1_r2_c4_rr6 = t0_r2_c4_rr12 + t0_r2_c4_rr13;
  assign t1_r2_c4_rr7 = t0_r2_c4_rr14;

  assign t2_r2_c4_rr0 = t1_r2_c4_rr0 + t1_r2_c4_rr1;
  assign t2_r2_c4_rr1 = t1_r2_c4_rr2 + t1_r2_c4_rr3;
  assign t2_r2_c4_rr2 = t1_r2_c4_rr4 + t1_r2_c4_rr5;
  assign t2_r2_c4_rr3 = t1_r2_c4_rr6 + t1_r2_c4_rr7;

  assign t3_r2_c4_rr0 = t2_r2_c4_rr0 + t2_r2_c4_rr1;
  assign t3_r2_c4_rr1 = t2_r2_c4_rr2 + t2_r2_c4_rr3;

  assign t4_r2_c4_rr0 = t3_r2_c4_rr0 + t3_r2_c4_rr1;

  assign c_2_4 = t4_r2_c4_rr0;
  assign t0_r2_c5_rr0 = a_2_0 * b_0_5;
  assign t0_r2_c5_rr1 = a_2_1 * b_1_5;
  assign t0_r2_c5_rr2 = a_2_2 * b_2_5;
  assign t0_r2_c5_rr3 = a_2_3 * b_3_5;
  assign t0_r2_c5_rr4 = a_2_4 * b_4_5;
  assign t0_r2_c5_rr5 = a_2_5 * b_5_5;
  assign t0_r2_c5_rr6 = a_2_6 * b_6_5;
  assign t0_r2_c5_rr7 = a_2_7 * b_7_5;
  assign t0_r2_c5_rr8 = a_2_8 * b_8_5;
  assign t0_r2_c5_rr9 = a_2_9 * b_9_5;
  assign t0_r2_c5_rr10 = a_2_10 * b_10_5;
  assign t0_r2_c5_rr11 = a_2_11 * b_11_5;
  assign t0_r2_c5_rr12 = a_2_12 * b_12_5;
  assign t0_r2_c5_rr13 = a_2_13 * b_13_5;
  assign t0_r2_c5_rr14 = a_2_14 * b_14_5;
  assign t1_r2_c5_rr0 = t0_r2_c5_rr0 + t0_r2_c5_rr1;
  assign t1_r2_c5_rr1 = t0_r2_c5_rr2 + t0_r2_c5_rr3;
  assign t1_r2_c5_rr2 = t0_r2_c5_rr4 + t0_r2_c5_rr5;
  assign t1_r2_c5_rr3 = t0_r2_c5_rr6 + t0_r2_c5_rr7;
  assign t1_r2_c5_rr4 = t0_r2_c5_rr8 + t0_r2_c5_rr9;
  assign t1_r2_c5_rr5 = t0_r2_c5_rr10 + t0_r2_c5_rr11;
  assign t1_r2_c5_rr6 = t0_r2_c5_rr12 + t0_r2_c5_rr13;
  assign t1_r2_c5_rr7 = t0_r2_c5_rr14;

  assign t2_r2_c5_rr0 = t1_r2_c5_rr0 + t1_r2_c5_rr1;
  assign t2_r2_c5_rr1 = t1_r2_c5_rr2 + t1_r2_c5_rr3;
  assign t2_r2_c5_rr2 = t1_r2_c5_rr4 + t1_r2_c5_rr5;
  assign t2_r2_c5_rr3 = t1_r2_c5_rr6 + t1_r2_c5_rr7;

  assign t3_r2_c5_rr0 = t2_r2_c5_rr0 + t2_r2_c5_rr1;
  assign t3_r2_c5_rr1 = t2_r2_c5_rr2 + t2_r2_c5_rr3;

  assign t4_r2_c5_rr0 = t3_r2_c5_rr0 + t3_r2_c5_rr1;

  assign c_2_5 = t4_r2_c5_rr0;
  assign t0_r2_c6_rr0 = a_2_0 * b_0_6;
  assign t0_r2_c6_rr1 = a_2_1 * b_1_6;
  assign t0_r2_c6_rr2 = a_2_2 * b_2_6;
  assign t0_r2_c6_rr3 = a_2_3 * b_3_6;
  assign t0_r2_c6_rr4 = a_2_4 * b_4_6;
  assign t0_r2_c6_rr5 = a_2_5 * b_5_6;
  assign t0_r2_c6_rr6 = a_2_6 * b_6_6;
  assign t0_r2_c6_rr7 = a_2_7 * b_7_6;
  assign t0_r2_c6_rr8 = a_2_8 * b_8_6;
  assign t0_r2_c6_rr9 = a_2_9 * b_9_6;
  assign t0_r2_c6_rr10 = a_2_10 * b_10_6;
  assign t0_r2_c6_rr11 = a_2_11 * b_11_6;
  assign t0_r2_c6_rr12 = a_2_12 * b_12_6;
  assign t0_r2_c6_rr13 = a_2_13 * b_13_6;
  assign t0_r2_c6_rr14 = a_2_14 * b_14_6;
  assign t1_r2_c6_rr0 = t0_r2_c6_rr0 + t0_r2_c6_rr1;
  assign t1_r2_c6_rr1 = t0_r2_c6_rr2 + t0_r2_c6_rr3;
  assign t1_r2_c6_rr2 = t0_r2_c6_rr4 + t0_r2_c6_rr5;
  assign t1_r2_c6_rr3 = t0_r2_c6_rr6 + t0_r2_c6_rr7;
  assign t1_r2_c6_rr4 = t0_r2_c6_rr8 + t0_r2_c6_rr9;
  assign t1_r2_c6_rr5 = t0_r2_c6_rr10 + t0_r2_c6_rr11;
  assign t1_r2_c6_rr6 = t0_r2_c6_rr12 + t0_r2_c6_rr13;
  assign t1_r2_c6_rr7 = t0_r2_c6_rr14;

  assign t2_r2_c6_rr0 = t1_r2_c6_rr0 + t1_r2_c6_rr1;
  assign t2_r2_c6_rr1 = t1_r2_c6_rr2 + t1_r2_c6_rr3;
  assign t2_r2_c6_rr2 = t1_r2_c6_rr4 + t1_r2_c6_rr5;
  assign t2_r2_c6_rr3 = t1_r2_c6_rr6 + t1_r2_c6_rr7;

  assign t3_r2_c6_rr0 = t2_r2_c6_rr0 + t2_r2_c6_rr1;
  assign t3_r2_c6_rr1 = t2_r2_c6_rr2 + t2_r2_c6_rr3;

  assign t4_r2_c6_rr0 = t3_r2_c6_rr0 + t3_r2_c6_rr1;

  assign c_2_6 = t4_r2_c6_rr0;
  assign t0_r2_c7_rr0 = a_2_0 * b_0_7;
  assign t0_r2_c7_rr1 = a_2_1 * b_1_7;
  assign t0_r2_c7_rr2 = a_2_2 * b_2_7;
  assign t0_r2_c7_rr3 = a_2_3 * b_3_7;
  assign t0_r2_c7_rr4 = a_2_4 * b_4_7;
  assign t0_r2_c7_rr5 = a_2_5 * b_5_7;
  assign t0_r2_c7_rr6 = a_2_6 * b_6_7;
  assign t0_r2_c7_rr7 = a_2_7 * b_7_7;
  assign t0_r2_c7_rr8 = a_2_8 * b_8_7;
  assign t0_r2_c7_rr9 = a_2_9 * b_9_7;
  assign t0_r2_c7_rr10 = a_2_10 * b_10_7;
  assign t0_r2_c7_rr11 = a_2_11 * b_11_7;
  assign t0_r2_c7_rr12 = a_2_12 * b_12_7;
  assign t0_r2_c7_rr13 = a_2_13 * b_13_7;
  assign t0_r2_c7_rr14 = a_2_14 * b_14_7;
  assign t1_r2_c7_rr0 = t0_r2_c7_rr0 + t0_r2_c7_rr1;
  assign t1_r2_c7_rr1 = t0_r2_c7_rr2 + t0_r2_c7_rr3;
  assign t1_r2_c7_rr2 = t0_r2_c7_rr4 + t0_r2_c7_rr5;
  assign t1_r2_c7_rr3 = t0_r2_c7_rr6 + t0_r2_c7_rr7;
  assign t1_r2_c7_rr4 = t0_r2_c7_rr8 + t0_r2_c7_rr9;
  assign t1_r2_c7_rr5 = t0_r2_c7_rr10 + t0_r2_c7_rr11;
  assign t1_r2_c7_rr6 = t0_r2_c7_rr12 + t0_r2_c7_rr13;
  assign t1_r2_c7_rr7 = t0_r2_c7_rr14;

  assign t2_r2_c7_rr0 = t1_r2_c7_rr0 + t1_r2_c7_rr1;
  assign t2_r2_c7_rr1 = t1_r2_c7_rr2 + t1_r2_c7_rr3;
  assign t2_r2_c7_rr2 = t1_r2_c7_rr4 + t1_r2_c7_rr5;
  assign t2_r2_c7_rr3 = t1_r2_c7_rr6 + t1_r2_c7_rr7;

  assign t3_r2_c7_rr0 = t2_r2_c7_rr0 + t2_r2_c7_rr1;
  assign t3_r2_c7_rr1 = t2_r2_c7_rr2 + t2_r2_c7_rr3;

  assign t4_r2_c7_rr0 = t3_r2_c7_rr0 + t3_r2_c7_rr1;

  assign c_2_7 = t4_r2_c7_rr0;
  assign t0_r2_c8_rr0 = a_2_0 * b_0_8;
  assign t0_r2_c8_rr1 = a_2_1 * b_1_8;
  assign t0_r2_c8_rr2 = a_2_2 * b_2_8;
  assign t0_r2_c8_rr3 = a_2_3 * b_3_8;
  assign t0_r2_c8_rr4 = a_2_4 * b_4_8;
  assign t0_r2_c8_rr5 = a_2_5 * b_5_8;
  assign t0_r2_c8_rr6 = a_2_6 * b_6_8;
  assign t0_r2_c8_rr7 = a_2_7 * b_7_8;
  assign t0_r2_c8_rr8 = a_2_8 * b_8_8;
  assign t0_r2_c8_rr9 = a_2_9 * b_9_8;
  assign t0_r2_c8_rr10 = a_2_10 * b_10_8;
  assign t0_r2_c8_rr11 = a_2_11 * b_11_8;
  assign t0_r2_c8_rr12 = a_2_12 * b_12_8;
  assign t0_r2_c8_rr13 = a_2_13 * b_13_8;
  assign t0_r2_c8_rr14 = a_2_14 * b_14_8;
  assign t1_r2_c8_rr0 = t0_r2_c8_rr0 + t0_r2_c8_rr1;
  assign t1_r2_c8_rr1 = t0_r2_c8_rr2 + t0_r2_c8_rr3;
  assign t1_r2_c8_rr2 = t0_r2_c8_rr4 + t0_r2_c8_rr5;
  assign t1_r2_c8_rr3 = t0_r2_c8_rr6 + t0_r2_c8_rr7;
  assign t1_r2_c8_rr4 = t0_r2_c8_rr8 + t0_r2_c8_rr9;
  assign t1_r2_c8_rr5 = t0_r2_c8_rr10 + t0_r2_c8_rr11;
  assign t1_r2_c8_rr6 = t0_r2_c8_rr12 + t0_r2_c8_rr13;
  assign t1_r2_c8_rr7 = t0_r2_c8_rr14;

  assign t2_r2_c8_rr0 = t1_r2_c8_rr0 + t1_r2_c8_rr1;
  assign t2_r2_c8_rr1 = t1_r2_c8_rr2 + t1_r2_c8_rr3;
  assign t2_r2_c8_rr2 = t1_r2_c8_rr4 + t1_r2_c8_rr5;
  assign t2_r2_c8_rr3 = t1_r2_c8_rr6 + t1_r2_c8_rr7;

  assign t3_r2_c8_rr0 = t2_r2_c8_rr0 + t2_r2_c8_rr1;
  assign t3_r2_c8_rr1 = t2_r2_c8_rr2 + t2_r2_c8_rr3;

  assign t4_r2_c8_rr0 = t3_r2_c8_rr0 + t3_r2_c8_rr1;

  assign c_2_8 = t4_r2_c8_rr0;
  assign t0_r2_c9_rr0 = a_2_0 * b_0_9;
  assign t0_r2_c9_rr1 = a_2_1 * b_1_9;
  assign t0_r2_c9_rr2 = a_2_2 * b_2_9;
  assign t0_r2_c9_rr3 = a_2_3 * b_3_9;
  assign t0_r2_c9_rr4 = a_2_4 * b_4_9;
  assign t0_r2_c9_rr5 = a_2_5 * b_5_9;
  assign t0_r2_c9_rr6 = a_2_6 * b_6_9;
  assign t0_r2_c9_rr7 = a_2_7 * b_7_9;
  assign t0_r2_c9_rr8 = a_2_8 * b_8_9;
  assign t0_r2_c9_rr9 = a_2_9 * b_9_9;
  assign t0_r2_c9_rr10 = a_2_10 * b_10_9;
  assign t0_r2_c9_rr11 = a_2_11 * b_11_9;
  assign t0_r2_c9_rr12 = a_2_12 * b_12_9;
  assign t0_r2_c9_rr13 = a_2_13 * b_13_9;
  assign t0_r2_c9_rr14 = a_2_14 * b_14_9;
  assign t1_r2_c9_rr0 = t0_r2_c9_rr0 + t0_r2_c9_rr1;
  assign t1_r2_c9_rr1 = t0_r2_c9_rr2 + t0_r2_c9_rr3;
  assign t1_r2_c9_rr2 = t0_r2_c9_rr4 + t0_r2_c9_rr5;
  assign t1_r2_c9_rr3 = t0_r2_c9_rr6 + t0_r2_c9_rr7;
  assign t1_r2_c9_rr4 = t0_r2_c9_rr8 + t0_r2_c9_rr9;
  assign t1_r2_c9_rr5 = t0_r2_c9_rr10 + t0_r2_c9_rr11;
  assign t1_r2_c9_rr6 = t0_r2_c9_rr12 + t0_r2_c9_rr13;
  assign t1_r2_c9_rr7 = t0_r2_c9_rr14;

  assign t2_r2_c9_rr0 = t1_r2_c9_rr0 + t1_r2_c9_rr1;
  assign t2_r2_c9_rr1 = t1_r2_c9_rr2 + t1_r2_c9_rr3;
  assign t2_r2_c9_rr2 = t1_r2_c9_rr4 + t1_r2_c9_rr5;
  assign t2_r2_c9_rr3 = t1_r2_c9_rr6 + t1_r2_c9_rr7;

  assign t3_r2_c9_rr0 = t2_r2_c9_rr0 + t2_r2_c9_rr1;
  assign t3_r2_c9_rr1 = t2_r2_c9_rr2 + t2_r2_c9_rr3;

  assign t4_r2_c9_rr0 = t3_r2_c9_rr0 + t3_r2_c9_rr1;

  assign c_2_9 = t4_r2_c9_rr0;
  assign t0_r2_c10_rr0 = a_2_0 * b_0_10;
  assign t0_r2_c10_rr1 = a_2_1 * b_1_10;
  assign t0_r2_c10_rr2 = a_2_2 * b_2_10;
  assign t0_r2_c10_rr3 = a_2_3 * b_3_10;
  assign t0_r2_c10_rr4 = a_2_4 * b_4_10;
  assign t0_r2_c10_rr5 = a_2_5 * b_5_10;
  assign t0_r2_c10_rr6 = a_2_6 * b_6_10;
  assign t0_r2_c10_rr7 = a_2_7 * b_7_10;
  assign t0_r2_c10_rr8 = a_2_8 * b_8_10;
  assign t0_r2_c10_rr9 = a_2_9 * b_9_10;
  assign t0_r2_c10_rr10 = a_2_10 * b_10_10;
  assign t0_r2_c10_rr11 = a_2_11 * b_11_10;
  assign t0_r2_c10_rr12 = a_2_12 * b_12_10;
  assign t0_r2_c10_rr13 = a_2_13 * b_13_10;
  assign t0_r2_c10_rr14 = a_2_14 * b_14_10;
  assign t1_r2_c10_rr0 = t0_r2_c10_rr0 + t0_r2_c10_rr1;
  assign t1_r2_c10_rr1 = t0_r2_c10_rr2 + t0_r2_c10_rr3;
  assign t1_r2_c10_rr2 = t0_r2_c10_rr4 + t0_r2_c10_rr5;
  assign t1_r2_c10_rr3 = t0_r2_c10_rr6 + t0_r2_c10_rr7;
  assign t1_r2_c10_rr4 = t0_r2_c10_rr8 + t0_r2_c10_rr9;
  assign t1_r2_c10_rr5 = t0_r2_c10_rr10 + t0_r2_c10_rr11;
  assign t1_r2_c10_rr6 = t0_r2_c10_rr12 + t0_r2_c10_rr13;
  assign t1_r2_c10_rr7 = t0_r2_c10_rr14;

  assign t2_r2_c10_rr0 = t1_r2_c10_rr0 + t1_r2_c10_rr1;
  assign t2_r2_c10_rr1 = t1_r2_c10_rr2 + t1_r2_c10_rr3;
  assign t2_r2_c10_rr2 = t1_r2_c10_rr4 + t1_r2_c10_rr5;
  assign t2_r2_c10_rr3 = t1_r2_c10_rr6 + t1_r2_c10_rr7;

  assign t3_r2_c10_rr0 = t2_r2_c10_rr0 + t2_r2_c10_rr1;
  assign t3_r2_c10_rr1 = t2_r2_c10_rr2 + t2_r2_c10_rr3;

  assign t4_r2_c10_rr0 = t3_r2_c10_rr0 + t3_r2_c10_rr1;

  assign c_2_10 = t4_r2_c10_rr0;
  assign t0_r2_c11_rr0 = a_2_0 * b_0_11;
  assign t0_r2_c11_rr1 = a_2_1 * b_1_11;
  assign t0_r2_c11_rr2 = a_2_2 * b_2_11;
  assign t0_r2_c11_rr3 = a_2_3 * b_3_11;
  assign t0_r2_c11_rr4 = a_2_4 * b_4_11;
  assign t0_r2_c11_rr5 = a_2_5 * b_5_11;
  assign t0_r2_c11_rr6 = a_2_6 * b_6_11;
  assign t0_r2_c11_rr7 = a_2_7 * b_7_11;
  assign t0_r2_c11_rr8 = a_2_8 * b_8_11;
  assign t0_r2_c11_rr9 = a_2_9 * b_9_11;
  assign t0_r2_c11_rr10 = a_2_10 * b_10_11;
  assign t0_r2_c11_rr11 = a_2_11 * b_11_11;
  assign t0_r2_c11_rr12 = a_2_12 * b_12_11;
  assign t0_r2_c11_rr13 = a_2_13 * b_13_11;
  assign t0_r2_c11_rr14 = a_2_14 * b_14_11;
  assign t1_r2_c11_rr0 = t0_r2_c11_rr0 + t0_r2_c11_rr1;
  assign t1_r2_c11_rr1 = t0_r2_c11_rr2 + t0_r2_c11_rr3;
  assign t1_r2_c11_rr2 = t0_r2_c11_rr4 + t0_r2_c11_rr5;
  assign t1_r2_c11_rr3 = t0_r2_c11_rr6 + t0_r2_c11_rr7;
  assign t1_r2_c11_rr4 = t0_r2_c11_rr8 + t0_r2_c11_rr9;
  assign t1_r2_c11_rr5 = t0_r2_c11_rr10 + t0_r2_c11_rr11;
  assign t1_r2_c11_rr6 = t0_r2_c11_rr12 + t0_r2_c11_rr13;
  assign t1_r2_c11_rr7 = t0_r2_c11_rr14;

  assign t2_r2_c11_rr0 = t1_r2_c11_rr0 + t1_r2_c11_rr1;
  assign t2_r2_c11_rr1 = t1_r2_c11_rr2 + t1_r2_c11_rr3;
  assign t2_r2_c11_rr2 = t1_r2_c11_rr4 + t1_r2_c11_rr5;
  assign t2_r2_c11_rr3 = t1_r2_c11_rr6 + t1_r2_c11_rr7;

  assign t3_r2_c11_rr0 = t2_r2_c11_rr0 + t2_r2_c11_rr1;
  assign t3_r2_c11_rr1 = t2_r2_c11_rr2 + t2_r2_c11_rr3;

  assign t4_r2_c11_rr0 = t3_r2_c11_rr0 + t3_r2_c11_rr1;

  assign c_2_11 = t4_r2_c11_rr0;
  assign t0_r2_c12_rr0 = a_2_0 * b_0_12;
  assign t0_r2_c12_rr1 = a_2_1 * b_1_12;
  assign t0_r2_c12_rr2 = a_2_2 * b_2_12;
  assign t0_r2_c12_rr3 = a_2_3 * b_3_12;
  assign t0_r2_c12_rr4 = a_2_4 * b_4_12;
  assign t0_r2_c12_rr5 = a_2_5 * b_5_12;
  assign t0_r2_c12_rr6 = a_2_6 * b_6_12;
  assign t0_r2_c12_rr7 = a_2_7 * b_7_12;
  assign t0_r2_c12_rr8 = a_2_8 * b_8_12;
  assign t0_r2_c12_rr9 = a_2_9 * b_9_12;
  assign t0_r2_c12_rr10 = a_2_10 * b_10_12;
  assign t0_r2_c12_rr11 = a_2_11 * b_11_12;
  assign t0_r2_c12_rr12 = a_2_12 * b_12_12;
  assign t0_r2_c12_rr13 = a_2_13 * b_13_12;
  assign t0_r2_c12_rr14 = a_2_14 * b_14_12;
  assign t1_r2_c12_rr0 = t0_r2_c12_rr0 + t0_r2_c12_rr1;
  assign t1_r2_c12_rr1 = t0_r2_c12_rr2 + t0_r2_c12_rr3;
  assign t1_r2_c12_rr2 = t0_r2_c12_rr4 + t0_r2_c12_rr5;
  assign t1_r2_c12_rr3 = t0_r2_c12_rr6 + t0_r2_c12_rr7;
  assign t1_r2_c12_rr4 = t0_r2_c12_rr8 + t0_r2_c12_rr9;
  assign t1_r2_c12_rr5 = t0_r2_c12_rr10 + t0_r2_c12_rr11;
  assign t1_r2_c12_rr6 = t0_r2_c12_rr12 + t0_r2_c12_rr13;
  assign t1_r2_c12_rr7 = t0_r2_c12_rr14;

  assign t2_r2_c12_rr0 = t1_r2_c12_rr0 + t1_r2_c12_rr1;
  assign t2_r2_c12_rr1 = t1_r2_c12_rr2 + t1_r2_c12_rr3;
  assign t2_r2_c12_rr2 = t1_r2_c12_rr4 + t1_r2_c12_rr5;
  assign t2_r2_c12_rr3 = t1_r2_c12_rr6 + t1_r2_c12_rr7;

  assign t3_r2_c12_rr0 = t2_r2_c12_rr0 + t2_r2_c12_rr1;
  assign t3_r2_c12_rr1 = t2_r2_c12_rr2 + t2_r2_c12_rr3;

  assign t4_r2_c12_rr0 = t3_r2_c12_rr0 + t3_r2_c12_rr1;

  assign c_2_12 = t4_r2_c12_rr0;
  assign t0_r2_c13_rr0 = a_2_0 * b_0_13;
  assign t0_r2_c13_rr1 = a_2_1 * b_1_13;
  assign t0_r2_c13_rr2 = a_2_2 * b_2_13;
  assign t0_r2_c13_rr3 = a_2_3 * b_3_13;
  assign t0_r2_c13_rr4 = a_2_4 * b_4_13;
  assign t0_r2_c13_rr5 = a_2_5 * b_5_13;
  assign t0_r2_c13_rr6 = a_2_6 * b_6_13;
  assign t0_r2_c13_rr7 = a_2_7 * b_7_13;
  assign t0_r2_c13_rr8 = a_2_8 * b_8_13;
  assign t0_r2_c13_rr9 = a_2_9 * b_9_13;
  assign t0_r2_c13_rr10 = a_2_10 * b_10_13;
  assign t0_r2_c13_rr11 = a_2_11 * b_11_13;
  assign t0_r2_c13_rr12 = a_2_12 * b_12_13;
  assign t0_r2_c13_rr13 = a_2_13 * b_13_13;
  assign t0_r2_c13_rr14 = a_2_14 * b_14_13;
  assign t1_r2_c13_rr0 = t0_r2_c13_rr0 + t0_r2_c13_rr1;
  assign t1_r2_c13_rr1 = t0_r2_c13_rr2 + t0_r2_c13_rr3;
  assign t1_r2_c13_rr2 = t0_r2_c13_rr4 + t0_r2_c13_rr5;
  assign t1_r2_c13_rr3 = t0_r2_c13_rr6 + t0_r2_c13_rr7;
  assign t1_r2_c13_rr4 = t0_r2_c13_rr8 + t0_r2_c13_rr9;
  assign t1_r2_c13_rr5 = t0_r2_c13_rr10 + t0_r2_c13_rr11;
  assign t1_r2_c13_rr6 = t0_r2_c13_rr12 + t0_r2_c13_rr13;
  assign t1_r2_c13_rr7 = t0_r2_c13_rr14;

  assign t2_r2_c13_rr0 = t1_r2_c13_rr0 + t1_r2_c13_rr1;
  assign t2_r2_c13_rr1 = t1_r2_c13_rr2 + t1_r2_c13_rr3;
  assign t2_r2_c13_rr2 = t1_r2_c13_rr4 + t1_r2_c13_rr5;
  assign t2_r2_c13_rr3 = t1_r2_c13_rr6 + t1_r2_c13_rr7;

  assign t3_r2_c13_rr0 = t2_r2_c13_rr0 + t2_r2_c13_rr1;
  assign t3_r2_c13_rr1 = t2_r2_c13_rr2 + t2_r2_c13_rr3;

  assign t4_r2_c13_rr0 = t3_r2_c13_rr0 + t3_r2_c13_rr1;

  assign c_2_13 = t4_r2_c13_rr0;
  assign t0_r2_c14_rr0 = a_2_0 * b_0_14;
  assign t0_r2_c14_rr1 = a_2_1 * b_1_14;
  assign t0_r2_c14_rr2 = a_2_2 * b_2_14;
  assign t0_r2_c14_rr3 = a_2_3 * b_3_14;
  assign t0_r2_c14_rr4 = a_2_4 * b_4_14;
  assign t0_r2_c14_rr5 = a_2_5 * b_5_14;
  assign t0_r2_c14_rr6 = a_2_6 * b_6_14;
  assign t0_r2_c14_rr7 = a_2_7 * b_7_14;
  assign t0_r2_c14_rr8 = a_2_8 * b_8_14;
  assign t0_r2_c14_rr9 = a_2_9 * b_9_14;
  assign t0_r2_c14_rr10 = a_2_10 * b_10_14;
  assign t0_r2_c14_rr11 = a_2_11 * b_11_14;
  assign t0_r2_c14_rr12 = a_2_12 * b_12_14;
  assign t0_r2_c14_rr13 = a_2_13 * b_13_14;
  assign t0_r2_c14_rr14 = a_2_14 * b_14_14;
  assign t1_r2_c14_rr0 = t0_r2_c14_rr0 + t0_r2_c14_rr1;
  assign t1_r2_c14_rr1 = t0_r2_c14_rr2 + t0_r2_c14_rr3;
  assign t1_r2_c14_rr2 = t0_r2_c14_rr4 + t0_r2_c14_rr5;
  assign t1_r2_c14_rr3 = t0_r2_c14_rr6 + t0_r2_c14_rr7;
  assign t1_r2_c14_rr4 = t0_r2_c14_rr8 + t0_r2_c14_rr9;
  assign t1_r2_c14_rr5 = t0_r2_c14_rr10 + t0_r2_c14_rr11;
  assign t1_r2_c14_rr6 = t0_r2_c14_rr12 + t0_r2_c14_rr13;
  assign t1_r2_c14_rr7 = t0_r2_c14_rr14;

  assign t2_r2_c14_rr0 = t1_r2_c14_rr0 + t1_r2_c14_rr1;
  assign t2_r2_c14_rr1 = t1_r2_c14_rr2 + t1_r2_c14_rr3;
  assign t2_r2_c14_rr2 = t1_r2_c14_rr4 + t1_r2_c14_rr5;
  assign t2_r2_c14_rr3 = t1_r2_c14_rr6 + t1_r2_c14_rr7;

  assign t3_r2_c14_rr0 = t2_r2_c14_rr0 + t2_r2_c14_rr1;
  assign t3_r2_c14_rr1 = t2_r2_c14_rr2 + t2_r2_c14_rr3;

  assign t4_r2_c14_rr0 = t3_r2_c14_rr0 + t3_r2_c14_rr1;

  assign c_2_14 = t4_r2_c14_rr0;
  assign t0_r3_c0_rr0 = a_3_0 * b_0_0;
  assign t0_r3_c0_rr1 = a_3_1 * b_1_0;
  assign t0_r3_c0_rr2 = a_3_2 * b_2_0;
  assign t0_r3_c0_rr3 = a_3_3 * b_3_0;
  assign t0_r3_c0_rr4 = a_3_4 * b_4_0;
  assign t0_r3_c0_rr5 = a_3_5 * b_5_0;
  assign t0_r3_c0_rr6 = a_3_6 * b_6_0;
  assign t0_r3_c0_rr7 = a_3_7 * b_7_0;
  assign t0_r3_c0_rr8 = a_3_8 * b_8_0;
  assign t0_r3_c0_rr9 = a_3_9 * b_9_0;
  assign t0_r3_c0_rr10 = a_3_10 * b_10_0;
  assign t0_r3_c0_rr11 = a_3_11 * b_11_0;
  assign t0_r3_c0_rr12 = a_3_12 * b_12_0;
  assign t0_r3_c0_rr13 = a_3_13 * b_13_0;
  assign t0_r3_c0_rr14 = a_3_14 * b_14_0;
  assign t1_r3_c0_rr0 = t0_r3_c0_rr0 + t0_r3_c0_rr1;
  assign t1_r3_c0_rr1 = t0_r3_c0_rr2 + t0_r3_c0_rr3;
  assign t1_r3_c0_rr2 = t0_r3_c0_rr4 + t0_r3_c0_rr5;
  assign t1_r3_c0_rr3 = t0_r3_c0_rr6 + t0_r3_c0_rr7;
  assign t1_r3_c0_rr4 = t0_r3_c0_rr8 + t0_r3_c0_rr9;
  assign t1_r3_c0_rr5 = t0_r3_c0_rr10 + t0_r3_c0_rr11;
  assign t1_r3_c0_rr6 = t0_r3_c0_rr12 + t0_r3_c0_rr13;
  assign t1_r3_c0_rr7 = t0_r3_c0_rr14;

  assign t2_r3_c0_rr0 = t1_r3_c0_rr0 + t1_r3_c0_rr1;
  assign t2_r3_c0_rr1 = t1_r3_c0_rr2 + t1_r3_c0_rr3;
  assign t2_r3_c0_rr2 = t1_r3_c0_rr4 + t1_r3_c0_rr5;
  assign t2_r3_c0_rr3 = t1_r3_c0_rr6 + t1_r3_c0_rr7;

  assign t3_r3_c0_rr0 = t2_r3_c0_rr0 + t2_r3_c0_rr1;
  assign t3_r3_c0_rr1 = t2_r3_c0_rr2 + t2_r3_c0_rr3;

  assign t4_r3_c0_rr0 = t3_r3_c0_rr0 + t3_r3_c0_rr1;

  assign c_3_0 = t4_r3_c0_rr0;
  assign t0_r3_c1_rr0 = a_3_0 * b_0_1;
  assign t0_r3_c1_rr1 = a_3_1 * b_1_1;
  assign t0_r3_c1_rr2 = a_3_2 * b_2_1;
  assign t0_r3_c1_rr3 = a_3_3 * b_3_1;
  assign t0_r3_c1_rr4 = a_3_4 * b_4_1;
  assign t0_r3_c1_rr5 = a_3_5 * b_5_1;
  assign t0_r3_c1_rr6 = a_3_6 * b_6_1;
  assign t0_r3_c1_rr7 = a_3_7 * b_7_1;
  assign t0_r3_c1_rr8 = a_3_8 * b_8_1;
  assign t0_r3_c1_rr9 = a_3_9 * b_9_1;
  assign t0_r3_c1_rr10 = a_3_10 * b_10_1;
  assign t0_r3_c1_rr11 = a_3_11 * b_11_1;
  assign t0_r3_c1_rr12 = a_3_12 * b_12_1;
  assign t0_r3_c1_rr13 = a_3_13 * b_13_1;
  assign t0_r3_c1_rr14 = a_3_14 * b_14_1;
  assign t1_r3_c1_rr0 = t0_r3_c1_rr0 + t0_r3_c1_rr1;
  assign t1_r3_c1_rr1 = t0_r3_c1_rr2 + t0_r3_c1_rr3;
  assign t1_r3_c1_rr2 = t0_r3_c1_rr4 + t0_r3_c1_rr5;
  assign t1_r3_c1_rr3 = t0_r3_c1_rr6 + t0_r3_c1_rr7;
  assign t1_r3_c1_rr4 = t0_r3_c1_rr8 + t0_r3_c1_rr9;
  assign t1_r3_c1_rr5 = t0_r3_c1_rr10 + t0_r3_c1_rr11;
  assign t1_r3_c1_rr6 = t0_r3_c1_rr12 + t0_r3_c1_rr13;
  assign t1_r3_c1_rr7 = t0_r3_c1_rr14;

  assign t2_r3_c1_rr0 = t1_r3_c1_rr0 + t1_r3_c1_rr1;
  assign t2_r3_c1_rr1 = t1_r3_c1_rr2 + t1_r3_c1_rr3;
  assign t2_r3_c1_rr2 = t1_r3_c1_rr4 + t1_r3_c1_rr5;
  assign t2_r3_c1_rr3 = t1_r3_c1_rr6 + t1_r3_c1_rr7;

  assign t3_r3_c1_rr0 = t2_r3_c1_rr0 + t2_r3_c1_rr1;
  assign t3_r3_c1_rr1 = t2_r3_c1_rr2 + t2_r3_c1_rr3;

  assign t4_r3_c1_rr0 = t3_r3_c1_rr0 + t3_r3_c1_rr1;

  assign c_3_1 = t4_r3_c1_rr0;
  assign t0_r3_c2_rr0 = a_3_0 * b_0_2;
  assign t0_r3_c2_rr1 = a_3_1 * b_1_2;
  assign t0_r3_c2_rr2 = a_3_2 * b_2_2;
  assign t0_r3_c2_rr3 = a_3_3 * b_3_2;
  assign t0_r3_c2_rr4 = a_3_4 * b_4_2;
  assign t0_r3_c2_rr5 = a_3_5 * b_5_2;
  assign t0_r3_c2_rr6 = a_3_6 * b_6_2;
  assign t0_r3_c2_rr7 = a_3_7 * b_7_2;
  assign t0_r3_c2_rr8 = a_3_8 * b_8_2;
  assign t0_r3_c2_rr9 = a_3_9 * b_9_2;
  assign t0_r3_c2_rr10 = a_3_10 * b_10_2;
  assign t0_r3_c2_rr11 = a_3_11 * b_11_2;
  assign t0_r3_c2_rr12 = a_3_12 * b_12_2;
  assign t0_r3_c2_rr13 = a_3_13 * b_13_2;
  assign t0_r3_c2_rr14 = a_3_14 * b_14_2;
  assign t1_r3_c2_rr0 = t0_r3_c2_rr0 + t0_r3_c2_rr1;
  assign t1_r3_c2_rr1 = t0_r3_c2_rr2 + t0_r3_c2_rr3;
  assign t1_r3_c2_rr2 = t0_r3_c2_rr4 + t0_r3_c2_rr5;
  assign t1_r3_c2_rr3 = t0_r3_c2_rr6 + t0_r3_c2_rr7;
  assign t1_r3_c2_rr4 = t0_r3_c2_rr8 + t0_r3_c2_rr9;
  assign t1_r3_c2_rr5 = t0_r3_c2_rr10 + t0_r3_c2_rr11;
  assign t1_r3_c2_rr6 = t0_r3_c2_rr12 + t0_r3_c2_rr13;
  assign t1_r3_c2_rr7 = t0_r3_c2_rr14;

  assign t2_r3_c2_rr0 = t1_r3_c2_rr0 + t1_r3_c2_rr1;
  assign t2_r3_c2_rr1 = t1_r3_c2_rr2 + t1_r3_c2_rr3;
  assign t2_r3_c2_rr2 = t1_r3_c2_rr4 + t1_r3_c2_rr5;
  assign t2_r3_c2_rr3 = t1_r3_c2_rr6 + t1_r3_c2_rr7;

  assign t3_r3_c2_rr0 = t2_r3_c2_rr0 + t2_r3_c2_rr1;
  assign t3_r3_c2_rr1 = t2_r3_c2_rr2 + t2_r3_c2_rr3;

  assign t4_r3_c2_rr0 = t3_r3_c2_rr0 + t3_r3_c2_rr1;

  assign c_3_2 = t4_r3_c2_rr0;
  assign t0_r3_c3_rr0 = a_3_0 * b_0_3;
  assign t0_r3_c3_rr1 = a_3_1 * b_1_3;
  assign t0_r3_c3_rr2 = a_3_2 * b_2_3;
  assign t0_r3_c3_rr3 = a_3_3 * b_3_3;
  assign t0_r3_c3_rr4 = a_3_4 * b_4_3;
  assign t0_r3_c3_rr5 = a_3_5 * b_5_3;
  assign t0_r3_c3_rr6 = a_3_6 * b_6_3;
  assign t0_r3_c3_rr7 = a_3_7 * b_7_3;
  assign t0_r3_c3_rr8 = a_3_8 * b_8_3;
  assign t0_r3_c3_rr9 = a_3_9 * b_9_3;
  assign t0_r3_c3_rr10 = a_3_10 * b_10_3;
  assign t0_r3_c3_rr11 = a_3_11 * b_11_3;
  assign t0_r3_c3_rr12 = a_3_12 * b_12_3;
  assign t0_r3_c3_rr13 = a_3_13 * b_13_3;
  assign t0_r3_c3_rr14 = a_3_14 * b_14_3;
  assign t1_r3_c3_rr0 = t0_r3_c3_rr0 + t0_r3_c3_rr1;
  assign t1_r3_c3_rr1 = t0_r3_c3_rr2 + t0_r3_c3_rr3;
  assign t1_r3_c3_rr2 = t0_r3_c3_rr4 + t0_r3_c3_rr5;
  assign t1_r3_c3_rr3 = t0_r3_c3_rr6 + t0_r3_c3_rr7;
  assign t1_r3_c3_rr4 = t0_r3_c3_rr8 + t0_r3_c3_rr9;
  assign t1_r3_c3_rr5 = t0_r3_c3_rr10 + t0_r3_c3_rr11;
  assign t1_r3_c3_rr6 = t0_r3_c3_rr12 + t0_r3_c3_rr13;
  assign t1_r3_c3_rr7 = t0_r3_c3_rr14;

  assign t2_r3_c3_rr0 = t1_r3_c3_rr0 + t1_r3_c3_rr1;
  assign t2_r3_c3_rr1 = t1_r3_c3_rr2 + t1_r3_c3_rr3;
  assign t2_r3_c3_rr2 = t1_r3_c3_rr4 + t1_r3_c3_rr5;
  assign t2_r3_c3_rr3 = t1_r3_c3_rr6 + t1_r3_c3_rr7;

  assign t3_r3_c3_rr0 = t2_r3_c3_rr0 + t2_r3_c3_rr1;
  assign t3_r3_c3_rr1 = t2_r3_c3_rr2 + t2_r3_c3_rr3;

  assign t4_r3_c3_rr0 = t3_r3_c3_rr0 + t3_r3_c3_rr1;

  assign c_3_3 = t4_r3_c3_rr0;
  assign t0_r3_c4_rr0 = a_3_0 * b_0_4;
  assign t0_r3_c4_rr1 = a_3_1 * b_1_4;
  assign t0_r3_c4_rr2 = a_3_2 * b_2_4;
  assign t0_r3_c4_rr3 = a_3_3 * b_3_4;
  assign t0_r3_c4_rr4 = a_3_4 * b_4_4;
  assign t0_r3_c4_rr5 = a_3_5 * b_5_4;
  assign t0_r3_c4_rr6 = a_3_6 * b_6_4;
  assign t0_r3_c4_rr7 = a_3_7 * b_7_4;
  assign t0_r3_c4_rr8 = a_3_8 * b_8_4;
  assign t0_r3_c4_rr9 = a_3_9 * b_9_4;
  assign t0_r3_c4_rr10 = a_3_10 * b_10_4;
  assign t0_r3_c4_rr11 = a_3_11 * b_11_4;
  assign t0_r3_c4_rr12 = a_3_12 * b_12_4;
  assign t0_r3_c4_rr13 = a_3_13 * b_13_4;
  assign t0_r3_c4_rr14 = a_3_14 * b_14_4;
  assign t1_r3_c4_rr0 = t0_r3_c4_rr0 + t0_r3_c4_rr1;
  assign t1_r3_c4_rr1 = t0_r3_c4_rr2 + t0_r3_c4_rr3;
  assign t1_r3_c4_rr2 = t0_r3_c4_rr4 + t0_r3_c4_rr5;
  assign t1_r3_c4_rr3 = t0_r3_c4_rr6 + t0_r3_c4_rr7;
  assign t1_r3_c4_rr4 = t0_r3_c4_rr8 + t0_r3_c4_rr9;
  assign t1_r3_c4_rr5 = t0_r3_c4_rr10 + t0_r3_c4_rr11;
  assign t1_r3_c4_rr6 = t0_r3_c4_rr12 + t0_r3_c4_rr13;
  assign t1_r3_c4_rr7 = t0_r3_c4_rr14;

  assign t2_r3_c4_rr0 = t1_r3_c4_rr0 + t1_r3_c4_rr1;
  assign t2_r3_c4_rr1 = t1_r3_c4_rr2 + t1_r3_c4_rr3;
  assign t2_r3_c4_rr2 = t1_r3_c4_rr4 + t1_r3_c4_rr5;
  assign t2_r3_c4_rr3 = t1_r3_c4_rr6 + t1_r3_c4_rr7;

  assign t3_r3_c4_rr0 = t2_r3_c4_rr0 + t2_r3_c4_rr1;
  assign t3_r3_c4_rr1 = t2_r3_c4_rr2 + t2_r3_c4_rr3;

  assign t4_r3_c4_rr0 = t3_r3_c4_rr0 + t3_r3_c4_rr1;

  assign c_3_4 = t4_r3_c4_rr0;
  assign t0_r3_c5_rr0 = a_3_0 * b_0_5;
  assign t0_r3_c5_rr1 = a_3_1 * b_1_5;
  assign t0_r3_c5_rr2 = a_3_2 * b_2_5;
  assign t0_r3_c5_rr3 = a_3_3 * b_3_5;
  assign t0_r3_c5_rr4 = a_3_4 * b_4_5;
  assign t0_r3_c5_rr5 = a_3_5 * b_5_5;
  assign t0_r3_c5_rr6 = a_3_6 * b_6_5;
  assign t0_r3_c5_rr7 = a_3_7 * b_7_5;
  assign t0_r3_c5_rr8 = a_3_8 * b_8_5;
  assign t0_r3_c5_rr9 = a_3_9 * b_9_5;
  assign t0_r3_c5_rr10 = a_3_10 * b_10_5;
  assign t0_r3_c5_rr11 = a_3_11 * b_11_5;
  assign t0_r3_c5_rr12 = a_3_12 * b_12_5;
  assign t0_r3_c5_rr13 = a_3_13 * b_13_5;
  assign t0_r3_c5_rr14 = a_3_14 * b_14_5;
  assign t1_r3_c5_rr0 = t0_r3_c5_rr0 + t0_r3_c5_rr1;
  assign t1_r3_c5_rr1 = t0_r3_c5_rr2 + t0_r3_c5_rr3;
  assign t1_r3_c5_rr2 = t0_r3_c5_rr4 + t0_r3_c5_rr5;
  assign t1_r3_c5_rr3 = t0_r3_c5_rr6 + t0_r3_c5_rr7;
  assign t1_r3_c5_rr4 = t0_r3_c5_rr8 + t0_r3_c5_rr9;
  assign t1_r3_c5_rr5 = t0_r3_c5_rr10 + t0_r3_c5_rr11;
  assign t1_r3_c5_rr6 = t0_r3_c5_rr12 + t0_r3_c5_rr13;
  assign t1_r3_c5_rr7 = t0_r3_c5_rr14;

  assign t2_r3_c5_rr0 = t1_r3_c5_rr0 + t1_r3_c5_rr1;
  assign t2_r3_c5_rr1 = t1_r3_c5_rr2 + t1_r3_c5_rr3;
  assign t2_r3_c5_rr2 = t1_r3_c5_rr4 + t1_r3_c5_rr5;
  assign t2_r3_c5_rr3 = t1_r3_c5_rr6 + t1_r3_c5_rr7;

  assign t3_r3_c5_rr0 = t2_r3_c5_rr0 + t2_r3_c5_rr1;
  assign t3_r3_c5_rr1 = t2_r3_c5_rr2 + t2_r3_c5_rr3;

  assign t4_r3_c5_rr0 = t3_r3_c5_rr0 + t3_r3_c5_rr1;

  assign c_3_5 = t4_r3_c5_rr0;
  assign t0_r3_c6_rr0 = a_3_0 * b_0_6;
  assign t0_r3_c6_rr1 = a_3_1 * b_1_6;
  assign t0_r3_c6_rr2 = a_3_2 * b_2_6;
  assign t0_r3_c6_rr3 = a_3_3 * b_3_6;
  assign t0_r3_c6_rr4 = a_3_4 * b_4_6;
  assign t0_r3_c6_rr5 = a_3_5 * b_5_6;
  assign t0_r3_c6_rr6 = a_3_6 * b_6_6;
  assign t0_r3_c6_rr7 = a_3_7 * b_7_6;
  assign t0_r3_c6_rr8 = a_3_8 * b_8_6;
  assign t0_r3_c6_rr9 = a_3_9 * b_9_6;
  assign t0_r3_c6_rr10 = a_3_10 * b_10_6;
  assign t0_r3_c6_rr11 = a_3_11 * b_11_6;
  assign t0_r3_c6_rr12 = a_3_12 * b_12_6;
  assign t0_r3_c6_rr13 = a_3_13 * b_13_6;
  assign t0_r3_c6_rr14 = a_3_14 * b_14_6;
  assign t1_r3_c6_rr0 = t0_r3_c6_rr0 + t0_r3_c6_rr1;
  assign t1_r3_c6_rr1 = t0_r3_c6_rr2 + t0_r3_c6_rr3;
  assign t1_r3_c6_rr2 = t0_r3_c6_rr4 + t0_r3_c6_rr5;
  assign t1_r3_c6_rr3 = t0_r3_c6_rr6 + t0_r3_c6_rr7;
  assign t1_r3_c6_rr4 = t0_r3_c6_rr8 + t0_r3_c6_rr9;
  assign t1_r3_c6_rr5 = t0_r3_c6_rr10 + t0_r3_c6_rr11;
  assign t1_r3_c6_rr6 = t0_r3_c6_rr12 + t0_r3_c6_rr13;
  assign t1_r3_c6_rr7 = t0_r3_c6_rr14;

  assign t2_r3_c6_rr0 = t1_r3_c6_rr0 + t1_r3_c6_rr1;
  assign t2_r3_c6_rr1 = t1_r3_c6_rr2 + t1_r3_c6_rr3;
  assign t2_r3_c6_rr2 = t1_r3_c6_rr4 + t1_r3_c6_rr5;
  assign t2_r3_c6_rr3 = t1_r3_c6_rr6 + t1_r3_c6_rr7;

  assign t3_r3_c6_rr0 = t2_r3_c6_rr0 + t2_r3_c6_rr1;
  assign t3_r3_c6_rr1 = t2_r3_c6_rr2 + t2_r3_c6_rr3;

  assign t4_r3_c6_rr0 = t3_r3_c6_rr0 + t3_r3_c6_rr1;

  assign c_3_6 = t4_r3_c6_rr0;
  assign t0_r3_c7_rr0 = a_3_0 * b_0_7;
  assign t0_r3_c7_rr1 = a_3_1 * b_1_7;
  assign t0_r3_c7_rr2 = a_3_2 * b_2_7;
  assign t0_r3_c7_rr3 = a_3_3 * b_3_7;
  assign t0_r3_c7_rr4 = a_3_4 * b_4_7;
  assign t0_r3_c7_rr5 = a_3_5 * b_5_7;
  assign t0_r3_c7_rr6 = a_3_6 * b_6_7;
  assign t0_r3_c7_rr7 = a_3_7 * b_7_7;
  assign t0_r3_c7_rr8 = a_3_8 * b_8_7;
  assign t0_r3_c7_rr9 = a_3_9 * b_9_7;
  assign t0_r3_c7_rr10 = a_3_10 * b_10_7;
  assign t0_r3_c7_rr11 = a_3_11 * b_11_7;
  assign t0_r3_c7_rr12 = a_3_12 * b_12_7;
  assign t0_r3_c7_rr13 = a_3_13 * b_13_7;
  assign t0_r3_c7_rr14 = a_3_14 * b_14_7;
  assign t1_r3_c7_rr0 = t0_r3_c7_rr0 + t0_r3_c7_rr1;
  assign t1_r3_c7_rr1 = t0_r3_c7_rr2 + t0_r3_c7_rr3;
  assign t1_r3_c7_rr2 = t0_r3_c7_rr4 + t0_r3_c7_rr5;
  assign t1_r3_c7_rr3 = t0_r3_c7_rr6 + t0_r3_c7_rr7;
  assign t1_r3_c7_rr4 = t0_r3_c7_rr8 + t0_r3_c7_rr9;
  assign t1_r3_c7_rr5 = t0_r3_c7_rr10 + t0_r3_c7_rr11;
  assign t1_r3_c7_rr6 = t0_r3_c7_rr12 + t0_r3_c7_rr13;
  assign t1_r3_c7_rr7 = t0_r3_c7_rr14;

  assign t2_r3_c7_rr0 = t1_r3_c7_rr0 + t1_r3_c7_rr1;
  assign t2_r3_c7_rr1 = t1_r3_c7_rr2 + t1_r3_c7_rr3;
  assign t2_r3_c7_rr2 = t1_r3_c7_rr4 + t1_r3_c7_rr5;
  assign t2_r3_c7_rr3 = t1_r3_c7_rr6 + t1_r3_c7_rr7;

  assign t3_r3_c7_rr0 = t2_r3_c7_rr0 + t2_r3_c7_rr1;
  assign t3_r3_c7_rr1 = t2_r3_c7_rr2 + t2_r3_c7_rr3;

  assign t4_r3_c7_rr0 = t3_r3_c7_rr0 + t3_r3_c7_rr1;

  assign c_3_7 = t4_r3_c7_rr0;
  assign t0_r3_c8_rr0 = a_3_0 * b_0_8;
  assign t0_r3_c8_rr1 = a_3_1 * b_1_8;
  assign t0_r3_c8_rr2 = a_3_2 * b_2_8;
  assign t0_r3_c8_rr3 = a_3_3 * b_3_8;
  assign t0_r3_c8_rr4 = a_3_4 * b_4_8;
  assign t0_r3_c8_rr5 = a_3_5 * b_5_8;
  assign t0_r3_c8_rr6 = a_3_6 * b_6_8;
  assign t0_r3_c8_rr7 = a_3_7 * b_7_8;
  assign t0_r3_c8_rr8 = a_3_8 * b_8_8;
  assign t0_r3_c8_rr9 = a_3_9 * b_9_8;
  assign t0_r3_c8_rr10 = a_3_10 * b_10_8;
  assign t0_r3_c8_rr11 = a_3_11 * b_11_8;
  assign t0_r3_c8_rr12 = a_3_12 * b_12_8;
  assign t0_r3_c8_rr13 = a_3_13 * b_13_8;
  assign t0_r3_c8_rr14 = a_3_14 * b_14_8;
  assign t1_r3_c8_rr0 = t0_r3_c8_rr0 + t0_r3_c8_rr1;
  assign t1_r3_c8_rr1 = t0_r3_c8_rr2 + t0_r3_c8_rr3;
  assign t1_r3_c8_rr2 = t0_r3_c8_rr4 + t0_r3_c8_rr5;
  assign t1_r3_c8_rr3 = t0_r3_c8_rr6 + t0_r3_c8_rr7;
  assign t1_r3_c8_rr4 = t0_r3_c8_rr8 + t0_r3_c8_rr9;
  assign t1_r3_c8_rr5 = t0_r3_c8_rr10 + t0_r3_c8_rr11;
  assign t1_r3_c8_rr6 = t0_r3_c8_rr12 + t0_r3_c8_rr13;
  assign t1_r3_c8_rr7 = t0_r3_c8_rr14;

  assign t2_r3_c8_rr0 = t1_r3_c8_rr0 + t1_r3_c8_rr1;
  assign t2_r3_c8_rr1 = t1_r3_c8_rr2 + t1_r3_c8_rr3;
  assign t2_r3_c8_rr2 = t1_r3_c8_rr4 + t1_r3_c8_rr5;
  assign t2_r3_c8_rr3 = t1_r3_c8_rr6 + t1_r3_c8_rr7;

  assign t3_r3_c8_rr0 = t2_r3_c8_rr0 + t2_r3_c8_rr1;
  assign t3_r3_c8_rr1 = t2_r3_c8_rr2 + t2_r3_c8_rr3;

  assign t4_r3_c8_rr0 = t3_r3_c8_rr0 + t3_r3_c8_rr1;

  assign c_3_8 = t4_r3_c8_rr0;
  assign t0_r3_c9_rr0 = a_3_0 * b_0_9;
  assign t0_r3_c9_rr1 = a_3_1 * b_1_9;
  assign t0_r3_c9_rr2 = a_3_2 * b_2_9;
  assign t0_r3_c9_rr3 = a_3_3 * b_3_9;
  assign t0_r3_c9_rr4 = a_3_4 * b_4_9;
  assign t0_r3_c9_rr5 = a_3_5 * b_5_9;
  assign t0_r3_c9_rr6 = a_3_6 * b_6_9;
  assign t0_r3_c9_rr7 = a_3_7 * b_7_9;
  assign t0_r3_c9_rr8 = a_3_8 * b_8_9;
  assign t0_r3_c9_rr9 = a_3_9 * b_9_9;
  assign t0_r3_c9_rr10 = a_3_10 * b_10_9;
  assign t0_r3_c9_rr11 = a_3_11 * b_11_9;
  assign t0_r3_c9_rr12 = a_3_12 * b_12_9;
  assign t0_r3_c9_rr13 = a_3_13 * b_13_9;
  assign t0_r3_c9_rr14 = a_3_14 * b_14_9;
  assign t1_r3_c9_rr0 = t0_r3_c9_rr0 + t0_r3_c9_rr1;
  assign t1_r3_c9_rr1 = t0_r3_c9_rr2 + t0_r3_c9_rr3;
  assign t1_r3_c9_rr2 = t0_r3_c9_rr4 + t0_r3_c9_rr5;
  assign t1_r3_c9_rr3 = t0_r3_c9_rr6 + t0_r3_c9_rr7;
  assign t1_r3_c9_rr4 = t0_r3_c9_rr8 + t0_r3_c9_rr9;
  assign t1_r3_c9_rr5 = t0_r3_c9_rr10 + t0_r3_c9_rr11;
  assign t1_r3_c9_rr6 = t0_r3_c9_rr12 + t0_r3_c9_rr13;
  assign t1_r3_c9_rr7 = t0_r3_c9_rr14;

  assign t2_r3_c9_rr0 = t1_r3_c9_rr0 + t1_r3_c9_rr1;
  assign t2_r3_c9_rr1 = t1_r3_c9_rr2 + t1_r3_c9_rr3;
  assign t2_r3_c9_rr2 = t1_r3_c9_rr4 + t1_r3_c9_rr5;
  assign t2_r3_c9_rr3 = t1_r3_c9_rr6 + t1_r3_c9_rr7;

  assign t3_r3_c9_rr0 = t2_r3_c9_rr0 + t2_r3_c9_rr1;
  assign t3_r3_c9_rr1 = t2_r3_c9_rr2 + t2_r3_c9_rr3;

  assign t4_r3_c9_rr0 = t3_r3_c9_rr0 + t3_r3_c9_rr1;

  assign c_3_9 = t4_r3_c9_rr0;
  assign t0_r3_c10_rr0 = a_3_0 * b_0_10;
  assign t0_r3_c10_rr1 = a_3_1 * b_1_10;
  assign t0_r3_c10_rr2 = a_3_2 * b_2_10;
  assign t0_r3_c10_rr3 = a_3_3 * b_3_10;
  assign t0_r3_c10_rr4 = a_3_4 * b_4_10;
  assign t0_r3_c10_rr5 = a_3_5 * b_5_10;
  assign t0_r3_c10_rr6 = a_3_6 * b_6_10;
  assign t0_r3_c10_rr7 = a_3_7 * b_7_10;
  assign t0_r3_c10_rr8 = a_3_8 * b_8_10;
  assign t0_r3_c10_rr9 = a_3_9 * b_9_10;
  assign t0_r3_c10_rr10 = a_3_10 * b_10_10;
  assign t0_r3_c10_rr11 = a_3_11 * b_11_10;
  assign t0_r3_c10_rr12 = a_3_12 * b_12_10;
  assign t0_r3_c10_rr13 = a_3_13 * b_13_10;
  assign t0_r3_c10_rr14 = a_3_14 * b_14_10;
  assign t1_r3_c10_rr0 = t0_r3_c10_rr0 + t0_r3_c10_rr1;
  assign t1_r3_c10_rr1 = t0_r3_c10_rr2 + t0_r3_c10_rr3;
  assign t1_r3_c10_rr2 = t0_r3_c10_rr4 + t0_r3_c10_rr5;
  assign t1_r3_c10_rr3 = t0_r3_c10_rr6 + t0_r3_c10_rr7;
  assign t1_r3_c10_rr4 = t0_r3_c10_rr8 + t0_r3_c10_rr9;
  assign t1_r3_c10_rr5 = t0_r3_c10_rr10 + t0_r3_c10_rr11;
  assign t1_r3_c10_rr6 = t0_r3_c10_rr12 + t0_r3_c10_rr13;
  assign t1_r3_c10_rr7 = t0_r3_c10_rr14;

  assign t2_r3_c10_rr0 = t1_r3_c10_rr0 + t1_r3_c10_rr1;
  assign t2_r3_c10_rr1 = t1_r3_c10_rr2 + t1_r3_c10_rr3;
  assign t2_r3_c10_rr2 = t1_r3_c10_rr4 + t1_r3_c10_rr5;
  assign t2_r3_c10_rr3 = t1_r3_c10_rr6 + t1_r3_c10_rr7;

  assign t3_r3_c10_rr0 = t2_r3_c10_rr0 + t2_r3_c10_rr1;
  assign t3_r3_c10_rr1 = t2_r3_c10_rr2 + t2_r3_c10_rr3;

  assign t4_r3_c10_rr0 = t3_r3_c10_rr0 + t3_r3_c10_rr1;

  assign c_3_10 = t4_r3_c10_rr0;
  assign t0_r3_c11_rr0 = a_3_0 * b_0_11;
  assign t0_r3_c11_rr1 = a_3_1 * b_1_11;
  assign t0_r3_c11_rr2 = a_3_2 * b_2_11;
  assign t0_r3_c11_rr3 = a_3_3 * b_3_11;
  assign t0_r3_c11_rr4 = a_3_4 * b_4_11;
  assign t0_r3_c11_rr5 = a_3_5 * b_5_11;
  assign t0_r3_c11_rr6 = a_3_6 * b_6_11;
  assign t0_r3_c11_rr7 = a_3_7 * b_7_11;
  assign t0_r3_c11_rr8 = a_3_8 * b_8_11;
  assign t0_r3_c11_rr9 = a_3_9 * b_9_11;
  assign t0_r3_c11_rr10 = a_3_10 * b_10_11;
  assign t0_r3_c11_rr11 = a_3_11 * b_11_11;
  assign t0_r3_c11_rr12 = a_3_12 * b_12_11;
  assign t0_r3_c11_rr13 = a_3_13 * b_13_11;
  assign t0_r3_c11_rr14 = a_3_14 * b_14_11;
  assign t1_r3_c11_rr0 = t0_r3_c11_rr0 + t0_r3_c11_rr1;
  assign t1_r3_c11_rr1 = t0_r3_c11_rr2 + t0_r3_c11_rr3;
  assign t1_r3_c11_rr2 = t0_r3_c11_rr4 + t0_r3_c11_rr5;
  assign t1_r3_c11_rr3 = t0_r3_c11_rr6 + t0_r3_c11_rr7;
  assign t1_r3_c11_rr4 = t0_r3_c11_rr8 + t0_r3_c11_rr9;
  assign t1_r3_c11_rr5 = t0_r3_c11_rr10 + t0_r3_c11_rr11;
  assign t1_r3_c11_rr6 = t0_r3_c11_rr12 + t0_r3_c11_rr13;
  assign t1_r3_c11_rr7 = t0_r3_c11_rr14;

  assign t2_r3_c11_rr0 = t1_r3_c11_rr0 + t1_r3_c11_rr1;
  assign t2_r3_c11_rr1 = t1_r3_c11_rr2 + t1_r3_c11_rr3;
  assign t2_r3_c11_rr2 = t1_r3_c11_rr4 + t1_r3_c11_rr5;
  assign t2_r3_c11_rr3 = t1_r3_c11_rr6 + t1_r3_c11_rr7;

  assign t3_r3_c11_rr0 = t2_r3_c11_rr0 + t2_r3_c11_rr1;
  assign t3_r3_c11_rr1 = t2_r3_c11_rr2 + t2_r3_c11_rr3;

  assign t4_r3_c11_rr0 = t3_r3_c11_rr0 + t3_r3_c11_rr1;

  assign c_3_11 = t4_r3_c11_rr0;
  assign t0_r3_c12_rr0 = a_3_0 * b_0_12;
  assign t0_r3_c12_rr1 = a_3_1 * b_1_12;
  assign t0_r3_c12_rr2 = a_3_2 * b_2_12;
  assign t0_r3_c12_rr3 = a_3_3 * b_3_12;
  assign t0_r3_c12_rr4 = a_3_4 * b_4_12;
  assign t0_r3_c12_rr5 = a_3_5 * b_5_12;
  assign t0_r3_c12_rr6 = a_3_6 * b_6_12;
  assign t0_r3_c12_rr7 = a_3_7 * b_7_12;
  assign t0_r3_c12_rr8 = a_3_8 * b_8_12;
  assign t0_r3_c12_rr9 = a_3_9 * b_9_12;
  assign t0_r3_c12_rr10 = a_3_10 * b_10_12;
  assign t0_r3_c12_rr11 = a_3_11 * b_11_12;
  assign t0_r3_c12_rr12 = a_3_12 * b_12_12;
  assign t0_r3_c12_rr13 = a_3_13 * b_13_12;
  assign t0_r3_c12_rr14 = a_3_14 * b_14_12;
  assign t1_r3_c12_rr0 = t0_r3_c12_rr0 + t0_r3_c12_rr1;
  assign t1_r3_c12_rr1 = t0_r3_c12_rr2 + t0_r3_c12_rr3;
  assign t1_r3_c12_rr2 = t0_r3_c12_rr4 + t0_r3_c12_rr5;
  assign t1_r3_c12_rr3 = t0_r3_c12_rr6 + t0_r3_c12_rr7;
  assign t1_r3_c12_rr4 = t0_r3_c12_rr8 + t0_r3_c12_rr9;
  assign t1_r3_c12_rr5 = t0_r3_c12_rr10 + t0_r3_c12_rr11;
  assign t1_r3_c12_rr6 = t0_r3_c12_rr12 + t0_r3_c12_rr13;
  assign t1_r3_c12_rr7 = t0_r3_c12_rr14;

  assign t2_r3_c12_rr0 = t1_r3_c12_rr0 + t1_r3_c12_rr1;
  assign t2_r3_c12_rr1 = t1_r3_c12_rr2 + t1_r3_c12_rr3;
  assign t2_r3_c12_rr2 = t1_r3_c12_rr4 + t1_r3_c12_rr5;
  assign t2_r3_c12_rr3 = t1_r3_c12_rr6 + t1_r3_c12_rr7;

  assign t3_r3_c12_rr0 = t2_r3_c12_rr0 + t2_r3_c12_rr1;
  assign t3_r3_c12_rr1 = t2_r3_c12_rr2 + t2_r3_c12_rr3;

  assign t4_r3_c12_rr0 = t3_r3_c12_rr0 + t3_r3_c12_rr1;

  assign c_3_12 = t4_r3_c12_rr0;
  assign t0_r3_c13_rr0 = a_3_0 * b_0_13;
  assign t0_r3_c13_rr1 = a_3_1 * b_1_13;
  assign t0_r3_c13_rr2 = a_3_2 * b_2_13;
  assign t0_r3_c13_rr3 = a_3_3 * b_3_13;
  assign t0_r3_c13_rr4 = a_3_4 * b_4_13;
  assign t0_r3_c13_rr5 = a_3_5 * b_5_13;
  assign t0_r3_c13_rr6 = a_3_6 * b_6_13;
  assign t0_r3_c13_rr7 = a_3_7 * b_7_13;
  assign t0_r3_c13_rr8 = a_3_8 * b_8_13;
  assign t0_r3_c13_rr9 = a_3_9 * b_9_13;
  assign t0_r3_c13_rr10 = a_3_10 * b_10_13;
  assign t0_r3_c13_rr11 = a_3_11 * b_11_13;
  assign t0_r3_c13_rr12 = a_3_12 * b_12_13;
  assign t0_r3_c13_rr13 = a_3_13 * b_13_13;
  assign t0_r3_c13_rr14 = a_3_14 * b_14_13;
  assign t1_r3_c13_rr0 = t0_r3_c13_rr0 + t0_r3_c13_rr1;
  assign t1_r3_c13_rr1 = t0_r3_c13_rr2 + t0_r3_c13_rr3;
  assign t1_r3_c13_rr2 = t0_r3_c13_rr4 + t0_r3_c13_rr5;
  assign t1_r3_c13_rr3 = t0_r3_c13_rr6 + t0_r3_c13_rr7;
  assign t1_r3_c13_rr4 = t0_r3_c13_rr8 + t0_r3_c13_rr9;
  assign t1_r3_c13_rr5 = t0_r3_c13_rr10 + t0_r3_c13_rr11;
  assign t1_r3_c13_rr6 = t0_r3_c13_rr12 + t0_r3_c13_rr13;
  assign t1_r3_c13_rr7 = t0_r3_c13_rr14;

  assign t2_r3_c13_rr0 = t1_r3_c13_rr0 + t1_r3_c13_rr1;
  assign t2_r3_c13_rr1 = t1_r3_c13_rr2 + t1_r3_c13_rr3;
  assign t2_r3_c13_rr2 = t1_r3_c13_rr4 + t1_r3_c13_rr5;
  assign t2_r3_c13_rr3 = t1_r3_c13_rr6 + t1_r3_c13_rr7;

  assign t3_r3_c13_rr0 = t2_r3_c13_rr0 + t2_r3_c13_rr1;
  assign t3_r3_c13_rr1 = t2_r3_c13_rr2 + t2_r3_c13_rr3;

  assign t4_r3_c13_rr0 = t3_r3_c13_rr0 + t3_r3_c13_rr1;

  assign c_3_13 = t4_r3_c13_rr0;
  assign t0_r3_c14_rr0 = a_3_0 * b_0_14;
  assign t0_r3_c14_rr1 = a_3_1 * b_1_14;
  assign t0_r3_c14_rr2 = a_3_2 * b_2_14;
  assign t0_r3_c14_rr3 = a_3_3 * b_3_14;
  assign t0_r3_c14_rr4 = a_3_4 * b_4_14;
  assign t0_r3_c14_rr5 = a_3_5 * b_5_14;
  assign t0_r3_c14_rr6 = a_3_6 * b_6_14;
  assign t0_r3_c14_rr7 = a_3_7 * b_7_14;
  assign t0_r3_c14_rr8 = a_3_8 * b_8_14;
  assign t0_r3_c14_rr9 = a_3_9 * b_9_14;
  assign t0_r3_c14_rr10 = a_3_10 * b_10_14;
  assign t0_r3_c14_rr11 = a_3_11 * b_11_14;
  assign t0_r3_c14_rr12 = a_3_12 * b_12_14;
  assign t0_r3_c14_rr13 = a_3_13 * b_13_14;
  assign t0_r3_c14_rr14 = a_3_14 * b_14_14;
  assign t1_r3_c14_rr0 = t0_r3_c14_rr0 + t0_r3_c14_rr1;
  assign t1_r3_c14_rr1 = t0_r3_c14_rr2 + t0_r3_c14_rr3;
  assign t1_r3_c14_rr2 = t0_r3_c14_rr4 + t0_r3_c14_rr5;
  assign t1_r3_c14_rr3 = t0_r3_c14_rr6 + t0_r3_c14_rr7;
  assign t1_r3_c14_rr4 = t0_r3_c14_rr8 + t0_r3_c14_rr9;
  assign t1_r3_c14_rr5 = t0_r3_c14_rr10 + t0_r3_c14_rr11;
  assign t1_r3_c14_rr6 = t0_r3_c14_rr12 + t0_r3_c14_rr13;
  assign t1_r3_c14_rr7 = t0_r3_c14_rr14;

  assign t2_r3_c14_rr0 = t1_r3_c14_rr0 + t1_r3_c14_rr1;
  assign t2_r3_c14_rr1 = t1_r3_c14_rr2 + t1_r3_c14_rr3;
  assign t2_r3_c14_rr2 = t1_r3_c14_rr4 + t1_r3_c14_rr5;
  assign t2_r3_c14_rr3 = t1_r3_c14_rr6 + t1_r3_c14_rr7;

  assign t3_r3_c14_rr0 = t2_r3_c14_rr0 + t2_r3_c14_rr1;
  assign t3_r3_c14_rr1 = t2_r3_c14_rr2 + t2_r3_c14_rr3;

  assign t4_r3_c14_rr0 = t3_r3_c14_rr0 + t3_r3_c14_rr1;

  assign c_3_14 = t4_r3_c14_rr0;
  assign t0_r4_c0_rr0 = a_4_0 * b_0_0;
  assign t0_r4_c0_rr1 = a_4_1 * b_1_0;
  assign t0_r4_c0_rr2 = a_4_2 * b_2_0;
  assign t0_r4_c0_rr3 = a_4_3 * b_3_0;
  assign t0_r4_c0_rr4 = a_4_4 * b_4_0;
  assign t0_r4_c0_rr5 = a_4_5 * b_5_0;
  assign t0_r4_c0_rr6 = a_4_6 * b_6_0;
  assign t0_r4_c0_rr7 = a_4_7 * b_7_0;
  assign t0_r4_c0_rr8 = a_4_8 * b_8_0;
  assign t0_r4_c0_rr9 = a_4_9 * b_9_0;
  assign t0_r4_c0_rr10 = a_4_10 * b_10_0;
  assign t0_r4_c0_rr11 = a_4_11 * b_11_0;
  assign t0_r4_c0_rr12 = a_4_12 * b_12_0;
  assign t0_r4_c0_rr13 = a_4_13 * b_13_0;
  assign t0_r4_c0_rr14 = a_4_14 * b_14_0;
  assign t1_r4_c0_rr0 = t0_r4_c0_rr0 + t0_r4_c0_rr1;
  assign t1_r4_c0_rr1 = t0_r4_c0_rr2 + t0_r4_c0_rr3;
  assign t1_r4_c0_rr2 = t0_r4_c0_rr4 + t0_r4_c0_rr5;
  assign t1_r4_c0_rr3 = t0_r4_c0_rr6 + t0_r4_c0_rr7;
  assign t1_r4_c0_rr4 = t0_r4_c0_rr8 + t0_r4_c0_rr9;
  assign t1_r4_c0_rr5 = t0_r4_c0_rr10 + t0_r4_c0_rr11;
  assign t1_r4_c0_rr6 = t0_r4_c0_rr12 + t0_r4_c0_rr13;
  assign t1_r4_c0_rr7 = t0_r4_c0_rr14;

  assign t2_r4_c0_rr0 = t1_r4_c0_rr0 + t1_r4_c0_rr1;
  assign t2_r4_c0_rr1 = t1_r4_c0_rr2 + t1_r4_c0_rr3;
  assign t2_r4_c0_rr2 = t1_r4_c0_rr4 + t1_r4_c0_rr5;
  assign t2_r4_c0_rr3 = t1_r4_c0_rr6 + t1_r4_c0_rr7;

  assign t3_r4_c0_rr0 = t2_r4_c0_rr0 + t2_r4_c0_rr1;
  assign t3_r4_c0_rr1 = t2_r4_c0_rr2 + t2_r4_c0_rr3;

  assign t4_r4_c0_rr0 = t3_r4_c0_rr0 + t3_r4_c0_rr1;

  assign c_4_0 = t4_r4_c0_rr0;
  assign t0_r4_c1_rr0 = a_4_0 * b_0_1;
  assign t0_r4_c1_rr1 = a_4_1 * b_1_1;
  assign t0_r4_c1_rr2 = a_4_2 * b_2_1;
  assign t0_r4_c1_rr3 = a_4_3 * b_3_1;
  assign t0_r4_c1_rr4 = a_4_4 * b_4_1;
  assign t0_r4_c1_rr5 = a_4_5 * b_5_1;
  assign t0_r4_c1_rr6 = a_4_6 * b_6_1;
  assign t0_r4_c1_rr7 = a_4_7 * b_7_1;
  assign t0_r4_c1_rr8 = a_4_8 * b_8_1;
  assign t0_r4_c1_rr9 = a_4_9 * b_9_1;
  assign t0_r4_c1_rr10 = a_4_10 * b_10_1;
  assign t0_r4_c1_rr11 = a_4_11 * b_11_1;
  assign t0_r4_c1_rr12 = a_4_12 * b_12_1;
  assign t0_r4_c1_rr13 = a_4_13 * b_13_1;
  assign t0_r4_c1_rr14 = a_4_14 * b_14_1;
  assign t1_r4_c1_rr0 = t0_r4_c1_rr0 + t0_r4_c1_rr1;
  assign t1_r4_c1_rr1 = t0_r4_c1_rr2 + t0_r4_c1_rr3;
  assign t1_r4_c1_rr2 = t0_r4_c1_rr4 + t0_r4_c1_rr5;
  assign t1_r4_c1_rr3 = t0_r4_c1_rr6 + t0_r4_c1_rr7;
  assign t1_r4_c1_rr4 = t0_r4_c1_rr8 + t0_r4_c1_rr9;
  assign t1_r4_c1_rr5 = t0_r4_c1_rr10 + t0_r4_c1_rr11;
  assign t1_r4_c1_rr6 = t0_r4_c1_rr12 + t0_r4_c1_rr13;
  assign t1_r4_c1_rr7 = t0_r4_c1_rr14;

  assign t2_r4_c1_rr0 = t1_r4_c1_rr0 + t1_r4_c1_rr1;
  assign t2_r4_c1_rr1 = t1_r4_c1_rr2 + t1_r4_c1_rr3;
  assign t2_r4_c1_rr2 = t1_r4_c1_rr4 + t1_r4_c1_rr5;
  assign t2_r4_c1_rr3 = t1_r4_c1_rr6 + t1_r4_c1_rr7;

  assign t3_r4_c1_rr0 = t2_r4_c1_rr0 + t2_r4_c1_rr1;
  assign t3_r4_c1_rr1 = t2_r4_c1_rr2 + t2_r4_c1_rr3;

  assign t4_r4_c1_rr0 = t3_r4_c1_rr0 + t3_r4_c1_rr1;

  assign c_4_1 = t4_r4_c1_rr0;
  assign t0_r4_c2_rr0 = a_4_0 * b_0_2;
  assign t0_r4_c2_rr1 = a_4_1 * b_1_2;
  assign t0_r4_c2_rr2 = a_4_2 * b_2_2;
  assign t0_r4_c2_rr3 = a_4_3 * b_3_2;
  assign t0_r4_c2_rr4 = a_4_4 * b_4_2;
  assign t0_r4_c2_rr5 = a_4_5 * b_5_2;
  assign t0_r4_c2_rr6 = a_4_6 * b_6_2;
  assign t0_r4_c2_rr7 = a_4_7 * b_7_2;
  assign t0_r4_c2_rr8 = a_4_8 * b_8_2;
  assign t0_r4_c2_rr9 = a_4_9 * b_9_2;
  assign t0_r4_c2_rr10 = a_4_10 * b_10_2;
  assign t0_r4_c2_rr11 = a_4_11 * b_11_2;
  assign t0_r4_c2_rr12 = a_4_12 * b_12_2;
  assign t0_r4_c2_rr13 = a_4_13 * b_13_2;
  assign t0_r4_c2_rr14 = a_4_14 * b_14_2;
  assign t1_r4_c2_rr0 = t0_r4_c2_rr0 + t0_r4_c2_rr1;
  assign t1_r4_c2_rr1 = t0_r4_c2_rr2 + t0_r4_c2_rr3;
  assign t1_r4_c2_rr2 = t0_r4_c2_rr4 + t0_r4_c2_rr5;
  assign t1_r4_c2_rr3 = t0_r4_c2_rr6 + t0_r4_c2_rr7;
  assign t1_r4_c2_rr4 = t0_r4_c2_rr8 + t0_r4_c2_rr9;
  assign t1_r4_c2_rr5 = t0_r4_c2_rr10 + t0_r4_c2_rr11;
  assign t1_r4_c2_rr6 = t0_r4_c2_rr12 + t0_r4_c2_rr13;
  assign t1_r4_c2_rr7 = t0_r4_c2_rr14;

  assign t2_r4_c2_rr0 = t1_r4_c2_rr0 + t1_r4_c2_rr1;
  assign t2_r4_c2_rr1 = t1_r4_c2_rr2 + t1_r4_c2_rr3;
  assign t2_r4_c2_rr2 = t1_r4_c2_rr4 + t1_r4_c2_rr5;
  assign t2_r4_c2_rr3 = t1_r4_c2_rr6 + t1_r4_c2_rr7;

  assign t3_r4_c2_rr0 = t2_r4_c2_rr0 + t2_r4_c2_rr1;
  assign t3_r4_c2_rr1 = t2_r4_c2_rr2 + t2_r4_c2_rr3;

  assign t4_r4_c2_rr0 = t3_r4_c2_rr0 + t3_r4_c2_rr1;

  assign c_4_2 = t4_r4_c2_rr0;
  assign t0_r4_c3_rr0 = a_4_0 * b_0_3;
  assign t0_r4_c3_rr1 = a_4_1 * b_1_3;
  assign t0_r4_c3_rr2 = a_4_2 * b_2_3;
  assign t0_r4_c3_rr3 = a_4_3 * b_3_3;
  assign t0_r4_c3_rr4 = a_4_4 * b_4_3;
  assign t0_r4_c3_rr5 = a_4_5 * b_5_3;
  assign t0_r4_c3_rr6 = a_4_6 * b_6_3;
  assign t0_r4_c3_rr7 = a_4_7 * b_7_3;
  assign t0_r4_c3_rr8 = a_4_8 * b_8_3;
  assign t0_r4_c3_rr9 = a_4_9 * b_9_3;
  assign t0_r4_c3_rr10 = a_4_10 * b_10_3;
  assign t0_r4_c3_rr11 = a_4_11 * b_11_3;
  assign t0_r4_c3_rr12 = a_4_12 * b_12_3;
  assign t0_r4_c3_rr13 = a_4_13 * b_13_3;
  assign t0_r4_c3_rr14 = a_4_14 * b_14_3;
  assign t1_r4_c3_rr0 = t0_r4_c3_rr0 + t0_r4_c3_rr1;
  assign t1_r4_c3_rr1 = t0_r4_c3_rr2 + t0_r4_c3_rr3;
  assign t1_r4_c3_rr2 = t0_r4_c3_rr4 + t0_r4_c3_rr5;
  assign t1_r4_c3_rr3 = t0_r4_c3_rr6 + t0_r4_c3_rr7;
  assign t1_r4_c3_rr4 = t0_r4_c3_rr8 + t0_r4_c3_rr9;
  assign t1_r4_c3_rr5 = t0_r4_c3_rr10 + t0_r4_c3_rr11;
  assign t1_r4_c3_rr6 = t0_r4_c3_rr12 + t0_r4_c3_rr13;
  assign t1_r4_c3_rr7 = t0_r4_c3_rr14;

  assign t2_r4_c3_rr0 = t1_r4_c3_rr0 + t1_r4_c3_rr1;
  assign t2_r4_c3_rr1 = t1_r4_c3_rr2 + t1_r4_c3_rr3;
  assign t2_r4_c3_rr2 = t1_r4_c3_rr4 + t1_r4_c3_rr5;
  assign t2_r4_c3_rr3 = t1_r4_c3_rr6 + t1_r4_c3_rr7;

  assign t3_r4_c3_rr0 = t2_r4_c3_rr0 + t2_r4_c3_rr1;
  assign t3_r4_c3_rr1 = t2_r4_c3_rr2 + t2_r4_c3_rr3;

  assign t4_r4_c3_rr0 = t3_r4_c3_rr0 + t3_r4_c3_rr1;

  assign c_4_3 = t4_r4_c3_rr0;
  assign t0_r4_c4_rr0 = a_4_0 * b_0_4;
  assign t0_r4_c4_rr1 = a_4_1 * b_1_4;
  assign t0_r4_c4_rr2 = a_4_2 * b_2_4;
  assign t0_r4_c4_rr3 = a_4_3 * b_3_4;
  assign t0_r4_c4_rr4 = a_4_4 * b_4_4;
  assign t0_r4_c4_rr5 = a_4_5 * b_5_4;
  assign t0_r4_c4_rr6 = a_4_6 * b_6_4;
  assign t0_r4_c4_rr7 = a_4_7 * b_7_4;
  assign t0_r4_c4_rr8 = a_4_8 * b_8_4;
  assign t0_r4_c4_rr9 = a_4_9 * b_9_4;
  assign t0_r4_c4_rr10 = a_4_10 * b_10_4;
  assign t0_r4_c4_rr11 = a_4_11 * b_11_4;
  assign t0_r4_c4_rr12 = a_4_12 * b_12_4;
  assign t0_r4_c4_rr13 = a_4_13 * b_13_4;
  assign t0_r4_c4_rr14 = a_4_14 * b_14_4;
  assign t1_r4_c4_rr0 = t0_r4_c4_rr0 + t0_r4_c4_rr1;
  assign t1_r4_c4_rr1 = t0_r4_c4_rr2 + t0_r4_c4_rr3;
  assign t1_r4_c4_rr2 = t0_r4_c4_rr4 + t0_r4_c4_rr5;
  assign t1_r4_c4_rr3 = t0_r4_c4_rr6 + t0_r4_c4_rr7;
  assign t1_r4_c4_rr4 = t0_r4_c4_rr8 + t0_r4_c4_rr9;
  assign t1_r4_c4_rr5 = t0_r4_c4_rr10 + t0_r4_c4_rr11;
  assign t1_r4_c4_rr6 = t0_r4_c4_rr12 + t0_r4_c4_rr13;
  assign t1_r4_c4_rr7 = t0_r4_c4_rr14;

  assign t2_r4_c4_rr0 = t1_r4_c4_rr0 + t1_r4_c4_rr1;
  assign t2_r4_c4_rr1 = t1_r4_c4_rr2 + t1_r4_c4_rr3;
  assign t2_r4_c4_rr2 = t1_r4_c4_rr4 + t1_r4_c4_rr5;
  assign t2_r4_c4_rr3 = t1_r4_c4_rr6 + t1_r4_c4_rr7;

  assign t3_r4_c4_rr0 = t2_r4_c4_rr0 + t2_r4_c4_rr1;
  assign t3_r4_c4_rr1 = t2_r4_c4_rr2 + t2_r4_c4_rr3;

  assign t4_r4_c4_rr0 = t3_r4_c4_rr0 + t3_r4_c4_rr1;

  assign c_4_4 = t4_r4_c4_rr0;
  assign t0_r4_c5_rr0 = a_4_0 * b_0_5;
  assign t0_r4_c5_rr1 = a_4_1 * b_1_5;
  assign t0_r4_c5_rr2 = a_4_2 * b_2_5;
  assign t0_r4_c5_rr3 = a_4_3 * b_3_5;
  assign t0_r4_c5_rr4 = a_4_4 * b_4_5;
  assign t0_r4_c5_rr5 = a_4_5 * b_5_5;
  assign t0_r4_c5_rr6 = a_4_6 * b_6_5;
  assign t0_r4_c5_rr7 = a_4_7 * b_7_5;
  assign t0_r4_c5_rr8 = a_4_8 * b_8_5;
  assign t0_r4_c5_rr9 = a_4_9 * b_9_5;
  assign t0_r4_c5_rr10 = a_4_10 * b_10_5;
  assign t0_r4_c5_rr11 = a_4_11 * b_11_5;
  assign t0_r4_c5_rr12 = a_4_12 * b_12_5;
  assign t0_r4_c5_rr13 = a_4_13 * b_13_5;
  assign t0_r4_c5_rr14 = a_4_14 * b_14_5;
  assign t1_r4_c5_rr0 = t0_r4_c5_rr0 + t0_r4_c5_rr1;
  assign t1_r4_c5_rr1 = t0_r4_c5_rr2 + t0_r4_c5_rr3;
  assign t1_r4_c5_rr2 = t0_r4_c5_rr4 + t0_r4_c5_rr5;
  assign t1_r4_c5_rr3 = t0_r4_c5_rr6 + t0_r4_c5_rr7;
  assign t1_r4_c5_rr4 = t0_r4_c5_rr8 + t0_r4_c5_rr9;
  assign t1_r4_c5_rr5 = t0_r4_c5_rr10 + t0_r4_c5_rr11;
  assign t1_r4_c5_rr6 = t0_r4_c5_rr12 + t0_r4_c5_rr13;
  assign t1_r4_c5_rr7 = t0_r4_c5_rr14;

  assign t2_r4_c5_rr0 = t1_r4_c5_rr0 + t1_r4_c5_rr1;
  assign t2_r4_c5_rr1 = t1_r4_c5_rr2 + t1_r4_c5_rr3;
  assign t2_r4_c5_rr2 = t1_r4_c5_rr4 + t1_r4_c5_rr5;
  assign t2_r4_c5_rr3 = t1_r4_c5_rr6 + t1_r4_c5_rr7;

  assign t3_r4_c5_rr0 = t2_r4_c5_rr0 + t2_r4_c5_rr1;
  assign t3_r4_c5_rr1 = t2_r4_c5_rr2 + t2_r4_c5_rr3;

  assign t4_r4_c5_rr0 = t3_r4_c5_rr0 + t3_r4_c5_rr1;

  assign c_4_5 = t4_r4_c5_rr0;
  assign t0_r4_c6_rr0 = a_4_0 * b_0_6;
  assign t0_r4_c6_rr1 = a_4_1 * b_1_6;
  assign t0_r4_c6_rr2 = a_4_2 * b_2_6;
  assign t0_r4_c6_rr3 = a_4_3 * b_3_6;
  assign t0_r4_c6_rr4 = a_4_4 * b_4_6;
  assign t0_r4_c6_rr5 = a_4_5 * b_5_6;
  assign t0_r4_c6_rr6 = a_4_6 * b_6_6;
  assign t0_r4_c6_rr7 = a_4_7 * b_7_6;
  assign t0_r4_c6_rr8 = a_4_8 * b_8_6;
  assign t0_r4_c6_rr9 = a_4_9 * b_9_6;
  assign t0_r4_c6_rr10 = a_4_10 * b_10_6;
  assign t0_r4_c6_rr11 = a_4_11 * b_11_6;
  assign t0_r4_c6_rr12 = a_4_12 * b_12_6;
  assign t0_r4_c6_rr13 = a_4_13 * b_13_6;
  assign t0_r4_c6_rr14 = a_4_14 * b_14_6;
  assign t1_r4_c6_rr0 = t0_r4_c6_rr0 + t0_r4_c6_rr1;
  assign t1_r4_c6_rr1 = t0_r4_c6_rr2 + t0_r4_c6_rr3;
  assign t1_r4_c6_rr2 = t0_r4_c6_rr4 + t0_r4_c6_rr5;
  assign t1_r4_c6_rr3 = t0_r4_c6_rr6 + t0_r4_c6_rr7;
  assign t1_r4_c6_rr4 = t0_r4_c6_rr8 + t0_r4_c6_rr9;
  assign t1_r4_c6_rr5 = t0_r4_c6_rr10 + t0_r4_c6_rr11;
  assign t1_r4_c6_rr6 = t0_r4_c6_rr12 + t0_r4_c6_rr13;
  assign t1_r4_c6_rr7 = t0_r4_c6_rr14;

  assign t2_r4_c6_rr0 = t1_r4_c6_rr0 + t1_r4_c6_rr1;
  assign t2_r4_c6_rr1 = t1_r4_c6_rr2 + t1_r4_c6_rr3;
  assign t2_r4_c6_rr2 = t1_r4_c6_rr4 + t1_r4_c6_rr5;
  assign t2_r4_c6_rr3 = t1_r4_c6_rr6 + t1_r4_c6_rr7;

  assign t3_r4_c6_rr0 = t2_r4_c6_rr0 + t2_r4_c6_rr1;
  assign t3_r4_c6_rr1 = t2_r4_c6_rr2 + t2_r4_c6_rr3;

  assign t4_r4_c6_rr0 = t3_r4_c6_rr0 + t3_r4_c6_rr1;

  assign c_4_6 = t4_r4_c6_rr0;
  assign t0_r4_c7_rr0 = a_4_0 * b_0_7;
  assign t0_r4_c7_rr1 = a_4_1 * b_1_7;
  assign t0_r4_c7_rr2 = a_4_2 * b_2_7;
  assign t0_r4_c7_rr3 = a_4_3 * b_3_7;
  assign t0_r4_c7_rr4 = a_4_4 * b_4_7;
  assign t0_r4_c7_rr5 = a_4_5 * b_5_7;
  assign t0_r4_c7_rr6 = a_4_6 * b_6_7;
  assign t0_r4_c7_rr7 = a_4_7 * b_7_7;
  assign t0_r4_c7_rr8 = a_4_8 * b_8_7;
  assign t0_r4_c7_rr9 = a_4_9 * b_9_7;
  assign t0_r4_c7_rr10 = a_4_10 * b_10_7;
  assign t0_r4_c7_rr11 = a_4_11 * b_11_7;
  assign t0_r4_c7_rr12 = a_4_12 * b_12_7;
  assign t0_r4_c7_rr13 = a_4_13 * b_13_7;
  assign t0_r4_c7_rr14 = a_4_14 * b_14_7;
  assign t1_r4_c7_rr0 = t0_r4_c7_rr0 + t0_r4_c7_rr1;
  assign t1_r4_c7_rr1 = t0_r4_c7_rr2 + t0_r4_c7_rr3;
  assign t1_r4_c7_rr2 = t0_r4_c7_rr4 + t0_r4_c7_rr5;
  assign t1_r4_c7_rr3 = t0_r4_c7_rr6 + t0_r4_c7_rr7;
  assign t1_r4_c7_rr4 = t0_r4_c7_rr8 + t0_r4_c7_rr9;
  assign t1_r4_c7_rr5 = t0_r4_c7_rr10 + t0_r4_c7_rr11;
  assign t1_r4_c7_rr6 = t0_r4_c7_rr12 + t0_r4_c7_rr13;
  assign t1_r4_c7_rr7 = t0_r4_c7_rr14;

  assign t2_r4_c7_rr0 = t1_r4_c7_rr0 + t1_r4_c7_rr1;
  assign t2_r4_c7_rr1 = t1_r4_c7_rr2 + t1_r4_c7_rr3;
  assign t2_r4_c7_rr2 = t1_r4_c7_rr4 + t1_r4_c7_rr5;
  assign t2_r4_c7_rr3 = t1_r4_c7_rr6 + t1_r4_c7_rr7;

  assign t3_r4_c7_rr0 = t2_r4_c7_rr0 + t2_r4_c7_rr1;
  assign t3_r4_c7_rr1 = t2_r4_c7_rr2 + t2_r4_c7_rr3;

  assign t4_r4_c7_rr0 = t3_r4_c7_rr0 + t3_r4_c7_rr1;

  assign c_4_7 = t4_r4_c7_rr0;
  assign t0_r4_c8_rr0 = a_4_0 * b_0_8;
  assign t0_r4_c8_rr1 = a_4_1 * b_1_8;
  assign t0_r4_c8_rr2 = a_4_2 * b_2_8;
  assign t0_r4_c8_rr3 = a_4_3 * b_3_8;
  assign t0_r4_c8_rr4 = a_4_4 * b_4_8;
  assign t0_r4_c8_rr5 = a_4_5 * b_5_8;
  assign t0_r4_c8_rr6 = a_4_6 * b_6_8;
  assign t0_r4_c8_rr7 = a_4_7 * b_7_8;
  assign t0_r4_c8_rr8 = a_4_8 * b_8_8;
  assign t0_r4_c8_rr9 = a_4_9 * b_9_8;
  assign t0_r4_c8_rr10 = a_4_10 * b_10_8;
  assign t0_r4_c8_rr11 = a_4_11 * b_11_8;
  assign t0_r4_c8_rr12 = a_4_12 * b_12_8;
  assign t0_r4_c8_rr13 = a_4_13 * b_13_8;
  assign t0_r4_c8_rr14 = a_4_14 * b_14_8;
  assign t1_r4_c8_rr0 = t0_r4_c8_rr0 + t0_r4_c8_rr1;
  assign t1_r4_c8_rr1 = t0_r4_c8_rr2 + t0_r4_c8_rr3;
  assign t1_r4_c8_rr2 = t0_r4_c8_rr4 + t0_r4_c8_rr5;
  assign t1_r4_c8_rr3 = t0_r4_c8_rr6 + t0_r4_c8_rr7;
  assign t1_r4_c8_rr4 = t0_r4_c8_rr8 + t0_r4_c8_rr9;
  assign t1_r4_c8_rr5 = t0_r4_c8_rr10 + t0_r4_c8_rr11;
  assign t1_r4_c8_rr6 = t0_r4_c8_rr12 + t0_r4_c8_rr13;
  assign t1_r4_c8_rr7 = t0_r4_c8_rr14;

  assign t2_r4_c8_rr0 = t1_r4_c8_rr0 + t1_r4_c8_rr1;
  assign t2_r4_c8_rr1 = t1_r4_c8_rr2 + t1_r4_c8_rr3;
  assign t2_r4_c8_rr2 = t1_r4_c8_rr4 + t1_r4_c8_rr5;
  assign t2_r4_c8_rr3 = t1_r4_c8_rr6 + t1_r4_c8_rr7;

  assign t3_r4_c8_rr0 = t2_r4_c8_rr0 + t2_r4_c8_rr1;
  assign t3_r4_c8_rr1 = t2_r4_c8_rr2 + t2_r4_c8_rr3;

  assign t4_r4_c8_rr0 = t3_r4_c8_rr0 + t3_r4_c8_rr1;

  assign c_4_8 = t4_r4_c8_rr0;
  assign t0_r4_c9_rr0 = a_4_0 * b_0_9;
  assign t0_r4_c9_rr1 = a_4_1 * b_1_9;
  assign t0_r4_c9_rr2 = a_4_2 * b_2_9;
  assign t0_r4_c9_rr3 = a_4_3 * b_3_9;
  assign t0_r4_c9_rr4 = a_4_4 * b_4_9;
  assign t0_r4_c9_rr5 = a_4_5 * b_5_9;
  assign t0_r4_c9_rr6 = a_4_6 * b_6_9;
  assign t0_r4_c9_rr7 = a_4_7 * b_7_9;
  assign t0_r4_c9_rr8 = a_4_8 * b_8_9;
  assign t0_r4_c9_rr9 = a_4_9 * b_9_9;
  assign t0_r4_c9_rr10 = a_4_10 * b_10_9;
  assign t0_r4_c9_rr11 = a_4_11 * b_11_9;
  assign t0_r4_c9_rr12 = a_4_12 * b_12_9;
  assign t0_r4_c9_rr13 = a_4_13 * b_13_9;
  assign t0_r4_c9_rr14 = a_4_14 * b_14_9;
  assign t1_r4_c9_rr0 = t0_r4_c9_rr0 + t0_r4_c9_rr1;
  assign t1_r4_c9_rr1 = t0_r4_c9_rr2 + t0_r4_c9_rr3;
  assign t1_r4_c9_rr2 = t0_r4_c9_rr4 + t0_r4_c9_rr5;
  assign t1_r4_c9_rr3 = t0_r4_c9_rr6 + t0_r4_c9_rr7;
  assign t1_r4_c9_rr4 = t0_r4_c9_rr8 + t0_r4_c9_rr9;
  assign t1_r4_c9_rr5 = t0_r4_c9_rr10 + t0_r4_c9_rr11;
  assign t1_r4_c9_rr6 = t0_r4_c9_rr12 + t0_r4_c9_rr13;
  assign t1_r4_c9_rr7 = t0_r4_c9_rr14;

  assign t2_r4_c9_rr0 = t1_r4_c9_rr0 + t1_r4_c9_rr1;
  assign t2_r4_c9_rr1 = t1_r4_c9_rr2 + t1_r4_c9_rr3;
  assign t2_r4_c9_rr2 = t1_r4_c9_rr4 + t1_r4_c9_rr5;
  assign t2_r4_c9_rr3 = t1_r4_c9_rr6 + t1_r4_c9_rr7;

  assign t3_r4_c9_rr0 = t2_r4_c9_rr0 + t2_r4_c9_rr1;
  assign t3_r4_c9_rr1 = t2_r4_c9_rr2 + t2_r4_c9_rr3;

  assign t4_r4_c9_rr0 = t3_r4_c9_rr0 + t3_r4_c9_rr1;

  assign c_4_9 = t4_r4_c9_rr0;
  assign t0_r4_c10_rr0 = a_4_0 * b_0_10;
  assign t0_r4_c10_rr1 = a_4_1 * b_1_10;
  assign t0_r4_c10_rr2 = a_4_2 * b_2_10;
  assign t0_r4_c10_rr3 = a_4_3 * b_3_10;
  assign t0_r4_c10_rr4 = a_4_4 * b_4_10;
  assign t0_r4_c10_rr5 = a_4_5 * b_5_10;
  assign t0_r4_c10_rr6 = a_4_6 * b_6_10;
  assign t0_r4_c10_rr7 = a_4_7 * b_7_10;
  assign t0_r4_c10_rr8 = a_4_8 * b_8_10;
  assign t0_r4_c10_rr9 = a_4_9 * b_9_10;
  assign t0_r4_c10_rr10 = a_4_10 * b_10_10;
  assign t0_r4_c10_rr11 = a_4_11 * b_11_10;
  assign t0_r4_c10_rr12 = a_4_12 * b_12_10;
  assign t0_r4_c10_rr13 = a_4_13 * b_13_10;
  assign t0_r4_c10_rr14 = a_4_14 * b_14_10;
  assign t1_r4_c10_rr0 = t0_r4_c10_rr0 + t0_r4_c10_rr1;
  assign t1_r4_c10_rr1 = t0_r4_c10_rr2 + t0_r4_c10_rr3;
  assign t1_r4_c10_rr2 = t0_r4_c10_rr4 + t0_r4_c10_rr5;
  assign t1_r4_c10_rr3 = t0_r4_c10_rr6 + t0_r4_c10_rr7;
  assign t1_r4_c10_rr4 = t0_r4_c10_rr8 + t0_r4_c10_rr9;
  assign t1_r4_c10_rr5 = t0_r4_c10_rr10 + t0_r4_c10_rr11;
  assign t1_r4_c10_rr6 = t0_r4_c10_rr12 + t0_r4_c10_rr13;
  assign t1_r4_c10_rr7 = t0_r4_c10_rr14;

  assign t2_r4_c10_rr0 = t1_r4_c10_rr0 + t1_r4_c10_rr1;
  assign t2_r4_c10_rr1 = t1_r4_c10_rr2 + t1_r4_c10_rr3;
  assign t2_r4_c10_rr2 = t1_r4_c10_rr4 + t1_r4_c10_rr5;
  assign t2_r4_c10_rr3 = t1_r4_c10_rr6 + t1_r4_c10_rr7;

  assign t3_r4_c10_rr0 = t2_r4_c10_rr0 + t2_r4_c10_rr1;
  assign t3_r4_c10_rr1 = t2_r4_c10_rr2 + t2_r4_c10_rr3;

  assign t4_r4_c10_rr0 = t3_r4_c10_rr0 + t3_r4_c10_rr1;

  assign c_4_10 = t4_r4_c10_rr0;
  assign t0_r4_c11_rr0 = a_4_0 * b_0_11;
  assign t0_r4_c11_rr1 = a_4_1 * b_1_11;
  assign t0_r4_c11_rr2 = a_4_2 * b_2_11;
  assign t0_r4_c11_rr3 = a_4_3 * b_3_11;
  assign t0_r4_c11_rr4 = a_4_4 * b_4_11;
  assign t0_r4_c11_rr5 = a_4_5 * b_5_11;
  assign t0_r4_c11_rr6 = a_4_6 * b_6_11;
  assign t0_r4_c11_rr7 = a_4_7 * b_7_11;
  assign t0_r4_c11_rr8 = a_4_8 * b_8_11;
  assign t0_r4_c11_rr9 = a_4_9 * b_9_11;
  assign t0_r4_c11_rr10 = a_4_10 * b_10_11;
  assign t0_r4_c11_rr11 = a_4_11 * b_11_11;
  assign t0_r4_c11_rr12 = a_4_12 * b_12_11;
  assign t0_r4_c11_rr13 = a_4_13 * b_13_11;
  assign t0_r4_c11_rr14 = a_4_14 * b_14_11;
  assign t1_r4_c11_rr0 = t0_r4_c11_rr0 + t0_r4_c11_rr1;
  assign t1_r4_c11_rr1 = t0_r4_c11_rr2 + t0_r4_c11_rr3;
  assign t1_r4_c11_rr2 = t0_r4_c11_rr4 + t0_r4_c11_rr5;
  assign t1_r4_c11_rr3 = t0_r4_c11_rr6 + t0_r4_c11_rr7;
  assign t1_r4_c11_rr4 = t0_r4_c11_rr8 + t0_r4_c11_rr9;
  assign t1_r4_c11_rr5 = t0_r4_c11_rr10 + t0_r4_c11_rr11;
  assign t1_r4_c11_rr6 = t0_r4_c11_rr12 + t0_r4_c11_rr13;
  assign t1_r4_c11_rr7 = t0_r4_c11_rr14;

  assign t2_r4_c11_rr0 = t1_r4_c11_rr0 + t1_r4_c11_rr1;
  assign t2_r4_c11_rr1 = t1_r4_c11_rr2 + t1_r4_c11_rr3;
  assign t2_r4_c11_rr2 = t1_r4_c11_rr4 + t1_r4_c11_rr5;
  assign t2_r4_c11_rr3 = t1_r4_c11_rr6 + t1_r4_c11_rr7;

  assign t3_r4_c11_rr0 = t2_r4_c11_rr0 + t2_r4_c11_rr1;
  assign t3_r4_c11_rr1 = t2_r4_c11_rr2 + t2_r4_c11_rr3;

  assign t4_r4_c11_rr0 = t3_r4_c11_rr0 + t3_r4_c11_rr1;

  assign c_4_11 = t4_r4_c11_rr0;
  assign t0_r4_c12_rr0 = a_4_0 * b_0_12;
  assign t0_r4_c12_rr1 = a_4_1 * b_1_12;
  assign t0_r4_c12_rr2 = a_4_2 * b_2_12;
  assign t0_r4_c12_rr3 = a_4_3 * b_3_12;
  assign t0_r4_c12_rr4 = a_4_4 * b_4_12;
  assign t0_r4_c12_rr5 = a_4_5 * b_5_12;
  assign t0_r4_c12_rr6 = a_4_6 * b_6_12;
  assign t0_r4_c12_rr7 = a_4_7 * b_7_12;
  assign t0_r4_c12_rr8 = a_4_8 * b_8_12;
  assign t0_r4_c12_rr9 = a_4_9 * b_9_12;
  assign t0_r4_c12_rr10 = a_4_10 * b_10_12;
  assign t0_r4_c12_rr11 = a_4_11 * b_11_12;
  assign t0_r4_c12_rr12 = a_4_12 * b_12_12;
  assign t0_r4_c12_rr13 = a_4_13 * b_13_12;
  assign t0_r4_c12_rr14 = a_4_14 * b_14_12;
  assign t1_r4_c12_rr0 = t0_r4_c12_rr0 + t0_r4_c12_rr1;
  assign t1_r4_c12_rr1 = t0_r4_c12_rr2 + t0_r4_c12_rr3;
  assign t1_r4_c12_rr2 = t0_r4_c12_rr4 + t0_r4_c12_rr5;
  assign t1_r4_c12_rr3 = t0_r4_c12_rr6 + t0_r4_c12_rr7;
  assign t1_r4_c12_rr4 = t0_r4_c12_rr8 + t0_r4_c12_rr9;
  assign t1_r4_c12_rr5 = t0_r4_c12_rr10 + t0_r4_c12_rr11;
  assign t1_r4_c12_rr6 = t0_r4_c12_rr12 + t0_r4_c12_rr13;
  assign t1_r4_c12_rr7 = t0_r4_c12_rr14;

  assign t2_r4_c12_rr0 = t1_r4_c12_rr0 + t1_r4_c12_rr1;
  assign t2_r4_c12_rr1 = t1_r4_c12_rr2 + t1_r4_c12_rr3;
  assign t2_r4_c12_rr2 = t1_r4_c12_rr4 + t1_r4_c12_rr5;
  assign t2_r4_c12_rr3 = t1_r4_c12_rr6 + t1_r4_c12_rr7;

  assign t3_r4_c12_rr0 = t2_r4_c12_rr0 + t2_r4_c12_rr1;
  assign t3_r4_c12_rr1 = t2_r4_c12_rr2 + t2_r4_c12_rr3;

  assign t4_r4_c12_rr0 = t3_r4_c12_rr0 + t3_r4_c12_rr1;

  assign c_4_12 = t4_r4_c12_rr0;
  assign t0_r4_c13_rr0 = a_4_0 * b_0_13;
  assign t0_r4_c13_rr1 = a_4_1 * b_1_13;
  assign t0_r4_c13_rr2 = a_4_2 * b_2_13;
  assign t0_r4_c13_rr3 = a_4_3 * b_3_13;
  assign t0_r4_c13_rr4 = a_4_4 * b_4_13;
  assign t0_r4_c13_rr5 = a_4_5 * b_5_13;
  assign t0_r4_c13_rr6 = a_4_6 * b_6_13;
  assign t0_r4_c13_rr7 = a_4_7 * b_7_13;
  assign t0_r4_c13_rr8 = a_4_8 * b_8_13;
  assign t0_r4_c13_rr9 = a_4_9 * b_9_13;
  assign t0_r4_c13_rr10 = a_4_10 * b_10_13;
  assign t0_r4_c13_rr11 = a_4_11 * b_11_13;
  assign t0_r4_c13_rr12 = a_4_12 * b_12_13;
  assign t0_r4_c13_rr13 = a_4_13 * b_13_13;
  assign t0_r4_c13_rr14 = a_4_14 * b_14_13;
  assign t1_r4_c13_rr0 = t0_r4_c13_rr0 + t0_r4_c13_rr1;
  assign t1_r4_c13_rr1 = t0_r4_c13_rr2 + t0_r4_c13_rr3;
  assign t1_r4_c13_rr2 = t0_r4_c13_rr4 + t0_r4_c13_rr5;
  assign t1_r4_c13_rr3 = t0_r4_c13_rr6 + t0_r4_c13_rr7;
  assign t1_r4_c13_rr4 = t0_r4_c13_rr8 + t0_r4_c13_rr9;
  assign t1_r4_c13_rr5 = t0_r4_c13_rr10 + t0_r4_c13_rr11;
  assign t1_r4_c13_rr6 = t0_r4_c13_rr12 + t0_r4_c13_rr13;
  assign t1_r4_c13_rr7 = t0_r4_c13_rr14;

  assign t2_r4_c13_rr0 = t1_r4_c13_rr0 + t1_r4_c13_rr1;
  assign t2_r4_c13_rr1 = t1_r4_c13_rr2 + t1_r4_c13_rr3;
  assign t2_r4_c13_rr2 = t1_r4_c13_rr4 + t1_r4_c13_rr5;
  assign t2_r4_c13_rr3 = t1_r4_c13_rr6 + t1_r4_c13_rr7;

  assign t3_r4_c13_rr0 = t2_r4_c13_rr0 + t2_r4_c13_rr1;
  assign t3_r4_c13_rr1 = t2_r4_c13_rr2 + t2_r4_c13_rr3;

  assign t4_r4_c13_rr0 = t3_r4_c13_rr0 + t3_r4_c13_rr1;

  assign c_4_13 = t4_r4_c13_rr0;
  assign t0_r4_c14_rr0 = a_4_0 * b_0_14;
  assign t0_r4_c14_rr1 = a_4_1 * b_1_14;
  assign t0_r4_c14_rr2 = a_4_2 * b_2_14;
  assign t0_r4_c14_rr3 = a_4_3 * b_3_14;
  assign t0_r4_c14_rr4 = a_4_4 * b_4_14;
  assign t0_r4_c14_rr5 = a_4_5 * b_5_14;
  assign t0_r4_c14_rr6 = a_4_6 * b_6_14;
  assign t0_r4_c14_rr7 = a_4_7 * b_7_14;
  assign t0_r4_c14_rr8 = a_4_8 * b_8_14;
  assign t0_r4_c14_rr9 = a_4_9 * b_9_14;
  assign t0_r4_c14_rr10 = a_4_10 * b_10_14;
  assign t0_r4_c14_rr11 = a_4_11 * b_11_14;
  assign t0_r4_c14_rr12 = a_4_12 * b_12_14;
  assign t0_r4_c14_rr13 = a_4_13 * b_13_14;
  assign t0_r4_c14_rr14 = a_4_14 * b_14_14;
  assign t1_r4_c14_rr0 = t0_r4_c14_rr0 + t0_r4_c14_rr1;
  assign t1_r4_c14_rr1 = t0_r4_c14_rr2 + t0_r4_c14_rr3;
  assign t1_r4_c14_rr2 = t0_r4_c14_rr4 + t0_r4_c14_rr5;
  assign t1_r4_c14_rr3 = t0_r4_c14_rr6 + t0_r4_c14_rr7;
  assign t1_r4_c14_rr4 = t0_r4_c14_rr8 + t0_r4_c14_rr9;
  assign t1_r4_c14_rr5 = t0_r4_c14_rr10 + t0_r4_c14_rr11;
  assign t1_r4_c14_rr6 = t0_r4_c14_rr12 + t0_r4_c14_rr13;
  assign t1_r4_c14_rr7 = t0_r4_c14_rr14;

  assign t2_r4_c14_rr0 = t1_r4_c14_rr0 + t1_r4_c14_rr1;
  assign t2_r4_c14_rr1 = t1_r4_c14_rr2 + t1_r4_c14_rr3;
  assign t2_r4_c14_rr2 = t1_r4_c14_rr4 + t1_r4_c14_rr5;
  assign t2_r4_c14_rr3 = t1_r4_c14_rr6 + t1_r4_c14_rr7;

  assign t3_r4_c14_rr0 = t2_r4_c14_rr0 + t2_r4_c14_rr1;
  assign t3_r4_c14_rr1 = t2_r4_c14_rr2 + t2_r4_c14_rr3;

  assign t4_r4_c14_rr0 = t3_r4_c14_rr0 + t3_r4_c14_rr1;

  assign c_4_14 = t4_r4_c14_rr0;
  assign t0_r5_c0_rr0 = a_5_0 * b_0_0;
  assign t0_r5_c0_rr1 = a_5_1 * b_1_0;
  assign t0_r5_c0_rr2 = a_5_2 * b_2_0;
  assign t0_r5_c0_rr3 = a_5_3 * b_3_0;
  assign t0_r5_c0_rr4 = a_5_4 * b_4_0;
  assign t0_r5_c0_rr5 = a_5_5 * b_5_0;
  assign t0_r5_c0_rr6 = a_5_6 * b_6_0;
  assign t0_r5_c0_rr7 = a_5_7 * b_7_0;
  assign t0_r5_c0_rr8 = a_5_8 * b_8_0;
  assign t0_r5_c0_rr9 = a_5_9 * b_9_0;
  assign t0_r5_c0_rr10 = a_5_10 * b_10_0;
  assign t0_r5_c0_rr11 = a_5_11 * b_11_0;
  assign t0_r5_c0_rr12 = a_5_12 * b_12_0;
  assign t0_r5_c0_rr13 = a_5_13 * b_13_0;
  assign t0_r5_c0_rr14 = a_5_14 * b_14_0;
  assign t1_r5_c0_rr0 = t0_r5_c0_rr0 + t0_r5_c0_rr1;
  assign t1_r5_c0_rr1 = t0_r5_c0_rr2 + t0_r5_c0_rr3;
  assign t1_r5_c0_rr2 = t0_r5_c0_rr4 + t0_r5_c0_rr5;
  assign t1_r5_c0_rr3 = t0_r5_c0_rr6 + t0_r5_c0_rr7;
  assign t1_r5_c0_rr4 = t0_r5_c0_rr8 + t0_r5_c0_rr9;
  assign t1_r5_c0_rr5 = t0_r5_c0_rr10 + t0_r5_c0_rr11;
  assign t1_r5_c0_rr6 = t0_r5_c0_rr12 + t0_r5_c0_rr13;
  assign t1_r5_c0_rr7 = t0_r5_c0_rr14;

  assign t2_r5_c0_rr0 = t1_r5_c0_rr0 + t1_r5_c0_rr1;
  assign t2_r5_c0_rr1 = t1_r5_c0_rr2 + t1_r5_c0_rr3;
  assign t2_r5_c0_rr2 = t1_r5_c0_rr4 + t1_r5_c0_rr5;
  assign t2_r5_c0_rr3 = t1_r5_c0_rr6 + t1_r5_c0_rr7;

  assign t3_r5_c0_rr0 = t2_r5_c0_rr0 + t2_r5_c0_rr1;
  assign t3_r5_c0_rr1 = t2_r5_c0_rr2 + t2_r5_c0_rr3;

  assign t4_r5_c0_rr0 = t3_r5_c0_rr0 + t3_r5_c0_rr1;

  assign c_5_0 = t4_r5_c0_rr0;
  assign t0_r5_c1_rr0 = a_5_0 * b_0_1;
  assign t0_r5_c1_rr1 = a_5_1 * b_1_1;
  assign t0_r5_c1_rr2 = a_5_2 * b_2_1;
  assign t0_r5_c1_rr3 = a_5_3 * b_3_1;
  assign t0_r5_c1_rr4 = a_5_4 * b_4_1;
  assign t0_r5_c1_rr5 = a_5_5 * b_5_1;
  assign t0_r5_c1_rr6 = a_5_6 * b_6_1;
  assign t0_r5_c1_rr7 = a_5_7 * b_7_1;
  assign t0_r5_c1_rr8 = a_5_8 * b_8_1;
  assign t0_r5_c1_rr9 = a_5_9 * b_9_1;
  assign t0_r5_c1_rr10 = a_5_10 * b_10_1;
  assign t0_r5_c1_rr11 = a_5_11 * b_11_1;
  assign t0_r5_c1_rr12 = a_5_12 * b_12_1;
  assign t0_r5_c1_rr13 = a_5_13 * b_13_1;
  assign t0_r5_c1_rr14 = a_5_14 * b_14_1;
  assign t1_r5_c1_rr0 = t0_r5_c1_rr0 + t0_r5_c1_rr1;
  assign t1_r5_c1_rr1 = t0_r5_c1_rr2 + t0_r5_c1_rr3;
  assign t1_r5_c1_rr2 = t0_r5_c1_rr4 + t0_r5_c1_rr5;
  assign t1_r5_c1_rr3 = t0_r5_c1_rr6 + t0_r5_c1_rr7;
  assign t1_r5_c1_rr4 = t0_r5_c1_rr8 + t0_r5_c1_rr9;
  assign t1_r5_c1_rr5 = t0_r5_c1_rr10 + t0_r5_c1_rr11;
  assign t1_r5_c1_rr6 = t0_r5_c1_rr12 + t0_r5_c1_rr13;
  assign t1_r5_c1_rr7 = t0_r5_c1_rr14;

  assign t2_r5_c1_rr0 = t1_r5_c1_rr0 + t1_r5_c1_rr1;
  assign t2_r5_c1_rr1 = t1_r5_c1_rr2 + t1_r5_c1_rr3;
  assign t2_r5_c1_rr2 = t1_r5_c1_rr4 + t1_r5_c1_rr5;
  assign t2_r5_c1_rr3 = t1_r5_c1_rr6 + t1_r5_c1_rr7;

  assign t3_r5_c1_rr0 = t2_r5_c1_rr0 + t2_r5_c1_rr1;
  assign t3_r5_c1_rr1 = t2_r5_c1_rr2 + t2_r5_c1_rr3;

  assign t4_r5_c1_rr0 = t3_r5_c1_rr0 + t3_r5_c1_rr1;

  assign c_5_1 = t4_r5_c1_rr0;
  assign t0_r5_c2_rr0 = a_5_0 * b_0_2;
  assign t0_r5_c2_rr1 = a_5_1 * b_1_2;
  assign t0_r5_c2_rr2 = a_5_2 * b_2_2;
  assign t0_r5_c2_rr3 = a_5_3 * b_3_2;
  assign t0_r5_c2_rr4 = a_5_4 * b_4_2;
  assign t0_r5_c2_rr5 = a_5_5 * b_5_2;
  assign t0_r5_c2_rr6 = a_5_6 * b_6_2;
  assign t0_r5_c2_rr7 = a_5_7 * b_7_2;
  assign t0_r5_c2_rr8 = a_5_8 * b_8_2;
  assign t0_r5_c2_rr9 = a_5_9 * b_9_2;
  assign t0_r5_c2_rr10 = a_5_10 * b_10_2;
  assign t0_r5_c2_rr11 = a_5_11 * b_11_2;
  assign t0_r5_c2_rr12 = a_5_12 * b_12_2;
  assign t0_r5_c2_rr13 = a_5_13 * b_13_2;
  assign t0_r5_c2_rr14 = a_5_14 * b_14_2;
  assign t1_r5_c2_rr0 = t0_r5_c2_rr0 + t0_r5_c2_rr1;
  assign t1_r5_c2_rr1 = t0_r5_c2_rr2 + t0_r5_c2_rr3;
  assign t1_r5_c2_rr2 = t0_r5_c2_rr4 + t0_r5_c2_rr5;
  assign t1_r5_c2_rr3 = t0_r5_c2_rr6 + t0_r5_c2_rr7;
  assign t1_r5_c2_rr4 = t0_r5_c2_rr8 + t0_r5_c2_rr9;
  assign t1_r5_c2_rr5 = t0_r5_c2_rr10 + t0_r5_c2_rr11;
  assign t1_r5_c2_rr6 = t0_r5_c2_rr12 + t0_r5_c2_rr13;
  assign t1_r5_c2_rr7 = t0_r5_c2_rr14;

  assign t2_r5_c2_rr0 = t1_r5_c2_rr0 + t1_r5_c2_rr1;
  assign t2_r5_c2_rr1 = t1_r5_c2_rr2 + t1_r5_c2_rr3;
  assign t2_r5_c2_rr2 = t1_r5_c2_rr4 + t1_r5_c2_rr5;
  assign t2_r5_c2_rr3 = t1_r5_c2_rr6 + t1_r5_c2_rr7;

  assign t3_r5_c2_rr0 = t2_r5_c2_rr0 + t2_r5_c2_rr1;
  assign t3_r5_c2_rr1 = t2_r5_c2_rr2 + t2_r5_c2_rr3;

  assign t4_r5_c2_rr0 = t3_r5_c2_rr0 + t3_r5_c2_rr1;

  assign c_5_2 = t4_r5_c2_rr0;
  assign t0_r5_c3_rr0 = a_5_0 * b_0_3;
  assign t0_r5_c3_rr1 = a_5_1 * b_1_3;
  assign t0_r5_c3_rr2 = a_5_2 * b_2_3;
  assign t0_r5_c3_rr3 = a_5_3 * b_3_3;
  assign t0_r5_c3_rr4 = a_5_4 * b_4_3;
  assign t0_r5_c3_rr5 = a_5_5 * b_5_3;
  assign t0_r5_c3_rr6 = a_5_6 * b_6_3;
  assign t0_r5_c3_rr7 = a_5_7 * b_7_3;
  assign t0_r5_c3_rr8 = a_5_8 * b_8_3;
  assign t0_r5_c3_rr9 = a_5_9 * b_9_3;
  assign t0_r5_c3_rr10 = a_5_10 * b_10_3;
  assign t0_r5_c3_rr11 = a_5_11 * b_11_3;
  assign t0_r5_c3_rr12 = a_5_12 * b_12_3;
  assign t0_r5_c3_rr13 = a_5_13 * b_13_3;
  assign t0_r5_c3_rr14 = a_5_14 * b_14_3;
  assign t1_r5_c3_rr0 = t0_r5_c3_rr0 + t0_r5_c3_rr1;
  assign t1_r5_c3_rr1 = t0_r5_c3_rr2 + t0_r5_c3_rr3;
  assign t1_r5_c3_rr2 = t0_r5_c3_rr4 + t0_r5_c3_rr5;
  assign t1_r5_c3_rr3 = t0_r5_c3_rr6 + t0_r5_c3_rr7;
  assign t1_r5_c3_rr4 = t0_r5_c3_rr8 + t0_r5_c3_rr9;
  assign t1_r5_c3_rr5 = t0_r5_c3_rr10 + t0_r5_c3_rr11;
  assign t1_r5_c3_rr6 = t0_r5_c3_rr12 + t0_r5_c3_rr13;
  assign t1_r5_c3_rr7 = t0_r5_c3_rr14;

  assign t2_r5_c3_rr0 = t1_r5_c3_rr0 + t1_r5_c3_rr1;
  assign t2_r5_c3_rr1 = t1_r5_c3_rr2 + t1_r5_c3_rr3;
  assign t2_r5_c3_rr2 = t1_r5_c3_rr4 + t1_r5_c3_rr5;
  assign t2_r5_c3_rr3 = t1_r5_c3_rr6 + t1_r5_c3_rr7;

  assign t3_r5_c3_rr0 = t2_r5_c3_rr0 + t2_r5_c3_rr1;
  assign t3_r5_c3_rr1 = t2_r5_c3_rr2 + t2_r5_c3_rr3;

  assign t4_r5_c3_rr0 = t3_r5_c3_rr0 + t3_r5_c3_rr1;

  assign c_5_3 = t4_r5_c3_rr0;
  assign t0_r5_c4_rr0 = a_5_0 * b_0_4;
  assign t0_r5_c4_rr1 = a_5_1 * b_1_4;
  assign t0_r5_c4_rr2 = a_5_2 * b_2_4;
  assign t0_r5_c4_rr3 = a_5_3 * b_3_4;
  assign t0_r5_c4_rr4 = a_5_4 * b_4_4;
  assign t0_r5_c4_rr5 = a_5_5 * b_5_4;
  assign t0_r5_c4_rr6 = a_5_6 * b_6_4;
  assign t0_r5_c4_rr7 = a_5_7 * b_7_4;
  assign t0_r5_c4_rr8 = a_5_8 * b_8_4;
  assign t0_r5_c4_rr9 = a_5_9 * b_9_4;
  assign t0_r5_c4_rr10 = a_5_10 * b_10_4;
  assign t0_r5_c4_rr11 = a_5_11 * b_11_4;
  assign t0_r5_c4_rr12 = a_5_12 * b_12_4;
  assign t0_r5_c4_rr13 = a_5_13 * b_13_4;
  assign t0_r5_c4_rr14 = a_5_14 * b_14_4;
  assign t1_r5_c4_rr0 = t0_r5_c4_rr0 + t0_r5_c4_rr1;
  assign t1_r5_c4_rr1 = t0_r5_c4_rr2 + t0_r5_c4_rr3;
  assign t1_r5_c4_rr2 = t0_r5_c4_rr4 + t0_r5_c4_rr5;
  assign t1_r5_c4_rr3 = t0_r5_c4_rr6 + t0_r5_c4_rr7;
  assign t1_r5_c4_rr4 = t0_r5_c4_rr8 + t0_r5_c4_rr9;
  assign t1_r5_c4_rr5 = t0_r5_c4_rr10 + t0_r5_c4_rr11;
  assign t1_r5_c4_rr6 = t0_r5_c4_rr12 + t0_r5_c4_rr13;
  assign t1_r5_c4_rr7 = t0_r5_c4_rr14;

  assign t2_r5_c4_rr0 = t1_r5_c4_rr0 + t1_r5_c4_rr1;
  assign t2_r5_c4_rr1 = t1_r5_c4_rr2 + t1_r5_c4_rr3;
  assign t2_r5_c4_rr2 = t1_r5_c4_rr4 + t1_r5_c4_rr5;
  assign t2_r5_c4_rr3 = t1_r5_c4_rr6 + t1_r5_c4_rr7;

  assign t3_r5_c4_rr0 = t2_r5_c4_rr0 + t2_r5_c4_rr1;
  assign t3_r5_c4_rr1 = t2_r5_c4_rr2 + t2_r5_c4_rr3;

  assign t4_r5_c4_rr0 = t3_r5_c4_rr0 + t3_r5_c4_rr1;

  assign c_5_4 = t4_r5_c4_rr0;
  assign t0_r5_c5_rr0 = a_5_0 * b_0_5;
  assign t0_r5_c5_rr1 = a_5_1 * b_1_5;
  assign t0_r5_c5_rr2 = a_5_2 * b_2_5;
  assign t0_r5_c5_rr3 = a_5_3 * b_3_5;
  assign t0_r5_c5_rr4 = a_5_4 * b_4_5;
  assign t0_r5_c5_rr5 = a_5_5 * b_5_5;
  assign t0_r5_c5_rr6 = a_5_6 * b_6_5;
  assign t0_r5_c5_rr7 = a_5_7 * b_7_5;
  assign t0_r5_c5_rr8 = a_5_8 * b_8_5;
  assign t0_r5_c5_rr9 = a_5_9 * b_9_5;
  assign t0_r5_c5_rr10 = a_5_10 * b_10_5;
  assign t0_r5_c5_rr11 = a_5_11 * b_11_5;
  assign t0_r5_c5_rr12 = a_5_12 * b_12_5;
  assign t0_r5_c5_rr13 = a_5_13 * b_13_5;
  assign t0_r5_c5_rr14 = a_5_14 * b_14_5;
  assign t1_r5_c5_rr0 = t0_r5_c5_rr0 + t0_r5_c5_rr1;
  assign t1_r5_c5_rr1 = t0_r5_c5_rr2 + t0_r5_c5_rr3;
  assign t1_r5_c5_rr2 = t0_r5_c5_rr4 + t0_r5_c5_rr5;
  assign t1_r5_c5_rr3 = t0_r5_c5_rr6 + t0_r5_c5_rr7;
  assign t1_r5_c5_rr4 = t0_r5_c5_rr8 + t0_r5_c5_rr9;
  assign t1_r5_c5_rr5 = t0_r5_c5_rr10 + t0_r5_c5_rr11;
  assign t1_r5_c5_rr6 = t0_r5_c5_rr12 + t0_r5_c5_rr13;
  assign t1_r5_c5_rr7 = t0_r5_c5_rr14;

  assign t2_r5_c5_rr0 = t1_r5_c5_rr0 + t1_r5_c5_rr1;
  assign t2_r5_c5_rr1 = t1_r5_c5_rr2 + t1_r5_c5_rr3;
  assign t2_r5_c5_rr2 = t1_r5_c5_rr4 + t1_r5_c5_rr5;
  assign t2_r5_c5_rr3 = t1_r5_c5_rr6 + t1_r5_c5_rr7;

  assign t3_r5_c5_rr0 = t2_r5_c5_rr0 + t2_r5_c5_rr1;
  assign t3_r5_c5_rr1 = t2_r5_c5_rr2 + t2_r5_c5_rr3;

  assign t4_r5_c5_rr0 = t3_r5_c5_rr0 + t3_r5_c5_rr1;

  assign c_5_5 = t4_r5_c5_rr0;
  assign t0_r5_c6_rr0 = a_5_0 * b_0_6;
  assign t0_r5_c6_rr1 = a_5_1 * b_1_6;
  assign t0_r5_c6_rr2 = a_5_2 * b_2_6;
  assign t0_r5_c6_rr3 = a_5_3 * b_3_6;
  assign t0_r5_c6_rr4 = a_5_4 * b_4_6;
  assign t0_r5_c6_rr5 = a_5_5 * b_5_6;
  assign t0_r5_c6_rr6 = a_5_6 * b_6_6;
  assign t0_r5_c6_rr7 = a_5_7 * b_7_6;
  assign t0_r5_c6_rr8 = a_5_8 * b_8_6;
  assign t0_r5_c6_rr9 = a_5_9 * b_9_6;
  assign t0_r5_c6_rr10 = a_5_10 * b_10_6;
  assign t0_r5_c6_rr11 = a_5_11 * b_11_6;
  assign t0_r5_c6_rr12 = a_5_12 * b_12_6;
  assign t0_r5_c6_rr13 = a_5_13 * b_13_6;
  assign t0_r5_c6_rr14 = a_5_14 * b_14_6;
  assign t1_r5_c6_rr0 = t0_r5_c6_rr0 + t0_r5_c6_rr1;
  assign t1_r5_c6_rr1 = t0_r5_c6_rr2 + t0_r5_c6_rr3;
  assign t1_r5_c6_rr2 = t0_r5_c6_rr4 + t0_r5_c6_rr5;
  assign t1_r5_c6_rr3 = t0_r5_c6_rr6 + t0_r5_c6_rr7;
  assign t1_r5_c6_rr4 = t0_r5_c6_rr8 + t0_r5_c6_rr9;
  assign t1_r5_c6_rr5 = t0_r5_c6_rr10 + t0_r5_c6_rr11;
  assign t1_r5_c6_rr6 = t0_r5_c6_rr12 + t0_r5_c6_rr13;
  assign t1_r5_c6_rr7 = t0_r5_c6_rr14;

  assign t2_r5_c6_rr0 = t1_r5_c6_rr0 + t1_r5_c6_rr1;
  assign t2_r5_c6_rr1 = t1_r5_c6_rr2 + t1_r5_c6_rr3;
  assign t2_r5_c6_rr2 = t1_r5_c6_rr4 + t1_r5_c6_rr5;
  assign t2_r5_c6_rr3 = t1_r5_c6_rr6 + t1_r5_c6_rr7;

  assign t3_r5_c6_rr0 = t2_r5_c6_rr0 + t2_r5_c6_rr1;
  assign t3_r5_c6_rr1 = t2_r5_c6_rr2 + t2_r5_c6_rr3;

  assign t4_r5_c6_rr0 = t3_r5_c6_rr0 + t3_r5_c6_rr1;

  assign c_5_6 = t4_r5_c6_rr0;
  assign t0_r5_c7_rr0 = a_5_0 * b_0_7;
  assign t0_r5_c7_rr1 = a_5_1 * b_1_7;
  assign t0_r5_c7_rr2 = a_5_2 * b_2_7;
  assign t0_r5_c7_rr3 = a_5_3 * b_3_7;
  assign t0_r5_c7_rr4 = a_5_4 * b_4_7;
  assign t0_r5_c7_rr5 = a_5_5 * b_5_7;
  assign t0_r5_c7_rr6 = a_5_6 * b_6_7;
  assign t0_r5_c7_rr7 = a_5_7 * b_7_7;
  assign t0_r5_c7_rr8 = a_5_8 * b_8_7;
  assign t0_r5_c7_rr9 = a_5_9 * b_9_7;
  assign t0_r5_c7_rr10 = a_5_10 * b_10_7;
  assign t0_r5_c7_rr11 = a_5_11 * b_11_7;
  assign t0_r5_c7_rr12 = a_5_12 * b_12_7;
  assign t0_r5_c7_rr13 = a_5_13 * b_13_7;
  assign t0_r5_c7_rr14 = a_5_14 * b_14_7;
  assign t1_r5_c7_rr0 = t0_r5_c7_rr0 + t0_r5_c7_rr1;
  assign t1_r5_c7_rr1 = t0_r5_c7_rr2 + t0_r5_c7_rr3;
  assign t1_r5_c7_rr2 = t0_r5_c7_rr4 + t0_r5_c7_rr5;
  assign t1_r5_c7_rr3 = t0_r5_c7_rr6 + t0_r5_c7_rr7;
  assign t1_r5_c7_rr4 = t0_r5_c7_rr8 + t0_r5_c7_rr9;
  assign t1_r5_c7_rr5 = t0_r5_c7_rr10 + t0_r5_c7_rr11;
  assign t1_r5_c7_rr6 = t0_r5_c7_rr12 + t0_r5_c7_rr13;
  assign t1_r5_c7_rr7 = t0_r5_c7_rr14;

  assign t2_r5_c7_rr0 = t1_r5_c7_rr0 + t1_r5_c7_rr1;
  assign t2_r5_c7_rr1 = t1_r5_c7_rr2 + t1_r5_c7_rr3;
  assign t2_r5_c7_rr2 = t1_r5_c7_rr4 + t1_r5_c7_rr5;
  assign t2_r5_c7_rr3 = t1_r5_c7_rr6 + t1_r5_c7_rr7;

  assign t3_r5_c7_rr0 = t2_r5_c7_rr0 + t2_r5_c7_rr1;
  assign t3_r5_c7_rr1 = t2_r5_c7_rr2 + t2_r5_c7_rr3;

  assign t4_r5_c7_rr0 = t3_r5_c7_rr0 + t3_r5_c7_rr1;

  assign c_5_7 = t4_r5_c7_rr0;
  assign t0_r5_c8_rr0 = a_5_0 * b_0_8;
  assign t0_r5_c8_rr1 = a_5_1 * b_1_8;
  assign t0_r5_c8_rr2 = a_5_2 * b_2_8;
  assign t0_r5_c8_rr3 = a_5_3 * b_3_8;
  assign t0_r5_c8_rr4 = a_5_4 * b_4_8;
  assign t0_r5_c8_rr5 = a_5_5 * b_5_8;
  assign t0_r5_c8_rr6 = a_5_6 * b_6_8;
  assign t0_r5_c8_rr7 = a_5_7 * b_7_8;
  assign t0_r5_c8_rr8 = a_5_8 * b_8_8;
  assign t0_r5_c8_rr9 = a_5_9 * b_9_8;
  assign t0_r5_c8_rr10 = a_5_10 * b_10_8;
  assign t0_r5_c8_rr11 = a_5_11 * b_11_8;
  assign t0_r5_c8_rr12 = a_5_12 * b_12_8;
  assign t0_r5_c8_rr13 = a_5_13 * b_13_8;
  assign t0_r5_c8_rr14 = a_5_14 * b_14_8;
  assign t1_r5_c8_rr0 = t0_r5_c8_rr0 + t0_r5_c8_rr1;
  assign t1_r5_c8_rr1 = t0_r5_c8_rr2 + t0_r5_c8_rr3;
  assign t1_r5_c8_rr2 = t0_r5_c8_rr4 + t0_r5_c8_rr5;
  assign t1_r5_c8_rr3 = t0_r5_c8_rr6 + t0_r5_c8_rr7;
  assign t1_r5_c8_rr4 = t0_r5_c8_rr8 + t0_r5_c8_rr9;
  assign t1_r5_c8_rr5 = t0_r5_c8_rr10 + t0_r5_c8_rr11;
  assign t1_r5_c8_rr6 = t0_r5_c8_rr12 + t0_r5_c8_rr13;
  assign t1_r5_c8_rr7 = t0_r5_c8_rr14;

  assign t2_r5_c8_rr0 = t1_r5_c8_rr0 + t1_r5_c8_rr1;
  assign t2_r5_c8_rr1 = t1_r5_c8_rr2 + t1_r5_c8_rr3;
  assign t2_r5_c8_rr2 = t1_r5_c8_rr4 + t1_r5_c8_rr5;
  assign t2_r5_c8_rr3 = t1_r5_c8_rr6 + t1_r5_c8_rr7;

  assign t3_r5_c8_rr0 = t2_r5_c8_rr0 + t2_r5_c8_rr1;
  assign t3_r5_c8_rr1 = t2_r5_c8_rr2 + t2_r5_c8_rr3;

  assign t4_r5_c8_rr0 = t3_r5_c8_rr0 + t3_r5_c8_rr1;

  assign c_5_8 = t4_r5_c8_rr0;
  assign t0_r5_c9_rr0 = a_5_0 * b_0_9;
  assign t0_r5_c9_rr1 = a_5_1 * b_1_9;
  assign t0_r5_c9_rr2 = a_5_2 * b_2_9;
  assign t0_r5_c9_rr3 = a_5_3 * b_3_9;
  assign t0_r5_c9_rr4 = a_5_4 * b_4_9;
  assign t0_r5_c9_rr5 = a_5_5 * b_5_9;
  assign t0_r5_c9_rr6 = a_5_6 * b_6_9;
  assign t0_r5_c9_rr7 = a_5_7 * b_7_9;
  assign t0_r5_c9_rr8 = a_5_8 * b_8_9;
  assign t0_r5_c9_rr9 = a_5_9 * b_9_9;
  assign t0_r5_c9_rr10 = a_5_10 * b_10_9;
  assign t0_r5_c9_rr11 = a_5_11 * b_11_9;
  assign t0_r5_c9_rr12 = a_5_12 * b_12_9;
  assign t0_r5_c9_rr13 = a_5_13 * b_13_9;
  assign t0_r5_c9_rr14 = a_5_14 * b_14_9;
  assign t1_r5_c9_rr0 = t0_r5_c9_rr0 + t0_r5_c9_rr1;
  assign t1_r5_c9_rr1 = t0_r5_c9_rr2 + t0_r5_c9_rr3;
  assign t1_r5_c9_rr2 = t0_r5_c9_rr4 + t0_r5_c9_rr5;
  assign t1_r5_c9_rr3 = t0_r5_c9_rr6 + t0_r5_c9_rr7;
  assign t1_r5_c9_rr4 = t0_r5_c9_rr8 + t0_r5_c9_rr9;
  assign t1_r5_c9_rr5 = t0_r5_c9_rr10 + t0_r5_c9_rr11;
  assign t1_r5_c9_rr6 = t0_r5_c9_rr12 + t0_r5_c9_rr13;
  assign t1_r5_c9_rr7 = t0_r5_c9_rr14;

  assign t2_r5_c9_rr0 = t1_r5_c9_rr0 + t1_r5_c9_rr1;
  assign t2_r5_c9_rr1 = t1_r5_c9_rr2 + t1_r5_c9_rr3;
  assign t2_r5_c9_rr2 = t1_r5_c9_rr4 + t1_r5_c9_rr5;
  assign t2_r5_c9_rr3 = t1_r5_c9_rr6 + t1_r5_c9_rr7;

  assign t3_r5_c9_rr0 = t2_r5_c9_rr0 + t2_r5_c9_rr1;
  assign t3_r5_c9_rr1 = t2_r5_c9_rr2 + t2_r5_c9_rr3;

  assign t4_r5_c9_rr0 = t3_r5_c9_rr0 + t3_r5_c9_rr1;

  assign c_5_9 = t4_r5_c9_rr0;
  assign t0_r5_c10_rr0 = a_5_0 * b_0_10;
  assign t0_r5_c10_rr1 = a_5_1 * b_1_10;
  assign t0_r5_c10_rr2 = a_5_2 * b_2_10;
  assign t0_r5_c10_rr3 = a_5_3 * b_3_10;
  assign t0_r5_c10_rr4 = a_5_4 * b_4_10;
  assign t0_r5_c10_rr5 = a_5_5 * b_5_10;
  assign t0_r5_c10_rr6 = a_5_6 * b_6_10;
  assign t0_r5_c10_rr7 = a_5_7 * b_7_10;
  assign t0_r5_c10_rr8 = a_5_8 * b_8_10;
  assign t0_r5_c10_rr9 = a_5_9 * b_9_10;
  assign t0_r5_c10_rr10 = a_5_10 * b_10_10;
  assign t0_r5_c10_rr11 = a_5_11 * b_11_10;
  assign t0_r5_c10_rr12 = a_5_12 * b_12_10;
  assign t0_r5_c10_rr13 = a_5_13 * b_13_10;
  assign t0_r5_c10_rr14 = a_5_14 * b_14_10;
  assign t1_r5_c10_rr0 = t0_r5_c10_rr0 + t0_r5_c10_rr1;
  assign t1_r5_c10_rr1 = t0_r5_c10_rr2 + t0_r5_c10_rr3;
  assign t1_r5_c10_rr2 = t0_r5_c10_rr4 + t0_r5_c10_rr5;
  assign t1_r5_c10_rr3 = t0_r5_c10_rr6 + t0_r5_c10_rr7;
  assign t1_r5_c10_rr4 = t0_r5_c10_rr8 + t0_r5_c10_rr9;
  assign t1_r5_c10_rr5 = t0_r5_c10_rr10 + t0_r5_c10_rr11;
  assign t1_r5_c10_rr6 = t0_r5_c10_rr12 + t0_r5_c10_rr13;
  assign t1_r5_c10_rr7 = t0_r5_c10_rr14;

  assign t2_r5_c10_rr0 = t1_r5_c10_rr0 + t1_r5_c10_rr1;
  assign t2_r5_c10_rr1 = t1_r5_c10_rr2 + t1_r5_c10_rr3;
  assign t2_r5_c10_rr2 = t1_r5_c10_rr4 + t1_r5_c10_rr5;
  assign t2_r5_c10_rr3 = t1_r5_c10_rr6 + t1_r5_c10_rr7;

  assign t3_r5_c10_rr0 = t2_r5_c10_rr0 + t2_r5_c10_rr1;
  assign t3_r5_c10_rr1 = t2_r5_c10_rr2 + t2_r5_c10_rr3;

  assign t4_r5_c10_rr0 = t3_r5_c10_rr0 + t3_r5_c10_rr1;

  assign c_5_10 = t4_r5_c10_rr0;
  assign t0_r5_c11_rr0 = a_5_0 * b_0_11;
  assign t0_r5_c11_rr1 = a_5_1 * b_1_11;
  assign t0_r5_c11_rr2 = a_5_2 * b_2_11;
  assign t0_r5_c11_rr3 = a_5_3 * b_3_11;
  assign t0_r5_c11_rr4 = a_5_4 * b_4_11;
  assign t0_r5_c11_rr5 = a_5_5 * b_5_11;
  assign t0_r5_c11_rr6 = a_5_6 * b_6_11;
  assign t0_r5_c11_rr7 = a_5_7 * b_7_11;
  assign t0_r5_c11_rr8 = a_5_8 * b_8_11;
  assign t0_r5_c11_rr9 = a_5_9 * b_9_11;
  assign t0_r5_c11_rr10 = a_5_10 * b_10_11;
  assign t0_r5_c11_rr11 = a_5_11 * b_11_11;
  assign t0_r5_c11_rr12 = a_5_12 * b_12_11;
  assign t0_r5_c11_rr13 = a_5_13 * b_13_11;
  assign t0_r5_c11_rr14 = a_5_14 * b_14_11;
  assign t1_r5_c11_rr0 = t0_r5_c11_rr0 + t0_r5_c11_rr1;
  assign t1_r5_c11_rr1 = t0_r5_c11_rr2 + t0_r5_c11_rr3;
  assign t1_r5_c11_rr2 = t0_r5_c11_rr4 + t0_r5_c11_rr5;
  assign t1_r5_c11_rr3 = t0_r5_c11_rr6 + t0_r5_c11_rr7;
  assign t1_r5_c11_rr4 = t0_r5_c11_rr8 + t0_r5_c11_rr9;
  assign t1_r5_c11_rr5 = t0_r5_c11_rr10 + t0_r5_c11_rr11;
  assign t1_r5_c11_rr6 = t0_r5_c11_rr12 + t0_r5_c11_rr13;
  assign t1_r5_c11_rr7 = t0_r5_c11_rr14;

  assign t2_r5_c11_rr0 = t1_r5_c11_rr0 + t1_r5_c11_rr1;
  assign t2_r5_c11_rr1 = t1_r5_c11_rr2 + t1_r5_c11_rr3;
  assign t2_r5_c11_rr2 = t1_r5_c11_rr4 + t1_r5_c11_rr5;
  assign t2_r5_c11_rr3 = t1_r5_c11_rr6 + t1_r5_c11_rr7;

  assign t3_r5_c11_rr0 = t2_r5_c11_rr0 + t2_r5_c11_rr1;
  assign t3_r5_c11_rr1 = t2_r5_c11_rr2 + t2_r5_c11_rr3;

  assign t4_r5_c11_rr0 = t3_r5_c11_rr0 + t3_r5_c11_rr1;

  assign c_5_11 = t4_r5_c11_rr0;
  assign t0_r5_c12_rr0 = a_5_0 * b_0_12;
  assign t0_r5_c12_rr1 = a_5_1 * b_1_12;
  assign t0_r5_c12_rr2 = a_5_2 * b_2_12;
  assign t0_r5_c12_rr3 = a_5_3 * b_3_12;
  assign t0_r5_c12_rr4 = a_5_4 * b_4_12;
  assign t0_r5_c12_rr5 = a_5_5 * b_5_12;
  assign t0_r5_c12_rr6 = a_5_6 * b_6_12;
  assign t0_r5_c12_rr7 = a_5_7 * b_7_12;
  assign t0_r5_c12_rr8 = a_5_8 * b_8_12;
  assign t0_r5_c12_rr9 = a_5_9 * b_9_12;
  assign t0_r5_c12_rr10 = a_5_10 * b_10_12;
  assign t0_r5_c12_rr11 = a_5_11 * b_11_12;
  assign t0_r5_c12_rr12 = a_5_12 * b_12_12;
  assign t0_r5_c12_rr13 = a_5_13 * b_13_12;
  assign t0_r5_c12_rr14 = a_5_14 * b_14_12;
  assign t1_r5_c12_rr0 = t0_r5_c12_rr0 + t0_r5_c12_rr1;
  assign t1_r5_c12_rr1 = t0_r5_c12_rr2 + t0_r5_c12_rr3;
  assign t1_r5_c12_rr2 = t0_r5_c12_rr4 + t0_r5_c12_rr5;
  assign t1_r5_c12_rr3 = t0_r5_c12_rr6 + t0_r5_c12_rr7;
  assign t1_r5_c12_rr4 = t0_r5_c12_rr8 + t0_r5_c12_rr9;
  assign t1_r5_c12_rr5 = t0_r5_c12_rr10 + t0_r5_c12_rr11;
  assign t1_r5_c12_rr6 = t0_r5_c12_rr12 + t0_r5_c12_rr13;
  assign t1_r5_c12_rr7 = t0_r5_c12_rr14;

  assign t2_r5_c12_rr0 = t1_r5_c12_rr0 + t1_r5_c12_rr1;
  assign t2_r5_c12_rr1 = t1_r5_c12_rr2 + t1_r5_c12_rr3;
  assign t2_r5_c12_rr2 = t1_r5_c12_rr4 + t1_r5_c12_rr5;
  assign t2_r5_c12_rr3 = t1_r5_c12_rr6 + t1_r5_c12_rr7;

  assign t3_r5_c12_rr0 = t2_r5_c12_rr0 + t2_r5_c12_rr1;
  assign t3_r5_c12_rr1 = t2_r5_c12_rr2 + t2_r5_c12_rr3;

  assign t4_r5_c12_rr0 = t3_r5_c12_rr0 + t3_r5_c12_rr1;

  assign c_5_12 = t4_r5_c12_rr0;
  assign t0_r5_c13_rr0 = a_5_0 * b_0_13;
  assign t0_r5_c13_rr1 = a_5_1 * b_1_13;
  assign t0_r5_c13_rr2 = a_5_2 * b_2_13;
  assign t0_r5_c13_rr3 = a_5_3 * b_3_13;
  assign t0_r5_c13_rr4 = a_5_4 * b_4_13;
  assign t0_r5_c13_rr5 = a_5_5 * b_5_13;
  assign t0_r5_c13_rr6 = a_5_6 * b_6_13;
  assign t0_r5_c13_rr7 = a_5_7 * b_7_13;
  assign t0_r5_c13_rr8 = a_5_8 * b_8_13;
  assign t0_r5_c13_rr9 = a_5_9 * b_9_13;
  assign t0_r5_c13_rr10 = a_5_10 * b_10_13;
  assign t0_r5_c13_rr11 = a_5_11 * b_11_13;
  assign t0_r5_c13_rr12 = a_5_12 * b_12_13;
  assign t0_r5_c13_rr13 = a_5_13 * b_13_13;
  assign t0_r5_c13_rr14 = a_5_14 * b_14_13;
  assign t1_r5_c13_rr0 = t0_r5_c13_rr0 + t0_r5_c13_rr1;
  assign t1_r5_c13_rr1 = t0_r5_c13_rr2 + t0_r5_c13_rr3;
  assign t1_r5_c13_rr2 = t0_r5_c13_rr4 + t0_r5_c13_rr5;
  assign t1_r5_c13_rr3 = t0_r5_c13_rr6 + t0_r5_c13_rr7;
  assign t1_r5_c13_rr4 = t0_r5_c13_rr8 + t0_r5_c13_rr9;
  assign t1_r5_c13_rr5 = t0_r5_c13_rr10 + t0_r5_c13_rr11;
  assign t1_r5_c13_rr6 = t0_r5_c13_rr12 + t0_r5_c13_rr13;
  assign t1_r5_c13_rr7 = t0_r5_c13_rr14;

  assign t2_r5_c13_rr0 = t1_r5_c13_rr0 + t1_r5_c13_rr1;
  assign t2_r5_c13_rr1 = t1_r5_c13_rr2 + t1_r5_c13_rr3;
  assign t2_r5_c13_rr2 = t1_r5_c13_rr4 + t1_r5_c13_rr5;
  assign t2_r5_c13_rr3 = t1_r5_c13_rr6 + t1_r5_c13_rr7;

  assign t3_r5_c13_rr0 = t2_r5_c13_rr0 + t2_r5_c13_rr1;
  assign t3_r5_c13_rr1 = t2_r5_c13_rr2 + t2_r5_c13_rr3;

  assign t4_r5_c13_rr0 = t3_r5_c13_rr0 + t3_r5_c13_rr1;

  assign c_5_13 = t4_r5_c13_rr0;
  assign t0_r5_c14_rr0 = a_5_0 * b_0_14;
  assign t0_r5_c14_rr1 = a_5_1 * b_1_14;
  assign t0_r5_c14_rr2 = a_5_2 * b_2_14;
  assign t0_r5_c14_rr3 = a_5_3 * b_3_14;
  assign t0_r5_c14_rr4 = a_5_4 * b_4_14;
  assign t0_r5_c14_rr5 = a_5_5 * b_5_14;
  assign t0_r5_c14_rr6 = a_5_6 * b_6_14;
  assign t0_r5_c14_rr7 = a_5_7 * b_7_14;
  assign t0_r5_c14_rr8 = a_5_8 * b_8_14;
  assign t0_r5_c14_rr9 = a_5_9 * b_9_14;
  assign t0_r5_c14_rr10 = a_5_10 * b_10_14;
  assign t0_r5_c14_rr11 = a_5_11 * b_11_14;
  assign t0_r5_c14_rr12 = a_5_12 * b_12_14;
  assign t0_r5_c14_rr13 = a_5_13 * b_13_14;
  assign t0_r5_c14_rr14 = a_5_14 * b_14_14;
  assign t1_r5_c14_rr0 = t0_r5_c14_rr0 + t0_r5_c14_rr1;
  assign t1_r5_c14_rr1 = t0_r5_c14_rr2 + t0_r5_c14_rr3;
  assign t1_r5_c14_rr2 = t0_r5_c14_rr4 + t0_r5_c14_rr5;
  assign t1_r5_c14_rr3 = t0_r5_c14_rr6 + t0_r5_c14_rr7;
  assign t1_r5_c14_rr4 = t0_r5_c14_rr8 + t0_r5_c14_rr9;
  assign t1_r5_c14_rr5 = t0_r5_c14_rr10 + t0_r5_c14_rr11;
  assign t1_r5_c14_rr6 = t0_r5_c14_rr12 + t0_r5_c14_rr13;
  assign t1_r5_c14_rr7 = t0_r5_c14_rr14;

  assign t2_r5_c14_rr0 = t1_r5_c14_rr0 + t1_r5_c14_rr1;
  assign t2_r5_c14_rr1 = t1_r5_c14_rr2 + t1_r5_c14_rr3;
  assign t2_r5_c14_rr2 = t1_r5_c14_rr4 + t1_r5_c14_rr5;
  assign t2_r5_c14_rr3 = t1_r5_c14_rr6 + t1_r5_c14_rr7;

  assign t3_r5_c14_rr0 = t2_r5_c14_rr0 + t2_r5_c14_rr1;
  assign t3_r5_c14_rr1 = t2_r5_c14_rr2 + t2_r5_c14_rr3;

  assign t4_r5_c14_rr0 = t3_r5_c14_rr0 + t3_r5_c14_rr1;

  assign c_5_14 = t4_r5_c14_rr0;
  assign t0_r6_c0_rr0 = a_6_0 * b_0_0;
  assign t0_r6_c0_rr1 = a_6_1 * b_1_0;
  assign t0_r6_c0_rr2 = a_6_2 * b_2_0;
  assign t0_r6_c0_rr3 = a_6_3 * b_3_0;
  assign t0_r6_c0_rr4 = a_6_4 * b_4_0;
  assign t0_r6_c0_rr5 = a_6_5 * b_5_0;
  assign t0_r6_c0_rr6 = a_6_6 * b_6_0;
  assign t0_r6_c0_rr7 = a_6_7 * b_7_0;
  assign t0_r6_c0_rr8 = a_6_8 * b_8_0;
  assign t0_r6_c0_rr9 = a_6_9 * b_9_0;
  assign t0_r6_c0_rr10 = a_6_10 * b_10_0;
  assign t0_r6_c0_rr11 = a_6_11 * b_11_0;
  assign t0_r6_c0_rr12 = a_6_12 * b_12_0;
  assign t0_r6_c0_rr13 = a_6_13 * b_13_0;
  assign t0_r6_c0_rr14 = a_6_14 * b_14_0;
  assign t1_r6_c0_rr0 = t0_r6_c0_rr0 + t0_r6_c0_rr1;
  assign t1_r6_c0_rr1 = t0_r6_c0_rr2 + t0_r6_c0_rr3;
  assign t1_r6_c0_rr2 = t0_r6_c0_rr4 + t0_r6_c0_rr5;
  assign t1_r6_c0_rr3 = t0_r6_c0_rr6 + t0_r6_c0_rr7;
  assign t1_r6_c0_rr4 = t0_r6_c0_rr8 + t0_r6_c0_rr9;
  assign t1_r6_c0_rr5 = t0_r6_c0_rr10 + t0_r6_c0_rr11;
  assign t1_r6_c0_rr6 = t0_r6_c0_rr12 + t0_r6_c0_rr13;
  assign t1_r6_c0_rr7 = t0_r6_c0_rr14;

  assign t2_r6_c0_rr0 = t1_r6_c0_rr0 + t1_r6_c0_rr1;
  assign t2_r6_c0_rr1 = t1_r6_c0_rr2 + t1_r6_c0_rr3;
  assign t2_r6_c0_rr2 = t1_r6_c0_rr4 + t1_r6_c0_rr5;
  assign t2_r6_c0_rr3 = t1_r6_c0_rr6 + t1_r6_c0_rr7;

  assign t3_r6_c0_rr0 = t2_r6_c0_rr0 + t2_r6_c0_rr1;
  assign t3_r6_c0_rr1 = t2_r6_c0_rr2 + t2_r6_c0_rr3;

  assign t4_r6_c0_rr0 = t3_r6_c0_rr0 + t3_r6_c0_rr1;

  assign c_6_0 = t4_r6_c0_rr0;
  assign t0_r6_c1_rr0 = a_6_0 * b_0_1;
  assign t0_r6_c1_rr1 = a_6_1 * b_1_1;
  assign t0_r6_c1_rr2 = a_6_2 * b_2_1;
  assign t0_r6_c1_rr3 = a_6_3 * b_3_1;
  assign t0_r6_c1_rr4 = a_6_4 * b_4_1;
  assign t0_r6_c1_rr5 = a_6_5 * b_5_1;
  assign t0_r6_c1_rr6 = a_6_6 * b_6_1;
  assign t0_r6_c1_rr7 = a_6_7 * b_7_1;
  assign t0_r6_c1_rr8 = a_6_8 * b_8_1;
  assign t0_r6_c1_rr9 = a_6_9 * b_9_1;
  assign t0_r6_c1_rr10 = a_6_10 * b_10_1;
  assign t0_r6_c1_rr11 = a_6_11 * b_11_1;
  assign t0_r6_c1_rr12 = a_6_12 * b_12_1;
  assign t0_r6_c1_rr13 = a_6_13 * b_13_1;
  assign t0_r6_c1_rr14 = a_6_14 * b_14_1;
  assign t1_r6_c1_rr0 = t0_r6_c1_rr0 + t0_r6_c1_rr1;
  assign t1_r6_c1_rr1 = t0_r6_c1_rr2 + t0_r6_c1_rr3;
  assign t1_r6_c1_rr2 = t0_r6_c1_rr4 + t0_r6_c1_rr5;
  assign t1_r6_c1_rr3 = t0_r6_c1_rr6 + t0_r6_c1_rr7;
  assign t1_r6_c1_rr4 = t0_r6_c1_rr8 + t0_r6_c1_rr9;
  assign t1_r6_c1_rr5 = t0_r6_c1_rr10 + t0_r6_c1_rr11;
  assign t1_r6_c1_rr6 = t0_r6_c1_rr12 + t0_r6_c1_rr13;
  assign t1_r6_c1_rr7 = t0_r6_c1_rr14;

  assign t2_r6_c1_rr0 = t1_r6_c1_rr0 + t1_r6_c1_rr1;
  assign t2_r6_c1_rr1 = t1_r6_c1_rr2 + t1_r6_c1_rr3;
  assign t2_r6_c1_rr2 = t1_r6_c1_rr4 + t1_r6_c1_rr5;
  assign t2_r6_c1_rr3 = t1_r6_c1_rr6 + t1_r6_c1_rr7;

  assign t3_r6_c1_rr0 = t2_r6_c1_rr0 + t2_r6_c1_rr1;
  assign t3_r6_c1_rr1 = t2_r6_c1_rr2 + t2_r6_c1_rr3;

  assign t4_r6_c1_rr0 = t3_r6_c1_rr0 + t3_r6_c1_rr1;

  assign c_6_1 = t4_r6_c1_rr0;
  assign t0_r6_c2_rr0 = a_6_0 * b_0_2;
  assign t0_r6_c2_rr1 = a_6_1 * b_1_2;
  assign t0_r6_c2_rr2 = a_6_2 * b_2_2;
  assign t0_r6_c2_rr3 = a_6_3 * b_3_2;
  assign t0_r6_c2_rr4 = a_6_4 * b_4_2;
  assign t0_r6_c2_rr5 = a_6_5 * b_5_2;
  assign t0_r6_c2_rr6 = a_6_6 * b_6_2;
  assign t0_r6_c2_rr7 = a_6_7 * b_7_2;
  assign t0_r6_c2_rr8 = a_6_8 * b_8_2;
  assign t0_r6_c2_rr9 = a_6_9 * b_9_2;
  assign t0_r6_c2_rr10 = a_6_10 * b_10_2;
  assign t0_r6_c2_rr11 = a_6_11 * b_11_2;
  assign t0_r6_c2_rr12 = a_6_12 * b_12_2;
  assign t0_r6_c2_rr13 = a_6_13 * b_13_2;
  assign t0_r6_c2_rr14 = a_6_14 * b_14_2;
  assign t1_r6_c2_rr0 = t0_r6_c2_rr0 + t0_r6_c2_rr1;
  assign t1_r6_c2_rr1 = t0_r6_c2_rr2 + t0_r6_c2_rr3;
  assign t1_r6_c2_rr2 = t0_r6_c2_rr4 + t0_r6_c2_rr5;
  assign t1_r6_c2_rr3 = t0_r6_c2_rr6 + t0_r6_c2_rr7;
  assign t1_r6_c2_rr4 = t0_r6_c2_rr8 + t0_r6_c2_rr9;
  assign t1_r6_c2_rr5 = t0_r6_c2_rr10 + t0_r6_c2_rr11;
  assign t1_r6_c2_rr6 = t0_r6_c2_rr12 + t0_r6_c2_rr13;
  assign t1_r6_c2_rr7 = t0_r6_c2_rr14;

  assign t2_r6_c2_rr0 = t1_r6_c2_rr0 + t1_r6_c2_rr1;
  assign t2_r6_c2_rr1 = t1_r6_c2_rr2 + t1_r6_c2_rr3;
  assign t2_r6_c2_rr2 = t1_r6_c2_rr4 + t1_r6_c2_rr5;
  assign t2_r6_c2_rr3 = t1_r6_c2_rr6 + t1_r6_c2_rr7;

  assign t3_r6_c2_rr0 = t2_r6_c2_rr0 + t2_r6_c2_rr1;
  assign t3_r6_c2_rr1 = t2_r6_c2_rr2 + t2_r6_c2_rr3;

  assign t4_r6_c2_rr0 = t3_r6_c2_rr0 + t3_r6_c2_rr1;

  assign c_6_2 = t4_r6_c2_rr0;
  assign t0_r6_c3_rr0 = a_6_0 * b_0_3;
  assign t0_r6_c3_rr1 = a_6_1 * b_1_3;
  assign t0_r6_c3_rr2 = a_6_2 * b_2_3;
  assign t0_r6_c3_rr3 = a_6_3 * b_3_3;
  assign t0_r6_c3_rr4 = a_6_4 * b_4_3;
  assign t0_r6_c3_rr5 = a_6_5 * b_5_3;
  assign t0_r6_c3_rr6 = a_6_6 * b_6_3;
  assign t0_r6_c3_rr7 = a_6_7 * b_7_3;
  assign t0_r6_c3_rr8 = a_6_8 * b_8_3;
  assign t0_r6_c3_rr9 = a_6_9 * b_9_3;
  assign t0_r6_c3_rr10 = a_6_10 * b_10_3;
  assign t0_r6_c3_rr11 = a_6_11 * b_11_3;
  assign t0_r6_c3_rr12 = a_6_12 * b_12_3;
  assign t0_r6_c3_rr13 = a_6_13 * b_13_3;
  assign t0_r6_c3_rr14 = a_6_14 * b_14_3;
  assign t1_r6_c3_rr0 = t0_r6_c3_rr0 + t0_r6_c3_rr1;
  assign t1_r6_c3_rr1 = t0_r6_c3_rr2 + t0_r6_c3_rr3;
  assign t1_r6_c3_rr2 = t0_r6_c3_rr4 + t0_r6_c3_rr5;
  assign t1_r6_c3_rr3 = t0_r6_c3_rr6 + t0_r6_c3_rr7;
  assign t1_r6_c3_rr4 = t0_r6_c3_rr8 + t0_r6_c3_rr9;
  assign t1_r6_c3_rr5 = t0_r6_c3_rr10 + t0_r6_c3_rr11;
  assign t1_r6_c3_rr6 = t0_r6_c3_rr12 + t0_r6_c3_rr13;
  assign t1_r6_c3_rr7 = t0_r6_c3_rr14;

  assign t2_r6_c3_rr0 = t1_r6_c3_rr0 + t1_r6_c3_rr1;
  assign t2_r6_c3_rr1 = t1_r6_c3_rr2 + t1_r6_c3_rr3;
  assign t2_r6_c3_rr2 = t1_r6_c3_rr4 + t1_r6_c3_rr5;
  assign t2_r6_c3_rr3 = t1_r6_c3_rr6 + t1_r6_c3_rr7;

  assign t3_r6_c3_rr0 = t2_r6_c3_rr0 + t2_r6_c3_rr1;
  assign t3_r6_c3_rr1 = t2_r6_c3_rr2 + t2_r6_c3_rr3;

  assign t4_r6_c3_rr0 = t3_r6_c3_rr0 + t3_r6_c3_rr1;

  assign c_6_3 = t4_r6_c3_rr0;
  assign t0_r6_c4_rr0 = a_6_0 * b_0_4;
  assign t0_r6_c4_rr1 = a_6_1 * b_1_4;
  assign t0_r6_c4_rr2 = a_6_2 * b_2_4;
  assign t0_r6_c4_rr3 = a_6_3 * b_3_4;
  assign t0_r6_c4_rr4 = a_6_4 * b_4_4;
  assign t0_r6_c4_rr5 = a_6_5 * b_5_4;
  assign t0_r6_c4_rr6 = a_6_6 * b_6_4;
  assign t0_r6_c4_rr7 = a_6_7 * b_7_4;
  assign t0_r6_c4_rr8 = a_6_8 * b_8_4;
  assign t0_r6_c4_rr9 = a_6_9 * b_9_4;
  assign t0_r6_c4_rr10 = a_6_10 * b_10_4;
  assign t0_r6_c4_rr11 = a_6_11 * b_11_4;
  assign t0_r6_c4_rr12 = a_6_12 * b_12_4;
  assign t0_r6_c4_rr13 = a_6_13 * b_13_4;
  assign t0_r6_c4_rr14 = a_6_14 * b_14_4;
  assign t1_r6_c4_rr0 = t0_r6_c4_rr0 + t0_r6_c4_rr1;
  assign t1_r6_c4_rr1 = t0_r6_c4_rr2 + t0_r6_c4_rr3;
  assign t1_r6_c4_rr2 = t0_r6_c4_rr4 + t0_r6_c4_rr5;
  assign t1_r6_c4_rr3 = t0_r6_c4_rr6 + t0_r6_c4_rr7;
  assign t1_r6_c4_rr4 = t0_r6_c4_rr8 + t0_r6_c4_rr9;
  assign t1_r6_c4_rr5 = t0_r6_c4_rr10 + t0_r6_c4_rr11;
  assign t1_r6_c4_rr6 = t0_r6_c4_rr12 + t0_r6_c4_rr13;
  assign t1_r6_c4_rr7 = t0_r6_c4_rr14;

  assign t2_r6_c4_rr0 = t1_r6_c4_rr0 + t1_r6_c4_rr1;
  assign t2_r6_c4_rr1 = t1_r6_c4_rr2 + t1_r6_c4_rr3;
  assign t2_r6_c4_rr2 = t1_r6_c4_rr4 + t1_r6_c4_rr5;
  assign t2_r6_c4_rr3 = t1_r6_c4_rr6 + t1_r6_c4_rr7;

  assign t3_r6_c4_rr0 = t2_r6_c4_rr0 + t2_r6_c4_rr1;
  assign t3_r6_c4_rr1 = t2_r6_c4_rr2 + t2_r6_c4_rr3;

  assign t4_r6_c4_rr0 = t3_r6_c4_rr0 + t3_r6_c4_rr1;

  assign c_6_4 = t4_r6_c4_rr0;
  assign t0_r6_c5_rr0 = a_6_0 * b_0_5;
  assign t0_r6_c5_rr1 = a_6_1 * b_1_5;
  assign t0_r6_c5_rr2 = a_6_2 * b_2_5;
  assign t0_r6_c5_rr3 = a_6_3 * b_3_5;
  assign t0_r6_c5_rr4 = a_6_4 * b_4_5;
  assign t0_r6_c5_rr5 = a_6_5 * b_5_5;
  assign t0_r6_c5_rr6 = a_6_6 * b_6_5;
  assign t0_r6_c5_rr7 = a_6_7 * b_7_5;
  assign t0_r6_c5_rr8 = a_6_8 * b_8_5;
  assign t0_r6_c5_rr9 = a_6_9 * b_9_5;
  assign t0_r6_c5_rr10 = a_6_10 * b_10_5;
  assign t0_r6_c5_rr11 = a_6_11 * b_11_5;
  assign t0_r6_c5_rr12 = a_6_12 * b_12_5;
  assign t0_r6_c5_rr13 = a_6_13 * b_13_5;
  assign t0_r6_c5_rr14 = a_6_14 * b_14_5;
  assign t1_r6_c5_rr0 = t0_r6_c5_rr0 + t0_r6_c5_rr1;
  assign t1_r6_c5_rr1 = t0_r6_c5_rr2 + t0_r6_c5_rr3;
  assign t1_r6_c5_rr2 = t0_r6_c5_rr4 + t0_r6_c5_rr5;
  assign t1_r6_c5_rr3 = t0_r6_c5_rr6 + t0_r6_c5_rr7;
  assign t1_r6_c5_rr4 = t0_r6_c5_rr8 + t0_r6_c5_rr9;
  assign t1_r6_c5_rr5 = t0_r6_c5_rr10 + t0_r6_c5_rr11;
  assign t1_r6_c5_rr6 = t0_r6_c5_rr12 + t0_r6_c5_rr13;
  assign t1_r6_c5_rr7 = t0_r6_c5_rr14;

  assign t2_r6_c5_rr0 = t1_r6_c5_rr0 + t1_r6_c5_rr1;
  assign t2_r6_c5_rr1 = t1_r6_c5_rr2 + t1_r6_c5_rr3;
  assign t2_r6_c5_rr2 = t1_r6_c5_rr4 + t1_r6_c5_rr5;
  assign t2_r6_c5_rr3 = t1_r6_c5_rr6 + t1_r6_c5_rr7;

  assign t3_r6_c5_rr0 = t2_r6_c5_rr0 + t2_r6_c5_rr1;
  assign t3_r6_c5_rr1 = t2_r6_c5_rr2 + t2_r6_c5_rr3;

  assign t4_r6_c5_rr0 = t3_r6_c5_rr0 + t3_r6_c5_rr1;

  assign c_6_5 = t4_r6_c5_rr0;
  assign t0_r6_c6_rr0 = a_6_0 * b_0_6;
  assign t0_r6_c6_rr1 = a_6_1 * b_1_6;
  assign t0_r6_c6_rr2 = a_6_2 * b_2_6;
  assign t0_r6_c6_rr3 = a_6_3 * b_3_6;
  assign t0_r6_c6_rr4 = a_6_4 * b_4_6;
  assign t0_r6_c6_rr5 = a_6_5 * b_5_6;
  assign t0_r6_c6_rr6 = a_6_6 * b_6_6;
  assign t0_r6_c6_rr7 = a_6_7 * b_7_6;
  assign t0_r6_c6_rr8 = a_6_8 * b_8_6;
  assign t0_r6_c6_rr9 = a_6_9 * b_9_6;
  assign t0_r6_c6_rr10 = a_6_10 * b_10_6;
  assign t0_r6_c6_rr11 = a_6_11 * b_11_6;
  assign t0_r6_c6_rr12 = a_6_12 * b_12_6;
  assign t0_r6_c6_rr13 = a_6_13 * b_13_6;
  assign t0_r6_c6_rr14 = a_6_14 * b_14_6;
  assign t1_r6_c6_rr0 = t0_r6_c6_rr0 + t0_r6_c6_rr1;
  assign t1_r6_c6_rr1 = t0_r6_c6_rr2 + t0_r6_c6_rr3;
  assign t1_r6_c6_rr2 = t0_r6_c6_rr4 + t0_r6_c6_rr5;
  assign t1_r6_c6_rr3 = t0_r6_c6_rr6 + t0_r6_c6_rr7;
  assign t1_r6_c6_rr4 = t0_r6_c6_rr8 + t0_r6_c6_rr9;
  assign t1_r6_c6_rr5 = t0_r6_c6_rr10 + t0_r6_c6_rr11;
  assign t1_r6_c6_rr6 = t0_r6_c6_rr12 + t0_r6_c6_rr13;
  assign t1_r6_c6_rr7 = t0_r6_c6_rr14;

  assign t2_r6_c6_rr0 = t1_r6_c6_rr0 + t1_r6_c6_rr1;
  assign t2_r6_c6_rr1 = t1_r6_c6_rr2 + t1_r6_c6_rr3;
  assign t2_r6_c6_rr2 = t1_r6_c6_rr4 + t1_r6_c6_rr5;
  assign t2_r6_c6_rr3 = t1_r6_c6_rr6 + t1_r6_c6_rr7;

  assign t3_r6_c6_rr0 = t2_r6_c6_rr0 + t2_r6_c6_rr1;
  assign t3_r6_c6_rr1 = t2_r6_c6_rr2 + t2_r6_c6_rr3;

  assign t4_r6_c6_rr0 = t3_r6_c6_rr0 + t3_r6_c6_rr1;

  assign c_6_6 = t4_r6_c6_rr0;
  assign t0_r6_c7_rr0 = a_6_0 * b_0_7;
  assign t0_r6_c7_rr1 = a_6_1 * b_1_7;
  assign t0_r6_c7_rr2 = a_6_2 * b_2_7;
  assign t0_r6_c7_rr3 = a_6_3 * b_3_7;
  assign t0_r6_c7_rr4 = a_6_4 * b_4_7;
  assign t0_r6_c7_rr5 = a_6_5 * b_5_7;
  assign t0_r6_c7_rr6 = a_6_6 * b_6_7;
  assign t0_r6_c7_rr7 = a_6_7 * b_7_7;
  assign t0_r6_c7_rr8 = a_6_8 * b_8_7;
  assign t0_r6_c7_rr9 = a_6_9 * b_9_7;
  assign t0_r6_c7_rr10 = a_6_10 * b_10_7;
  assign t0_r6_c7_rr11 = a_6_11 * b_11_7;
  assign t0_r6_c7_rr12 = a_6_12 * b_12_7;
  assign t0_r6_c7_rr13 = a_6_13 * b_13_7;
  assign t0_r6_c7_rr14 = a_6_14 * b_14_7;
  assign t1_r6_c7_rr0 = t0_r6_c7_rr0 + t0_r6_c7_rr1;
  assign t1_r6_c7_rr1 = t0_r6_c7_rr2 + t0_r6_c7_rr3;
  assign t1_r6_c7_rr2 = t0_r6_c7_rr4 + t0_r6_c7_rr5;
  assign t1_r6_c7_rr3 = t0_r6_c7_rr6 + t0_r6_c7_rr7;
  assign t1_r6_c7_rr4 = t0_r6_c7_rr8 + t0_r6_c7_rr9;
  assign t1_r6_c7_rr5 = t0_r6_c7_rr10 + t0_r6_c7_rr11;
  assign t1_r6_c7_rr6 = t0_r6_c7_rr12 + t0_r6_c7_rr13;
  assign t1_r6_c7_rr7 = t0_r6_c7_rr14;

  assign t2_r6_c7_rr0 = t1_r6_c7_rr0 + t1_r6_c7_rr1;
  assign t2_r6_c7_rr1 = t1_r6_c7_rr2 + t1_r6_c7_rr3;
  assign t2_r6_c7_rr2 = t1_r6_c7_rr4 + t1_r6_c7_rr5;
  assign t2_r6_c7_rr3 = t1_r6_c7_rr6 + t1_r6_c7_rr7;

  assign t3_r6_c7_rr0 = t2_r6_c7_rr0 + t2_r6_c7_rr1;
  assign t3_r6_c7_rr1 = t2_r6_c7_rr2 + t2_r6_c7_rr3;

  assign t4_r6_c7_rr0 = t3_r6_c7_rr0 + t3_r6_c7_rr1;

  assign c_6_7 = t4_r6_c7_rr0;
  assign t0_r6_c8_rr0 = a_6_0 * b_0_8;
  assign t0_r6_c8_rr1 = a_6_1 * b_1_8;
  assign t0_r6_c8_rr2 = a_6_2 * b_2_8;
  assign t0_r6_c8_rr3 = a_6_3 * b_3_8;
  assign t0_r6_c8_rr4 = a_6_4 * b_4_8;
  assign t0_r6_c8_rr5 = a_6_5 * b_5_8;
  assign t0_r6_c8_rr6 = a_6_6 * b_6_8;
  assign t0_r6_c8_rr7 = a_6_7 * b_7_8;
  assign t0_r6_c8_rr8 = a_6_8 * b_8_8;
  assign t0_r6_c8_rr9 = a_6_9 * b_9_8;
  assign t0_r6_c8_rr10 = a_6_10 * b_10_8;
  assign t0_r6_c8_rr11 = a_6_11 * b_11_8;
  assign t0_r6_c8_rr12 = a_6_12 * b_12_8;
  assign t0_r6_c8_rr13 = a_6_13 * b_13_8;
  assign t0_r6_c8_rr14 = a_6_14 * b_14_8;
  assign t1_r6_c8_rr0 = t0_r6_c8_rr0 + t0_r6_c8_rr1;
  assign t1_r6_c8_rr1 = t0_r6_c8_rr2 + t0_r6_c8_rr3;
  assign t1_r6_c8_rr2 = t0_r6_c8_rr4 + t0_r6_c8_rr5;
  assign t1_r6_c8_rr3 = t0_r6_c8_rr6 + t0_r6_c8_rr7;
  assign t1_r6_c8_rr4 = t0_r6_c8_rr8 + t0_r6_c8_rr9;
  assign t1_r6_c8_rr5 = t0_r6_c8_rr10 + t0_r6_c8_rr11;
  assign t1_r6_c8_rr6 = t0_r6_c8_rr12 + t0_r6_c8_rr13;
  assign t1_r6_c8_rr7 = t0_r6_c8_rr14;

  assign t2_r6_c8_rr0 = t1_r6_c8_rr0 + t1_r6_c8_rr1;
  assign t2_r6_c8_rr1 = t1_r6_c8_rr2 + t1_r6_c8_rr3;
  assign t2_r6_c8_rr2 = t1_r6_c8_rr4 + t1_r6_c8_rr5;
  assign t2_r6_c8_rr3 = t1_r6_c8_rr6 + t1_r6_c8_rr7;

  assign t3_r6_c8_rr0 = t2_r6_c8_rr0 + t2_r6_c8_rr1;
  assign t3_r6_c8_rr1 = t2_r6_c8_rr2 + t2_r6_c8_rr3;

  assign t4_r6_c8_rr0 = t3_r6_c8_rr0 + t3_r6_c8_rr1;

  assign c_6_8 = t4_r6_c8_rr0;
  assign t0_r6_c9_rr0 = a_6_0 * b_0_9;
  assign t0_r6_c9_rr1 = a_6_1 * b_1_9;
  assign t0_r6_c9_rr2 = a_6_2 * b_2_9;
  assign t0_r6_c9_rr3 = a_6_3 * b_3_9;
  assign t0_r6_c9_rr4 = a_6_4 * b_4_9;
  assign t0_r6_c9_rr5 = a_6_5 * b_5_9;
  assign t0_r6_c9_rr6 = a_6_6 * b_6_9;
  assign t0_r6_c9_rr7 = a_6_7 * b_7_9;
  assign t0_r6_c9_rr8 = a_6_8 * b_8_9;
  assign t0_r6_c9_rr9 = a_6_9 * b_9_9;
  assign t0_r6_c9_rr10 = a_6_10 * b_10_9;
  assign t0_r6_c9_rr11 = a_6_11 * b_11_9;
  assign t0_r6_c9_rr12 = a_6_12 * b_12_9;
  assign t0_r6_c9_rr13 = a_6_13 * b_13_9;
  assign t0_r6_c9_rr14 = a_6_14 * b_14_9;
  assign t1_r6_c9_rr0 = t0_r6_c9_rr0 + t0_r6_c9_rr1;
  assign t1_r6_c9_rr1 = t0_r6_c9_rr2 + t0_r6_c9_rr3;
  assign t1_r6_c9_rr2 = t0_r6_c9_rr4 + t0_r6_c9_rr5;
  assign t1_r6_c9_rr3 = t0_r6_c9_rr6 + t0_r6_c9_rr7;
  assign t1_r6_c9_rr4 = t0_r6_c9_rr8 + t0_r6_c9_rr9;
  assign t1_r6_c9_rr5 = t0_r6_c9_rr10 + t0_r6_c9_rr11;
  assign t1_r6_c9_rr6 = t0_r6_c9_rr12 + t0_r6_c9_rr13;
  assign t1_r6_c9_rr7 = t0_r6_c9_rr14;

  assign t2_r6_c9_rr0 = t1_r6_c9_rr0 + t1_r6_c9_rr1;
  assign t2_r6_c9_rr1 = t1_r6_c9_rr2 + t1_r6_c9_rr3;
  assign t2_r6_c9_rr2 = t1_r6_c9_rr4 + t1_r6_c9_rr5;
  assign t2_r6_c9_rr3 = t1_r6_c9_rr6 + t1_r6_c9_rr7;

  assign t3_r6_c9_rr0 = t2_r6_c9_rr0 + t2_r6_c9_rr1;
  assign t3_r6_c9_rr1 = t2_r6_c9_rr2 + t2_r6_c9_rr3;

  assign t4_r6_c9_rr0 = t3_r6_c9_rr0 + t3_r6_c9_rr1;

  assign c_6_9 = t4_r6_c9_rr0;
  assign t0_r6_c10_rr0 = a_6_0 * b_0_10;
  assign t0_r6_c10_rr1 = a_6_1 * b_1_10;
  assign t0_r6_c10_rr2 = a_6_2 * b_2_10;
  assign t0_r6_c10_rr3 = a_6_3 * b_3_10;
  assign t0_r6_c10_rr4 = a_6_4 * b_4_10;
  assign t0_r6_c10_rr5 = a_6_5 * b_5_10;
  assign t0_r6_c10_rr6 = a_6_6 * b_6_10;
  assign t0_r6_c10_rr7 = a_6_7 * b_7_10;
  assign t0_r6_c10_rr8 = a_6_8 * b_8_10;
  assign t0_r6_c10_rr9 = a_6_9 * b_9_10;
  assign t0_r6_c10_rr10 = a_6_10 * b_10_10;
  assign t0_r6_c10_rr11 = a_6_11 * b_11_10;
  assign t0_r6_c10_rr12 = a_6_12 * b_12_10;
  assign t0_r6_c10_rr13 = a_6_13 * b_13_10;
  assign t0_r6_c10_rr14 = a_6_14 * b_14_10;
  assign t1_r6_c10_rr0 = t0_r6_c10_rr0 + t0_r6_c10_rr1;
  assign t1_r6_c10_rr1 = t0_r6_c10_rr2 + t0_r6_c10_rr3;
  assign t1_r6_c10_rr2 = t0_r6_c10_rr4 + t0_r6_c10_rr5;
  assign t1_r6_c10_rr3 = t0_r6_c10_rr6 + t0_r6_c10_rr7;
  assign t1_r6_c10_rr4 = t0_r6_c10_rr8 + t0_r6_c10_rr9;
  assign t1_r6_c10_rr5 = t0_r6_c10_rr10 + t0_r6_c10_rr11;
  assign t1_r6_c10_rr6 = t0_r6_c10_rr12 + t0_r6_c10_rr13;
  assign t1_r6_c10_rr7 = t0_r6_c10_rr14;

  assign t2_r6_c10_rr0 = t1_r6_c10_rr0 + t1_r6_c10_rr1;
  assign t2_r6_c10_rr1 = t1_r6_c10_rr2 + t1_r6_c10_rr3;
  assign t2_r6_c10_rr2 = t1_r6_c10_rr4 + t1_r6_c10_rr5;
  assign t2_r6_c10_rr3 = t1_r6_c10_rr6 + t1_r6_c10_rr7;

  assign t3_r6_c10_rr0 = t2_r6_c10_rr0 + t2_r6_c10_rr1;
  assign t3_r6_c10_rr1 = t2_r6_c10_rr2 + t2_r6_c10_rr3;

  assign t4_r6_c10_rr0 = t3_r6_c10_rr0 + t3_r6_c10_rr1;

  assign c_6_10 = t4_r6_c10_rr0;
  assign t0_r6_c11_rr0 = a_6_0 * b_0_11;
  assign t0_r6_c11_rr1 = a_6_1 * b_1_11;
  assign t0_r6_c11_rr2 = a_6_2 * b_2_11;
  assign t0_r6_c11_rr3 = a_6_3 * b_3_11;
  assign t0_r6_c11_rr4 = a_6_4 * b_4_11;
  assign t0_r6_c11_rr5 = a_6_5 * b_5_11;
  assign t0_r6_c11_rr6 = a_6_6 * b_6_11;
  assign t0_r6_c11_rr7 = a_6_7 * b_7_11;
  assign t0_r6_c11_rr8 = a_6_8 * b_8_11;
  assign t0_r6_c11_rr9 = a_6_9 * b_9_11;
  assign t0_r6_c11_rr10 = a_6_10 * b_10_11;
  assign t0_r6_c11_rr11 = a_6_11 * b_11_11;
  assign t0_r6_c11_rr12 = a_6_12 * b_12_11;
  assign t0_r6_c11_rr13 = a_6_13 * b_13_11;
  assign t0_r6_c11_rr14 = a_6_14 * b_14_11;
  assign t1_r6_c11_rr0 = t0_r6_c11_rr0 + t0_r6_c11_rr1;
  assign t1_r6_c11_rr1 = t0_r6_c11_rr2 + t0_r6_c11_rr3;
  assign t1_r6_c11_rr2 = t0_r6_c11_rr4 + t0_r6_c11_rr5;
  assign t1_r6_c11_rr3 = t0_r6_c11_rr6 + t0_r6_c11_rr7;
  assign t1_r6_c11_rr4 = t0_r6_c11_rr8 + t0_r6_c11_rr9;
  assign t1_r6_c11_rr5 = t0_r6_c11_rr10 + t0_r6_c11_rr11;
  assign t1_r6_c11_rr6 = t0_r6_c11_rr12 + t0_r6_c11_rr13;
  assign t1_r6_c11_rr7 = t0_r6_c11_rr14;

  assign t2_r6_c11_rr0 = t1_r6_c11_rr0 + t1_r6_c11_rr1;
  assign t2_r6_c11_rr1 = t1_r6_c11_rr2 + t1_r6_c11_rr3;
  assign t2_r6_c11_rr2 = t1_r6_c11_rr4 + t1_r6_c11_rr5;
  assign t2_r6_c11_rr3 = t1_r6_c11_rr6 + t1_r6_c11_rr7;

  assign t3_r6_c11_rr0 = t2_r6_c11_rr0 + t2_r6_c11_rr1;
  assign t3_r6_c11_rr1 = t2_r6_c11_rr2 + t2_r6_c11_rr3;

  assign t4_r6_c11_rr0 = t3_r6_c11_rr0 + t3_r6_c11_rr1;

  assign c_6_11 = t4_r6_c11_rr0;
  assign t0_r6_c12_rr0 = a_6_0 * b_0_12;
  assign t0_r6_c12_rr1 = a_6_1 * b_1_12;
  assign t0_r6_c12_rr2 = a_6_2 * b_2_12;
  assign t0_r6_c12_rr3 = a_6_3 * b_3_12;
  assign t0_r6_c12_rr4 = a_6_4 * b_4_12;
  assign t0_r6_c12_rr5 = a_6_5 * b_5_12;
  assign t0_r6_c12_rr6 = a_6_6 * b_6_12;
  assign t0_r6_c12_rr7 = a_6_7 * b_7_12;
  assign t0_r6_c12_rr8 = a_6_8 * b_8_12;
  assign t0_r6_c12_rr9 = a_6_9 * b_9_12;
  assign t0_r6_c12_rr10 = a_6_10 * b_10_12;
  assign t0_r6_c12_rr11 = a_6_11 * b_11_12;
  assign t0_r6_c12_rr12 = a_6_12 * b_12_12;
  assign t0_r6_c12_rr13 = a_6_13 * b_13_12;
  assign t0_r6_c12_rr14 = a_6_14 * b_14_12;
  assign t1_r6_c12_rr0 = t0_r6_c12_rr0 + t0_r6_c12_rr1;
  assign t1_r6_c12_rr1 = t0_r6_c12_rr2 + t0_r6_c12_rr3;
  assign t1_r6_c12_rr2 = t0_r6_c12_rr4 + t0_r6_c12_rr5;
  assign t1_r6_c12_rr3 = t0_r6_c12_rr6 + t0_r6_c12_rr7;
  assign t1_r6_c12_rr4 = t0_r6_c12_rr8 + t0_r6_c12_rr9;
  assign t1_r6_c12_rr5 = t0_r6_c12_rr10 + t0_r6_c12_rr11;
  assign t1_r6_c12_rr6 = t0_r6_c12_rr12 + t0_r6_c12_rr13;
  assign t1_r6_c12_rr7 = t0_r6_c12_rr14;

  assign t2_r6_c12_rr0 = t1_r6_c12_rr0 + t1_r6_c12_rr1;
  assign t2_r6_c12_rr1 = t1_r6_c12_rr2 + t1_r6_c12_rr3;
  assign t2_r6_c12_rr2 = t1_r6_c12_rr4 + t1_r6_c12_rr5;
  assign t2_r6_c12_rr3 = t1_r6_c12_rr6 + t1_r6_c12_rr7;

  assign t3_r6_c12_rr0 = t2_r6_c12_rr0 + t2_r6_c12_rr1;
  assign t3_r6_c12_rr1 = t2_r6_c12_rr2 + t2_r6_c12_rr3;

  assign t4_r6_c12_rr0 = t3_r6_c12_rr0 + t3_r6_c12_rr1;

  assign c_6_12 = t4_r6_c12_rr0;
  assign t0_r6_c13_rr0 = a_6_0 * b_0_13;
  assign t0_r6_c13_rr1 = a_6_1 * b_1_13;
  assign t0_r6_c13_rr2 = a_6_2 * b_2_13;
  assign t0_r6_c13_rr3 = a_6_3 * b_3_13;
  assign t0_r6_c13_rr4 = a_6_4 * b_4_13;
  assign t0_r6_c13_rr5 = a_6_5 * b_5_13;
  assign t0_r6_c13_rr6 = a_6_6 * b_6_13;
  assign t0_r6_c13_rr7 = a_6_7 * b_7_13;
  assign t0_r6_c13_rr8 = a_6_8 * b_8_13;
  assign t0_r6_c13_rr9 = a_6_9 * b_9_13;
  assign t0_r6_c13_rr10 = a_6_10 * b_10_13;
  assign t0_r6_c13_rr11 = a_6_11 * b_11_13;
  assign t0_r6_c13_rr12 = a_6_12 * b_12_13;
  assign t0_r6_c13_rr13 = a_6_13 * b_13_13;
  assign t0_r6_c13_rr14 = a_6_14 * b_14_13;
  assign t1_r6_c13_rr0 = t0_r6_c13_rr0 + t0_r6_c13_rr1;
  assign t1_r6_c13_rr1 = t0_r6_c13_rr2 + t0_r6_c13_rr3;
  assign t1_r6_c13_rr2 = t0_r6_c13_rr4 + t0_r6_c13_rr5;
  assign t1_r6_c13_rr3 = t0_r6_c13_rr6 + t0_r6_c13_rr7;
  assign t1_r6_c13_rr4 = t0_r6_c13_rr8 + t0_r6_c13_rr9;
  assign t1_r6_c13_rr5 = t0_r6_c13_rr10 + t0_r6_c13_rr11;
  assign t1_r6_c13_rr6 = t0_r6_c13_rr12 + t0_r6_c13_rr13;
  assign t1_r6_c13_rr7 = t0_r6_c13_rr14;

  assign t2_r6_c13_rr0 = t1_r6_c13_rr0 + t1_r6_c13_rr1;
  assign t2_r6_c13_rr1 = t1_r6_c13_rr2 + t1_r6_c13_rr3;
  assign t2_r6_c13_rr2 = t1_r6_c13_rr4 + t1_r6_c13_rr5;
  assign t2_r6_c13_rr3 = t1_r6_c13_rr6 + t1_r6_c13_rr7;

  assign t3_r6_c13_rr0 = t2_r6_c13_rr0 + t2_r6_c13_rr1;
  assign t3_r6_c13_rr1 = t2_r6_c13_rr2 + t2_r6_c13_rr3;

  assign t4_r6_c13_rr0 = t3_r6_c13_rr0 + t3_r6_c13_rr1;

  assign c_6_13 = t4_r6_c13_rr0;
  assign t0_r6_c14_rr0 = a_6_0 * b_0_14;
  assign t0_r6_c14_rr1 = a_6_1 * b_1_14;
  assign t0_r6_c14_rr2 = a_6_2 * b_2_14;
  assign t0_r6_c14_rr3 = a_6_3 * b_3_14;
  assign t0_r6_c14_rr4 = a_6_4 * b_4_14;
  assign t0_r6_c14_rr5 = a_6_5 * b_5_14;
  assign t0_r6_c14_rr6 = a_6_6 * b_6_14;
  assign t0_r6_c14_rr7 = a_6_7 * b_7_14;
  assign t0_r6_c14_rr8 = a_6_8 * b_8_14;
  assign t0_r6_c14_rr9 = a_6_9 * b_9_14;
  assign t0_r6_c14_rr10 = a_6_10 * b_10_14;
  assign t0_r6_c14_rr11 = a_6_11 * b_11_14;
  assign t0_r6_c14_rr12 = a_6_12 * b_12_14;
  assign t0_r6_c14_rr13 = a_6_13 * b_13_14;
  assign t0_r6_c14_rr14 = a_6_14 * b_14_14;
  assign t1_r6_c14_rr0 = t0_r6_c14_rr0 + t0_r6_c14_rr1;
  assign t1_r6_c14_rr1 = t0_r6_c14_rr2 + t0_r6_c14_rr3;
  assign t1_r6_c14_rr2 = t0_r6_c14_rr4 + t0_r6_c14_rr5;
  assign t1_r6_c14_rr3 = t0_r6_c14_rr6 + t0_r6_c14_rr7;
  assign t1_r6_c14_rr4 = t0_r6_c14_rr8 + t0_r6_c14_rr9;
  assign t1_r6_c14_rr5 = t0_r6_c14_rr10 + t0_r6_c14_rr11;
  assign t1_r6_c14_rr6 = t0_r6_c14_rr12 + t0_r6_c14_rr13;
  assign t1_r6_c14_rr7 = t0_r6_c14_rr14;

  assign t2_r6_c14_rr0 = t1_r6_c14_rr0 + t1_r6_c14_rr1;
  assign t2_r6_c14_rr1 = t1_r6_c14_rr2 + t1_r6_c14_rr3;
  assign t2_r6_c14_rr2 = t1_r6_c14_rr4 + t1_r6_c14_rr5;
  assign t2_r6_c14_rr3 = t1_r6_c14_rr6 + t1_r6_c14_rr7;

  assign t3_r6_c14_rr0 = t2_r6_c14_rr0 + t2_r6_c14_rr1;
  assign t3_r6_c14_rr1 = t2_r6_c14_rr2 + t2_r6_c14_rr3;

  assign t4_r6_c14_rr0 = t3_r6_c14_rr0 + t3_r6_c14_rr1;

  assign c_6_14 = t4_r6_c14_rr0;
  assign t0_r7_c0_rr0 = a_7_0 * b_0_0;
  assign t0_r7_c0_rr1 = a_7_1 * b_1_0;
  assign t0_r7_c0_rr2 = a_7_2 * b_2_0;
  assign t0_r7_c0_rr3 = a_7_3 * b_3_0;
  assign t0_r7_c0_rr4 = a_7_4 * b_4_0;
  assign t0_r7_c0_rr5 = a_7_5 * b_5_0;
  assign t0_r7_c0_rr6 = a_7_6 * b_6_0;
  assign t0_r7_c0_rr7 = a_7_7 * b_7_0;
  assign t0_r7_c0_rr8 = a_7_8 * b_8_0;
  assign t0_r7_c0_rr9 = a_7_9 * b_9_0;
  assign t0_r7_c0_rr10 = a_7_10 * b_10_0;
  assign t0_r7_c0_rr11 = a_7_11 * b_11_0;
  assign t0_r7_c0_rr12 = a_7_12 * b_12_0;
  assign t0_r7_c0_rr13 = a_7_13 * b_13_0;
  assign t0_r7_c0_rr14 = a_7_14 * b_14_0;
  assign t1_r7_c0_rr0 = t0_r7_c0_rr0 + t0_r7_c0_rr1;
  assign t1_r7_c0_rr1 = t0_r7_c0_rr2 + t0_r7_c0_rr3;
  assign t1_r7_c0_rr2 = t0_r7_c0_rr4 + t0_r7_c0_rr5;
  assign t1_r7_c0_rr3 = t0_r7_c0_rr6 + t0_r7_c0_rr7;
  assign t1_r7_c0_rr4 = t0_r7_c0_rr8 + t0_r7_c0_rr9;
  assign t1_r7_c0_rr5 = t0_r7_c0_rr10 + t0_r7_c0_rr11;
  assign t1_r7_c0_rr6 = t0_r7_c0_rr12 + t0_r7_c0_rr13;
  assign t1_r7_c0_rr7 = t0_r7_c0_rr14;

  assign t2_r7_c0_rr0 = t1_r7_c0_rr0 + t1_r7_c0_rr1;
  assign t2_r7_c0_rr1 = t1_r7_c0_rr2 + t1_r7_c0_rr3;
  assign t2_r7_c0_rr2 = t1_r7_c0_rr4 + t1_r7_c0_rr5;
  assign t2_r7_c0_rr3 = t1_r7_c0_rr6 + t1_r7_c0_rr7;

  assign t3_r7_c0_rr0 = t2_r7_c0_rr0 + t2_r7_c0_rr1;
  assign t3_r7_c0_rr1 = t2_r7_c0_rr2 + t2_r7_c0_rr3;

  assign t4_r7_c0_rr0 = t3_r7_c0_rr0 + t3_r7_c0_rr1;

  assign c_7_0 = t4_r7_c0_rr0;
  assign t0_r7_c1_rr0 = a_7_0 * b_0_1;
  assign t0_r7_c1_rr1 = a_7_1 * b_1_1;
  assign t0_r7_c1_rr2 = a_7_2 * b_2_1;
  assign t0_r7_c1_rr3 = a_7_3 * b_3_1;
  assign t0_r7_c1_rr4 = a_7_4 * b_4_1;
  assign t0_r7_c1_rr5 = a_7_5 * b_5_1;
  assign t0_r7_c1_rr6 = a_7_6 * b_6_1;
  assign t0_r7_c1_rr7 = a_7_7 * b_7_1;
  assign t0_r7_c1_rr8 = a_7_8 * b_8_1;
  assign t0_r7_c1_rr9 = a_7_9 * b_9_1;
  assign t0_r7_c1_rr10 = a_7_10 * b_10_1;
  assign t0_r7_c1_rr11 = a_7_11 * b_11_1;
  assign t0_r7_c1_rr12 = a_7_12 * b_12_1;
  assign t0_r7_c1_rr13 = a_7_13 * b_13_1;
  assign t0_r7_c1_rr14 = a_7_14 * b_14_1;
  assign t1_r7_c1_rr0 = t0_r7_c1_rr0 + t0_r7_c1_rr1;
  assign t1_r7_c1_rr1 = t0_r7_c1_rr2 + t0_r7_c1_rr3;
  assign t1_r7_c1_rr2 = t0_r7_c1_rr4 + t0_r7_c1_rr5;
  assign t1_r7_c1_rr3 = t0_r7_c1_rr6 + t0_r7_c1_rr7;
  assign t1_r7_c1_rr4 = t0_r7_c1_rr8 + t0_r7_c1_rr9;
  assign t1_r7_c1_rr5 = t0_r7_c1_rr10 + t0_r7_c1_rr11;
  assign t1_r7_c1_rr6 = t0_r7_c1_rr12 + t0_r7_c1_rr13;
  assign t1_r7_c1_rr7 = t0_r7_c1_rr14;

  assign t2_r7_c1_rr0 = t1_r7_c1_rr0 + t1_r7_c1_rr1;
  assign t2_r7_c1_rr1 = t1_r7_c1_rr2 + t1_r7_c1_rr3;
  assign t2_r7_c1_rr2 = t1_r7_c1_rr4 + t1_r7_c1_rr5;
  assign t2_r7_c1_rr3 = t1_r7_c1_rr6 + t1_r7_c1_rr7;

  assign t3_r7_c1_rr0 = t2_r7_c1_rr0 + t2_r7_c1_rr1;
  assign t3_r7_c1_rr1 = t2_r7_c1_rr2 + t2_r7_c1_rr3;

  assign t4_r7_c1_rr0 = t3_r7_c1_rr0 + t3_r7_c1_rr1;

  assign c_7_1 = t4_r7_c1_rr0;
  assign t0_r7_c2_rr0 = a_7_0 * b_0_2;
  assign t0_r7_c2_rr1 = a_7_1 * b_1_2;
  assign t0_r7_c2_rr2 = a_7_2 * b_2_2;
  assign t0_r7_c2_rr3 = a_7_3 * b_3_2;
  assign t0_r7_c2_rr4 = a_7_4 * b_4_2;
  assign t0_r7_c2_rr5 = a_7_5 * b_5_2;
  assign t0_r7_c2_rr6 = a_7_6 * b_6_2;
  assign t0_r7_c2_rr7 = a_7_7 * b_7_2;
  assign t0_r7_c2_rr8 = a_7_8 * b_8_2;
  assign t0_r7_c2_rr9 = a_7_9 * b_9_2;
  assign t0_r7_c2_rr10 = a_7_10 * b_10_2;
  assign t0_r7_c2_rr11 = a_7_11 * b_11_2;
  assign t0_r7_c2_rr12 = a_7_12 * b_12_2;
  assign t0_r7_c2_rr13 = a_7_13 * b_13_2;
  assign t0_r7_c2_rr14 = a_7_14 * b_14_2;
  assign t1_r7_c2_rr0 = t0_r7_c2_rr0 + t0_r7_c2_rr1;
  assign t1_r7_c2_rr1 = t0_r7_c2_rr2 + t0_r7_c2_rr3;
  assign t1_r7_c2_rr2 = t0_r7_c2_rr4 + t0_r7_c2_rr5;
  assign t1_r7_c2_rr3 = t0_r7_c2_rr6 + t0_r7_c2_rr7;
  assign t1_r7_c2_rr4 = t0_r7_c2_rr8 + t0_r7_c2_rr9;
  assign t1_r7_c2_rr5 = t0_r7_c2_rr10 + t0_r7_c2_rr11;
  assign t1_r7_c2_rr6 = t0_r7_c2_rr12 + t0_r7_c2_rr13;
  assign t1_r7_c2_rr7 = t0_r7_c2_rr14;

  assign t2_r7_c2_rr0 = t1_r7_c2_rr0 + t1_r7_c2_rr1;
  assign t2_r7_c2_rr1 = t1_r7_c2_rr2 + t1_r7_c2_rr3;
  assign t2_r7_c2_rr2 = t1_r7_c2_rr4 + t1_r7_c2_rr5;
  assign t2_r7_c2_rr3 = t1_r7_c2_rr6 + t1_r7_c2_rr7;

  assign t3_r7_c2_rr0 = t2_r7_c2_rr0 + t2_r7_c2_rr1;
  assign t3_r7_c2_rr1 = t2_r7_c2_rr2 + t2_r7_c2_rr3;

  assign t4_r7_c2_rr0 = t3_r7_c2_rr0 + t3_r7_c2_rr1;

  assign c_7_2 = t4_r7_c2_rr0;
  assign t0_r7_c3_rr0 = a_7_0 * b_0_3;
  assign t0_r7_c3_rr1 = a_7_1 * b_1_3;
  assign t0_r7_c3_rr2 = a_7_2 * b_2_3;
  assign t0_r7_c3_rr3 = a_7_3 * b_3_3;
  assign t0_r7_c3_rr4 = a_7_4 * b_4_3;
  assign t0_r7_c3_rr5 = a_7_5 * b_5_3;
  assign t0_r7_c3_rr6 = a_7_6 * b_6_3;
  assign t0_r7_c3_rr7 = a_7_7 * b_7_3;
  assign t0_r7_c3_rr8 = a_7_8 * b_8_3;
  assign t0_r7_c3_rr9 = a_7_9 * b_9_3;
  assign t0_r7_c3_rr10 = a_7_10 * b_10_3;
  assign t0_r7_c3_rr11 = a_7_11 * b_11_3;
  assign t0_r7_c3_rr12 = a_7_12 * b_12_3;
  assign t0_r7_c3_rr13 = a_7_13 * b_13_3;
  assign t0_r7_c3_rr14 = a_7_14 * b_14_3;
  assign t1_r7_c3_rr0 = t0_r7_c3_rr0 + t0_r7_c3_rr1;
  assign t1_r7_c3_rr1 = t0_r7_c3_rr2 + t0_r7_c3_rr3;
  assign t1_r7_c3_rr2 = t0_r7_c3_rr4 + t0_r7_c3_rr5;
  assign t1_r7_c3_rr3 = t0_r7_c3_rr6 + t0_r7_c3_rr7;
  assign t1_r7_c3_rr4 = t0_r7_c3_rr8 + t0_r7_c3_rr9;
  assign t1_r7_c3_rr5 = t0_r7_c3_rr10 + t0_r7_c3_rr11;
  assign t1_r7_c3_rr6 = t0_r7_c3_rr12 + t0_r7_c3_rr13;
  assign t1_r7_c3_rr7 = t0_r7_c3_rr14;

  assign t2_r7_c3_rr0 = t1_r7_c3_rr0 + t1_r7_c3_rr1;
  assign t2_r7_c3_rr1 = t1_r7_c3_rr2 + t1_r7_c3_rr3;
  assign t2_r7_c3_rr2 = t1_r7_c3_rr4 + t1_r7_c3_rr5;
  assign t2_r7_c3_rr3 = t1_r7_c3_rr6 + t1_r7_c3_rr7;

  assign t3_r7_c3_rr0 = t2_r7_c3_rr0 + t2_r7_c3_rr1;
  assign t3_r7_c3_rr1 = t2_r7_c3_rr2 + t2_r7_c3_rr3;

  assign t4_r7_c3_rr0 = t3_r7_c3_rr0 + t3_r7_c3_rr1;

  assign c_7_3 = t4_r7_c3_rr0;
  assign t0_r7_c4_rr0 = a_7_0 * b_0_4;
  assign t0_r7_c4_rr1 = a_7_1 * b_1_4;
  assign t0_r7_c4_rr2 = a_7_2 * b_2_4;
  assign t0_r7_c4_rr3 = a_7_3 * b_3_4;
  assign t0_r7_c4_rr4 = a_7_4 * b_4_4;
  assign t0_r7_c4_rr5 = a_7_5 * b_5_4;
  assign t0_r7_c4_rr6 = a_7_6 * b_6_4;
  assign t0_r7_c4_rr7 = a_7_7 * b_7_4;
  assign t0_r7_c4_rr8 = a_7_8 * b_8_4;
  assign t0_r7_c4_rr9 = a_7_9 * b_9_4;
  assign t0_r7_c4_rr10 = a_7_10 * b_10_4;
  assign t0_r7_c4_rr11 = a_7_11 * b_11_4;
  assign t0_r7_c4_rr12 = a_7_12 * b_12_4;
  assign t0_r7_c4_rr13 = a_7_13 * b_13_4;
  assign t0_r7_c4_rr14 = a_7_14 * b_14_4;
  assign t1_r7_c4_rr0 = t0_r7_c4_rr0 + t0_r7_c4_rr1;
  assign t1_r7_c4_rr1 = t0_r7_c4_rr2 + t0_r7_c4_rr3;
  assign t1_r7_c4_rr2 = t0_r7_c4_rr4 + t0_r7_c4_rr5;
  assign t1_r7_c4_rr3 = t0_r7_c4_rr6 + t0_r7_c4_rr7;
  assign t1_r7_c4_rr4 = t0_r7_c4_rr8 + t0_r7_c4_rr9;
  assign t1_r7_c4_rr5 = t0_r7_c4_rr10 + t0_r7_c4_rr11;
  assign t1_r7_c4_rr6 = t0_r7_c4_rr12 + t0_r7_c4_rr13;
  assign t1_r7_c4_rr7 = t0_r7_c4_rr14;

  assign t2_r7_c4_rr0 = t1_r7_c4_rr0 + t1_r7_c4_rr1;
  assign t2_r7_c4_rr1 = t1_r7_c4_rr2 + t1_r7_c4_rr3;
  assign t2_r7_c4_rr2 = t1_r7_c4_rr4 + t1_r7_c4_rr5;
  assign t2_r7_c4_rr3 = t1_r7_c4_rr6 + t1_r7_c4_rr7;

  assign t3_r7_c4_rr0 = t2_r7_c4_rr0 + t2_r7_c4_rr1;
  assign t3_r7_c4_rr1 = t2_r7_c4_rr2 + t2_r7_c4_rr3;

  assign t4_r7_c4_rr0 = t3_r7_c4_rr0 + t3_r7_c4_rr1;

  assign c_7_4 = t4_r7_c4_rr0;
  assign t0_r7_c5_rr0 = a_7_0 * b_0_5;
  assign t0_r7_c5_rr1 = a_7_1 * b_1_5;
  assign t0_r7_c5_rr2 = a_7_2 * b_2_5;
  assign t0_r7_c5_rr3 = a_7_3 * b_3_5;
  assign t0_r7_c5_rr4 = a_7_4 * b_4_5;
  assign t0_r7_c5_rr5 = a_7_5 * b_5_5;
  assign t0_r7_c5_rr6 = a_7_6 * b_6_5;
  assign t0_r7_c5_rr7 = a_7_7 * b_7_5;
  assign t0_r7_c5_rr8 = a_7_8 * b_8_5;
  assign t0_r7_c5_rr9 = a_7_9 * b_9_5;
  assign t0_r7_c5_rr10 = a_7_10 * b_10_5;
  assign t0_r7_c5_rr11 = a_7_11 * b_11_5;
  assign t0_r7_c5_rr12 = a_7_12 * b_12_5;
  assign t0_r7_c5_rr13 = a_7_13 * b_13_5;
  assign t0_r7_c5_rr14 = a_7_14 * b_14_5;
  assign t1_r7_c5_rr0 = t0_r7_c5_rr0 + t0_r7_c5_rr1;
  assign t1_r7_c5_rr1 = t0_r7_c5_rr2 + t0_r7_c5_rr3;
  assign t1_r7_c5_rr2 = t0_r7_c5_rr4 + t0_r7_c5_rr5;
  assign t1_r7_c5_rr3 = t0_r7_c5_rr6 + t0_r7_c5_rr7;
  assign t1_r7_c5_rr4 = t0_r7_c5_rr8 + t0_r7_c5_rr9;
  assign t1_r7_c5_rr5 = t0_r7_c5_rr10 + t0_r7_c5_rr11;
  assign t1_r7_c5_rr6 = t0_r7_c5_rr12 + t0_r7_c5_rr13;
  assign t1_r7_c5_rr7 = t0_r7_c5_rr14;

  assign t2_r7_c5_rr0 = t1_r7_c5_rr0 + t1_r7_c5_rr1;
  assign t2_r7_c5_rr1 = t1_r7_c5_rr2 + t1_r7_c5_rr3;
  assign t2_r7_c5_rr2 = t1_r7_c5_rr4 + t1_r7_c5_rr5;
  assign t2_r7_c5_rr3 = t1_r7_c5_rr6 + t1_r7_c5_rr7;

  assign t3_r7_c5_rr0 = t2_r7_c5_rr0 + t2_r7_c5_rr1;
  assign t3_r7_c5_rr1 = t2_r7_c5_rr2 + t2_r7_c5_rr3;

  assign t4_r7_c5_rr0 = t3_r7_c5_rr0 + t3_r7_c5_rr1;

  assign c_7_5 = t4_r7_c5_rr0;
  assign t0_r7_c6_rr0 = a_7_0 * b_0_6;
  assign t0_r7_c6_rr1 = a_7_1 * b_1_6;
  assign t0_r7_c6_rr2 = a_7_2 * b_2_6;
  assign t0_r7_c6_rr3 = a_7_3 * b_3_6;
  assign t0_r7_c6_rr4 = a_7_4 * b_4_6;
  assign t0_r7_c6_rr5 = a_7_5 * b_5_6;
  assign t0_r7_c6_rr6 = a_7_6 * b_6_6;
  assign t0_r7_c6_rr7 = a_7_7 * b_7_6;
  assign t0_r7_c6_rr8 = a_7_8 * b_8_6;
  assign t0_r7_c6_rr9 = a_7_9 * b_9_6;
  assign t0_r7_c6_rr10 = a_7_10 * b_10_6;
  assign t0_r7_c6_rr11 = a_7_11 * b_11_6;
  assign t0_r7_c6_rr12 = a_7_12 * b_12_6;
  assign t0_r7_c6_rr13 = a_7_13 * b_13_6;
  assign t0_r7_c6_rr14 = a_7_14 * b_14_6;
  assign t1_r7_c6_rr0 = t0_r7_c6_rr0 + t0_r7_c6_rr1;
  assign t1_r7_c6_rr1 = t0_r7_c6_rr2 + t0_r7_c6_rr3;
  assign t1_r7_c6_rr2 = t0_r7_c6_rr4 + t0_r7_c6_rr5;
  assign t1_r7_c6_rr3 = t0_r7_c6_rr6 + t0_r7_c6_rr7;
  assign t1_r7_c6_rr4 = t0_r7_c6_rr8 + t0_r7_c6_rr9;
  assign t1_r7_c6_rr5 = t0_r7_c6_rr10 + t0_r7_c6_rr11;
  assign t1_r7_c6_rr6 = t0_r7_c6_rr12 + t0_r7_c6_rr13;
  assign t1_r7_c6_rr7 = t0_r7_c6_rr14;

  assign t2_r7_c6_rr0 = t1_r7_c6_rr0 + t1_r7_c6_rr1;
  assign t2_r7_c6_rr1 = t1_r7_c6_rr2 + t1_r7_c6_rr3;
  assign t2_r7_c6_rr2 = t1_r7_c6_rr4 + t1_r7_c6_rr5;
  assign t2_r7_c6_rr3 = t1_r7_c6_rr6 + t1_r7_c6_rr7;

  assign t3_r7_c6_rr0 = t2_r7_c6_rr0 + t2_r7_c6_rr1;
  assign t3_r7_c6_rr1 = t2_r7_c6_rr2 + t2_r7_c6_rr3;

  assign t4_r7_c6_rr0 = t3_r7_c6_rr0 + t3_r7_c6_rr1;

  assign c_7_6 = t4_r7_c6_rr0;
  assign t0_r7_c7_rr0 = a_7_0 * b_0_7;
  assign t0_r7_c7_rr1 = a_7_1 * b_1_7;
  assign t0_r7_c7_rr2 = a_7_2 * b_2_7;
  assign t0_r7_c7_rr3 = a_7_3 * b_3_7;
  assign t0_r7_c7_rr4 = a_7_4 * b_4_7;
  assign t0_r7_c7_rr5 = a_7_5 * b_5_7;
  assign t0_r7_c7_rr6 = a_7_6 * b_6_7;
  assign t0_r7_c7_rr7 = a_7_7 * b_7_7;
  assign t0_r7_c7_rr8 = a_7_8 * b_8_7;
  assign t0_r7_c7_rr9 = a_7_9 * b_9_7;
  assign t0_r7_c7_rr10 = a_7_10 * b_10_7;
  assign t0_r7_c7_rr11 = a_7_11 * b_11_7;
  assign t0_r7_c7_rr12 = a_7_12 * b_12_7;
  assign t0_r7_c7_rr13 = a_7_13 * b_13_7;
  assign t0_r7_c7_rr14 = a_7_14 * b_14_7;
  assign t1_r7_c7_rr0 = t0_r7_c7_rr0 + t0_r7_c7_rr1;
  assign t1_r7_c7_rr1 = t0_r7_c7_rr2 + t0_r7_c7_rr3;
  assign t1_r7_c7_rr2 = t0_r7_c7_rr4 + t0_r7_c7_rr5;
  assign t1_r7_c7_rr3 = t0_r7_c7_rr6 + t0_r7_c7_rr7;
  assign t1_r7_c7_rr4 = t0_r7_c7_rr8 + t0_r7_c7_rr9;
  assign t1_r7_c7_rr5 = t0_r7_c7_rr10 + t0_r7_c7_rr11;
  assign t1_r7_c7_rr6 = t0_r7_c7_rr12 + t0_r7_c7_rr13;
  assign t1_r7_c7_rr7 = t0_r7_c7_rr14;

  assign t2_r7_c7_rr0 = t1_r7_c7_rr0 + t1_r7_c7_rr1;
  assign t2_r7_c7_rr1 = t1_r7_c7_rr2 + t1_r7_c7_rr3;
  assign t2_r7_c7_rr2 = t1_r7_c7_rr4 + t1_r7_c7_rr5;
  assign t2_r7_c7_rr3 = t1_r7_c7_rr6 + t1_r7_c7_rr7;

  assign t3_r7_c7_rr0 = t2_r7_c7_rr0 + t2_r7_c7_rr1;
  assign t3_r7_c7_rr1 = t2_r7_c7_rr2 + t2_r7_c7_rr3;

  assign t4_r7_c7_rr0 = t3_r7_c7_rr0 + t3_r7_c7_rr1;

  assign c_7_7 = t4_r7_c7_rr0;
  assign t0_r7_c8_rr0 = a_7_0 * b_0_8;
  assign t0_r7_c8_rr1 = a_7_1 * b_1_8;
  assign t0_r7_c8_rr2 = a_7_2 * b_2_8;
  assign t0_r7_c8_rr3 = a_7_3 * b_3_8;
  assign t0_r7_c8_rr4 = a_7_4 * b_4_8;
  assign t0_r7_c8_rr5 = a_7_5 * b_5_8;
  assign t0_r7_c8_rr6 = a_7_6 * b_6_8;
  assign t0_r7_c8_rr7 = a_7_7 * b_7_8;
  assign t0_r7_c8_rr8 = a_7_8 * b_8_8;
  assign t0_r7_c8_rr9 = a_7_9 * b_9_8;
  assign t0_r7_c8_rr10 = a_7_10 * b_10_8;
  assign t0_r7_c8_rr11 = a_7_11 * b_11_8;
  assign t0_r7_c8_rr12 = a_7_12 * b_12_8;
  assign t0_r7_c8_rr13 = a_7_13 * b_13_8;
  assign t0_r7_c8_rr14 = a_7_14 * b_14_8;
  assign t1_r7_c8_rr0 = t0_r7_c8_rr0 + t0_r7_c8_rr1;
  assign t1_r7_c8_rr1 = t0_r7_c8_rr2 + t0_r7_c8_rr3;
  assign t1_r7_c8_rr2 = t0_r7_c8_rr4 + t0_r7_c8_rr5;
  assign t1_r7_c8_rr3 = t0_r7_c8_rr6 + t0_r7_c8_rr7;
  assign t1_r7_c8_rr4 = t0_r7_c8_rr8 + t0_r7_c8_rr9;
  assign t1_r7_c8_rr5 = t0_r7_c8_rr10 + t0_r7_c8_rr11;
  assign t1_r7_c8_rr6 = t0_r7_c8_rr12 + t0_r7_c8_rr13;
  assign t1_r7_c8_rr7 = t0_r7_c8_rr14;

  assign t2_r7_c8_rr0 = t1_r7_c8_rr0 + t1_r7_c8_rr1;
  assign t2_r7_c8_rr1 = t1_r7_c8_rr2 + t1_r7_c8_rr3;
  assign t2_r7_c8_rr2 = t1_r7_c8_rr4 + t1_r7_c8_rr5;
  assign t2_r7_c8_rr3 = t1_r7_c8_rr6 + t1_r7_c8_rr7;

  assign t3_r7_c8_rr0 = t2_r7_c8_rr0 + t2_r7_c8_rr1;
  assign t3_r7_c8_rr1 = t2_r7_c8_rr2 + t2_r7_c8_rr3;

  assign t4_r7_c8_rr0 = t3_r7_c8_rr0 + t3_r7_c8_rr1;

  assign c_7_8 = t4_r7_c8_rr0;
  assign t0_r7_c9_rr0 = a_7_0 * b_0_9;
  assign t0_r7_c9_rr1 = a_7_1 * b_1_9;
  assign t0_r7_c9_rr2 = a_7_2 * b_2_9;
  assign t0_r7_c9_rr3 = a_7_3 * b_3_9;
  assign t0_r7_c9_rr4 = a_7_4 * b_4_9;
  assign t0_r7_c9_rr5 = a_7_5 * b_5_9;
  assign t0_r7_c9_rr6 = a_7_6 * b_6_9;
  assign t0_r7_c9_rr7 = a_7_7 * b_7_9;
  assign t0_r7_c9_rr8 = a_7_8 * b_8_9;
  assign t0_r7_c9_rr9 = a_7_9 * b_9_9;
  assign t0_r7_c9_rr10 = a_7_10 * b_10_9;
  assign t0_r7_c9_rr11 = a_7_11 * b_11_9;
  assign t0_r7_c9_rr12 = a_7_12 * b_12_9;
  assign t0_r7_c9_rr13 = a_7_13 * b_13_9;
  assign t0_r7_c9_rr14 = a_7_14 * b_14_9;
  assign t1_r7_c9_rr0 = t0_r7_c9_rr0 + t0_r7_c9_rr1;
  assign t1_r7_c9_rr1 = t0_r7_c9_rr2 + t0_r7_c9_rr3;
  assign t1_r7_c9_rr2 = t0_r7_c9_rr4 + t0_r7_c9_rr5;
  assign t1_r7_c9_rr3 = t0_r7_c9_rr6 + t0_r7_c9_rr7;
  assign t1_r7_c9_rr4 = t0_r7_c9_rr8 + t0_r7_c9_rr9;
  assign t1_r7_c9_rr5 = t0_r7_c9_rr10 + t0_r7_c9_rr11;
  assign t1_r7_c9_rr6 = t0_r7_c9_rr12 + t0_r7_c9_rr13;
  assign t1_r7_c9_rr7 = t0_r7_c9_rr14;

  assign t2_r7_c9_rr0 = t1_r7_c9_rr0 + t1_r7_c9_rr1;
  assign t2_r7_c9_rr1 = t1_r7_c9_rr2 + t1_r7_c9_rr3;
  assign t2_r7_c9_rr2 = t1_r7_c9_rr4 + t1_r7_c9_rr5;
  assign t2_r7_c9_rr3 = t1_r7_c9_rr6 + t1_r7_c9_rr7;

  assign t3_r7_c9_rr0 = t2_r7_c9_rr0 + t2_r7_c9_rr1;
  assign t3_r7_c9_rr1 = t2_r7_c9_rr2 + t2_r7_c9_rr3;

  assign t4_r7_c9_rr0 = t3_r7_c9_rr0 + t3_r7_c9_rr1;

  assign c_7_9 = t4_r7_c9_rr0;
  assign t0_r7_c10_rr0 = a_7_0 * b_0_10;
  assign t0_r7_c10_rr1 = a_7_1 * b_1_10;
  assign t0_r7_c10_rr2 = a_7_2 * b_2_10;
  assign t0_r7_c10_rr3 = a_7_3 * b_3_10;
  assign t0_r7_c10_rr4 = a_7_4 * b_4_10;
  assign t0_r7_c10_rr5 = a_7_5 * b_5_10;
  assign t0_r7_c10_rr6 = a_7_6 * b_6_10;
  assign t0_r7_c10_rr7 = a_7_7 * b_7_10;
  assign t0_r7_c10_rr8 = a_7_8 * b_8_10;
  assign t0_r7_c10_rr9 = a_7_9 * b_9_10;
  assign t0_r7_c10_rr10 = a_7_10 * b_10_10;
  assign t0_r7_c10_rr11 = a_7_11 * b_11_10;
  assign t0_r7_c10_rr12 = a_7_12 * b_12_10;
  assign t0_r7_c10_rr13 = a_7_13 * b_13_10;
  assign t0_r7_c10_rr14 = a_7_14 * b_14_10;
  assign t1_r7_c10_rr0 = t0_r7_c10_rr0 + t0_r7_c10_rr1;
  assign t1_r7_c10_rr1 = t0_r7_c10_rr2 + t0_r7_c10_rr3;
  assign t1_r7_c10_rr2 = t0_r7_c10_rr4 + t0_r7_c10_rr5;
  assign t1_r7_c10_rr3 = t0_r7_c10_rr6 + t0_r7_c10_rr7;
  assign t1_r7_c10_rr4 = t0_r7_c10_rr8 + t0_r7_c10_rr9;
  assign t1_r7_c10_rr5 = t0_r7_c10_rr10 + t0_r7_c10_rr11;
  assign t1_r7_c10_rr6 = t0_r7_c10_rr12 + t0_r7_c10_rr13;
  assign t1_r7_c10_rr7 = t0_r7_c10_rr14;

  assign t2_r7_c10_rr0 = t1_r7_c10_rr0 + t1_r7_c10_rr1;
  assign t2_r7_c10_rr1 = t1_r7_c10_rr2 + t1_r7_c10_rr3;
  assign t2_r7_c10_rr2 = t1_r7_c10_rr4 + t1_r7_c10_rr5;
  assign t2_r7_c10_rr3 = t1_r7_c10_rr6 + t1_r7_c10_rr7;

  assign t3_r7_c10_rr0 = t2_r7_c10_rr0 + t2_r7_c10_rr1;
  assign t3_r7_c10_rr1 = t2_r7_c10_rr2 + t2_r7_c10_rr3;

  assign t4_r7_c10_rr0 = t3_r7_c10_rr0 + t3_r7_c10_rr1;

  assign c_7_10 = t4_r7_c10_rr0;
  assign t0_r7_c11_rr0 = a_7_0 * b_0_11;
  assign t0_r7_c11_rr1 = a_7_1 * b_1_11;
  assign t0_r7_c11_rr2 = a_7_2 * b_2_11;
  assign t0_r7_c11_rr3 = a_7_3 * b_3_11;
  assign t0_r7_c11_rr4 = a_7_4 * b_4_11;
  assign t0_r7_c11_rr5 = a_7_5 * b_5_11;
  assign t0_r7_c11_rr6 = a_7_6 * b_6_11;
  assign t0_r7_c11_rr7 = a_7_7 * b_7_11;
  assign t0_r7_c11_rr8 = a_7_8 * b_8_11;
  assign t0_r7_c11_rr9 = a_7_9 * b_9_11;
  assign t0_r7_c11_rr10 = a_7_10 * b_10_11;
  assign t0_r7_c11_rr11 = a_7_11 * b_11_11;
  assign t0_r7_c11_rr12 = a_7_12 * b_12_11;
  assign t0_r7_c11_rr13 = a_7_13 * b_13_11;
  assign t0_r7_c11_rr14 = a_7_14 * b_14_11;
  assign t1_r7_c11_rr0 = t0_r7_c11_rr0 + t0_r7_c11_rr1;
  assign t1_r7_c11_rr1 = t0_r7_c11_rr2 + t0_r7_c11_rr3;
  assign t1_r7_c11_rr2 = t0_r7_c11_rr4 + t0_r7_c11_rr5;
  assign t1_r7_c11_rr3 = t0_r7_c11_rr6 + t0_r7_c11_rr7;
  assign t1_r7_c11_rr4 = t0_r7_c11_rr8 + t0_r7_c11_rr9;
  assign t1_r7_c11_rr5 = t0_r7_c11_rr10 + t0_r7_c11_rr11;
  assign t1_r7_c11_rr6 = t0_r7_c11_rr12 + t0_r7_c11_rr13;
  assign t1_r7_c11_rr7 = t0_r7_c11_rr14;

  assign t2_r7_c11_rr0 = t1_r7_c11_rr0 + t1_r7_c11_rr1;
  assign t2_r7_c11_rr1 = t1_r7_c11_rr2 + t1_r7_c11_rr3;
  assign t2_r7_c11_rr2 = t1_r7_c11_rr4 + t1_r7_c11_rr5;
  assign t2_r7_c11_rr3 = t1_r7_c11_rr6 + t1_r7_c11_rr7;

  assign t3_r7_c11_rr0 = t2_r7_c11_rr0 + t2_r7_c11_rr1;
  assign t3_r7_c11_rr1 = t2_r7_c11_rr2 + t2_r7_c11_rr3;

  assign t4_r7_c11_rr0 = t3_r7_c11_rr0 + t3_r7_c11_rr1;

  assign c_7_11 = t4_r7_c11_rr0;
  assign t0_r7_c12_rr0 = a_7_0 * b_0_12;
  assign t0_r7_c12_rr1 = a_7_1 * b_1_12;
  assign t0_r7_c12_rr2 = a_7_2 * b_2_12;
  assign t0_r7_c12_rr3 = a_7_3 * b_3_12;
  assign t0_r7_c12_rr4 = a_7_4 * b_4_12;
  assign t0_r7_c12_rr5 = a_7_5 * b_5_12;
  assign t0_r7_c12_rr6 = a_7_6 * b_6_12;
  assign t0_r7_c12_rr7 = a_7_7 * b_7_12;
  assign t0_r7_c12_rr8 = a_7_8 * b_8_12;
  assign t0_r7_c12_rr9 = a_7_9 * b_9_12;
  assign t0_r7_c12_rr10 = a_7_10 * b_10_12;
  assign t0_r7_c12_rr11 = a_7_11 * b_11_12;
  assign t0_r7_c12_rr12 = a_7_12 * b_12_12;
  assign t0_r7_c12_rr13 = a_7_13 * b_13_12;
  assign t0_r7_c12_rr14 = a_7_14 * b_14_12;
  assign t1_r7_c12_rr0 = t0_r7_c12_rr0 + t0_r7_c12_rr1;
  assign t1_r7_c12_rr1 = t0_r7_c12_rr2 + t0_r7_c12_rr3;
  assign t1_r7_c12_rr2 = t0_r7_c12_rr4 + t0_r7_c12_rr5;
  assign t1_r7_c12_rr3 = t0_r7_c12_rr6 + t0_r7_c12_rr7;
  assign t1_r7_c12_rr4 = t0_r7_c12_rr8 + t0_r7_c12_rr9;
  assign t1_r7_c12_rr5 = t0_r7_c12_rr10 + t0_r7_c12_rr11;
  assign t1_r7_c12_rr6 = t0_r7_c12_rr12 + t0_r7_c12_rr13;
  assign t1_r7_c12_rr7 = t0_r7_c12_rr14;

  assign t2_r7_c12_rr0 = t1_r7_c12_rr0 + t1_r7_c12_rr1;
  assign t2_r7_c12_rr1 = t1_r7_c12_rr2 + t1_r7_c12_rr3;
  assign t2_r7_c12_rr2 = t1_r7_c12_rr4 + t1_r7_c12_rr5;
  assign t2_r7_c12_rr3 = t1_r7_c12_rr6 + t1_r7_c12_rr7;

  assign t3_r7_c12_rr0 = t2_r7_c12_rr0 + t2_r7_c12_rr1;
  assign t3_r7_c12_rr1 = t2_r7_c12_rr2 + t2_r7_c12_rr3;

  assign t4_r7_c12_rr0 = t3_r7_c12_rr0 + t3_r7_c12_rr1;

  assign c_7_12 = t4_r7_c12_rr0;
  assign t0_r7_c13_rr0 = a_7_0 * b_0_13;
  assign t0_r7_c13_rr1 = a_7_1 * b_1_13;
  assign t0_r7_c13_rr2 = a_7_2 * b_2_13;
  assign t0_r7_c13_rr3 = a_7_3 * b_3_13;
  assign t0_r7_c13_rr4 = a_7_4 * b_4_13;
  assign t0_r7_c13_rr5 = a_7_5 * b_5_13;
  assign t0_r7_c13_rr6 = a_7_6 * b_6_13;
  assign t0_r7_c13_rr7 = a_7_7 * b_7_13;
  assign t0_r7_c13_rr8 = a_7_8 * b_8_13;
  assign t0_r7_c13_rr9 = a_7_9 * b_9_13;
  assign t0_r7_c13_rr10 = a_7_10 * b_10_13;
  assign t0_r7_c13_rr11 = a_7_11 * b_11_13;
  assign t0_r7_c13_rr12 = a_7_12 * b_12_13;
  assign t0_r7_c13_rr13 = a_7_13 * b_13_13;
  assign t0_r7_c13_rr14 = a_7_14 * b_14_13;
  assign t1_r7_c13_rr0 = t0_r7_c13_rr0 + t0_r7_c13_rr1;
  assign t1_r7_c13_rr1 = t0_r7_c13_rr2 + t0_r7_c13_rr3;
  assign t1_r7_c13_rr2 = t0_r7_c13_rr4 + t0_r7_c13_rr5;
  assign t1_r7_c13_rr3 = t0_r7_c13_rr6 + t0_r7_c13_rr7;
  assign t1_r7_c13_rr4 = t0_r7_c13_rr8 + t0_r7_c13_rr9;
  assign t1_r7_c13_rr5 = t0_r7_c13_rr10 + t0_r7_c13_rr11;
  assign t1_r7_c13_rr6 = t0_r7_c13_rr12 + t0_r7_c13_rr13;
  assign t1_r7_c13_rr7 = t0_r7_c13_rr14;

  assign t2_r7_c13_rr0 = t1_r7_c13_rr0 + t1_r7_c13_rr1;
  assign t2_r7_c13_rr1 = t1_r7_c13_rr2 + t1_r7_c13_rr3;
  assign t2_r7_c13_rr2 = t1_r7_c13_rr4 + t1_r7_c13_rr5;
  assign t2_r7_c13_rr3 = t1_r7_c13_rr6 + t1_r7_c13_rr7;

  assign t3_r7_c13_rr0 = t2_r7_c13_rr0 + t2_r7_c13_rr1;
  assign t3_r7_c13_rr1 = t2_r7_c13_rr2 + t2_r7_c13_rr3;

  assign t4_r7_c13_rr0 = t3_r7_c13_rr0 + t3_r7_c13_rr1;

  assign c_7_13 = t4_r7_c13_rr0;
  assign t0_r7_c14_rr0 = a_7_0 * b_0_14;
  assign t0_r7_c14_rr1 = a_7_1 * b_1_14;
  assign t0_r7_c14_rr2 = a_7_2 * b_2_14;
  assign t0_r7_c14_rr3 = a_7_3 * b_3_14;
  assign t0_r7_c14_rr4 = a_7_4 * b_4_14;
  assign t0_r7_c14_rr5 = a_7_5 * b_5_14;
  assign t0_r7_c14_rr6 = a_7_6 * b_6_14;
  assign t0_r7_c14_rr7 = a_7_7 * b_7_14;
  assign t0_r7_c14_rr8 = a_7_8 * b_8_14;
  assign t0_r7_c14_rr9 = a_7_9 * b_9_14;
  assign t0_r7_c14_rr10 = a_7_10 * b_10_14;
  assign t0_r7_c14_rr11 = a_7_11 * b_11_14;
  assign t0_r7_c14_rr12 = a_7_12 * b_12_14;
  assign t0_r7_c14_rr13 = a_7_13 * b_13_14;
  assign t0_r7_c14_rr14 = a_7_14 * b_14_14;
  assign t1_r7_c14_rr0 = t0_r7_c14_rr0 + t0_r7_c14_rr1;
  assign t1_r7_c14_rr1 = t0_r7_c14_rr2 + t0_r7_c14_rr3;
  assign t1_r7_c14_rr2 = t0_r7_c14_rr4 + t0_r7_c14_rr5;
  assign t1_r7_c14_rr3 = t0_r7_c14_rr6 + t0_r7_c14_rr7;
  assign t1_r7_c14_rr4 = t0_r7_c14_rr8 + t0_r7_c14_rr9;
  assign t1_r7_c14_rr5 = t0_r7_c14_rr10 + t0_r7_c14_rr11;
  assign t1_r7_c14_rr6 = t0_r7_c14_rr12 + t0_r7_c14_rr13;
  assign t1_r7_c14_rr7 = t0_r7_c14_rr14;

  assign t2_r7_c14_rr0 = t1_r7_c14_rr0 + t1_r7_c14_rr1;
  assign t2_r7_c14_rr1 = t1_r7_c14_rr2 + t1_r7_c14_rr3;
  assign t2_r7_c14_rr2 = t1_r7_c14_rr4 + t1_r7_c14_rr5;
  assign t2_r7_c14_rr3 = t1_r7_c14_rr6 + t1_r7_c14_rr7;

  assign t3_r7_c14_rr0 = t2_r7_c14_rr0 + t2_r7_c14_rr1;
  assign t3_r7_c14_rr1 = t2_r7_c14_rr2 + t2_r7_c14_rr3;

  assign t4_r7_c14_rr0 = t3_r7_c14_rr0 + t3_r7_c14_rr1;

  assign c_7_14 = t4_r7_c14_rr0;
  assign t0_r8_c0_rr0 = a_8_0 * b_0_0;
  assign t0_r8_c0_rr1 = a_8_1 * b_1_0;
  assign t0_r8_c0_rr2 = a_8_2 * b_2_0;
  assign t0_r8_c0_rr3 = a_8_3 * b_3_0;
  assign t0_r8_c0_rr4 = a_8_4 * b_4_0;
  assign t0_r8_c0_rr5 = a_8_5 * b_5_0;
  assign t0_r8_c0_rr6 = a_8_6 * b_6_0;
  assign t0_r8_c0_rr7 = a_8_7 * b_7_0;
  assign t0_r8_c0_rr8 = a_8_8 * b_8_0;
  assign t0_r8_c0_rr9 = a_8_9 * b_9_0;
  assign t0_r8_c0_rr10 = a_8_10 * b_10_0;
  assign t0_r8_c0_rr11 = a_8_11 * b_11_0;
  assign t0_r8_c0_rr12 = a_8_12 * b_12_0;
  assign t0_r8_c0_rr13 = a_8_13 * b_13_0;
  assign t0_r8_c0_rr14 = a_8_14 * b_14_0;
  assign t1_r8_c0_rr0 = t0_r8_c0_rr0 + t0_r8_c0_rr1;
  assign t1_r8_c0_rr1 = t0_r8_c0_rr2 + t0_r8_c0_rr3;
  assign t1_r8_c0_rr2 = t0_r8_c0_rr4 + t0_r8_c0_rr5;
  assign t1_r8_c0_rr3 = t0_r8_c0_rr6 + t0_r8_c0_rr7;
  assign t1_r8_c0_rr4 = t0_r8_c0_rr8 + t0_r8_c0_rr9;
  assign t1_r8_c0_rr5 = t0_r8_c0_rr10 + t0_r8_c0_rr11;
  assign t1_r8_c0_rr6 = t0_r8_c0_rr12 + t0_r8_c0_rr13;
  assign t1_r8_c0_rr7 = t0_r8_c0_rr14;

  assign t2_r8_c0_rr0 = t1_r8_c0_rr0 + t1_r8_c0_rr1;
  assign t2_r8_c0_rr1 = t1_r8_c0_rr2 + t1_r8_c0_rr3;
  assign t2_r8_c0_rr2 = t1_r8_c0_rr4 + t1_r8_c0_rr5;
  assign t2_r8_c0_rr3 = t1_r8_c0_rr6 + t1_r8_c0_rr7;

  assign t3_r8_c0_rr0 = t2_r8_c0_rr0 + t2_r8_c0_rr1;
  assign t3_r8_c0_rr1 = t2_r8_c0_rr2 + t2_r8_c0_rr3;

  assign t4_r8_c0_rr0 = t3_r8_c0_rr0 + t3_r8_c0_rr1;

  assign c_8_0 = t4_r8_c0_rr0;
  assign t0_r8_c1_rr0 = a_8_0 * b_0_1;
  assign t0_r8_c1_rr1 = a_8_1 * b_1_1;
  assign t0_r8_c1_rr2 = a_8_2 * b_2_1;
  assign t0_r8_c1_rr3 = a_8_3 * b_3_1;
  assign t0_r8_c1_rr4 = a_8_4 * b_4_1;
  assign t0_r8_c1_rr5 = a_8_5 * b_5_1;
  assign t0_r8_c1_rr6 = a_8_6 * b_6_1;
  assign t0_r8_c1_rr7 = a_8_7 * b_7_1;
  assign t0_r8_c1_rr8 = a_8_8 * b_8_1;
  assign t0_r8_c1_rr9 = a_8_9 * b_9_1;
  assign t0_r8_c1_rr10 = a_8_10 * b_10_1;
  assign t0_r8_c1_rr11 = a_8_11 * b_11_1;
  assign t0_r8_c1_rr12 = a_8_12 * b_12_1;
  assign t0_r8_c1_rr13 = a_8_13 * b_13_1;
  assign t0_r8_c1_rr14 = a_8_14 * b_14_1;
  assign t1_r8_c1_rr0 = t0_r8_c1_rr0 + t0_r8_c1_rr1;
  assign t1_r8_c1_rr1 = t0_r8_c1_rr2 + t0_r8_c1_rr3;
  assign t1_r8_c1_rr2 = t0_r8_c1_rr4 + t0_r8_c1_rr5;
  assign t1_r8_c1_rr3 = t0_r8_c1_rr6 + t0_r8_c1_rr7;
  assign t1_r8_c1_rr4 = t0_r8_c1_rr8 + t0_r8_c1_rr9;
  assign t1_r8_c1_rr5 = t0_r8_c1_rr10 + t0_r8_c1_rr11;
  assign t1_r8_c1_rr6 = t0_r8_c1_rr12 + t0_r8_c1_rr13;
  assign t1_r8_c1_rr7 = t0_r8_c1_rr14;

  assign t2_r8_c1_rr0 = t1_r8_c1_rr0 + t1_r8_c1_rr1;
  assign t2_r8_c1_rr1 = t1_r8_c1_rr2 + t1_r8_c1_rr3;
  assign t2_r8_c1_rr2 = t1_r8_c1_rr4 + t1_r8_c1_rr5;
  assign t2_r8_c1_rr3 = t1_r8_c1_rr6 + t1_r8_c1_rr7;

  assign t3_r8_c1_rr0 = t2_r8_c1_rr0 + t2_r8_c1_rr1;
  assign t3_r8_c1_rr1 = t2_r8_c1_rr2 + t2_r8_c1_rr3;

  assign t4_r8_c1_rr0 = t3_r8_c1_rr0 + t3_r8_c1_rr1;

  assign c_8_1 = t4_r8_c1_rr0;
  assign t0_r8_c2_rr0 = a_8_0 * b_0_2;
  assign t0_r8_c2_rr1 = a_8_1 * b_1_2;
  assign t0_r8_c2_rr2 = a_8_2 * b_2_2;
  assign t0_r8_c2_rr3 = a_8_3 * b_3_2;
  assign t0_r8_c2_rr4 = a_8_4 * b_4_2;
  assign t0_r8_c2_rr5 = a_8_5 * b_5_2;
  assign t0_r8_c2_rr6 = a_8_6 * b_6_2;
  assign t0_r8_c2_rr7 = a_8_7 * b_7_2;
  assign t0_r8_c2_rr8 = a_8_8 * b_8_2;
  assign t0_r8_c2_rr9 = a_8_9 * b_9_2;
  assign t0_r8_c2_rr10 = a_8_10 * b_10_2;
  assign t0_r8_c2_rr11 = a_8_11 * b_11_2;
  assign t0_r8_c2_rr12 = a_8_12 * b_12_2;
  assign t0_r8_c2_rr13 = a_8_13 * b_13_2;
  assign t0_r8_c2_rr14 = a_8_14 * b_14_2;
  assign t1_r8_c2_rr0 = t0_r8_c2_rr0 + t0_r8_c2_rr1;
  assign t1_r8_c2_rr1 = t0_r8_c2_rr2 + t0_r8_c2_rr3;
  assign t1_r8_c2_rr2 = t0_r8_c2_rr4 + t0_r8_c2_rr5;
  assign t1_r8_c2_rr3 = t0_r8_c2_rr6 + t0_r8_c2_rr7;
  assign t1_r8_c2_rr4 = t0_r8_c2_rr8 + t0_r8_c2_rr9;
  assign t1_r8_c2_rr5 = t0_r8_c2_rr10 + t0_r8_c2_rr11;
  assign t1_r8_c2_rr6 = t0_r8_c2_rr12 + t0_r8_c2_rr13;
  assign t1_r8_c2_rr7 = t0_r8_c2_rr14;

  assign t2_r8_c2_rr0 = t1_r8_c2_rr0 + t1_r8_c2_rr1;
  assign t2_r8_c2_rr1 = t1_r8_c2_rr2 + t1_r8_c2_rr3;
  assign t2_r8_c2_rr2 = t1_r8_c2_rr4 + t1_r8_c2_rr5;
  assign t2_r8_c2_rr3 = t1_r8_c2_rr6 + t1_r8_c2_rr7;

  assign t3_r8_c2_rr0 = t2_r8_c2_rr0 + t2_r8_c2_rr1;
  assign t3_r8_c2_rr1 = t2_r8_c2_rr2 + t2_r8_c2_rr3;

  assign t4_r8_c2_rr0 = t3_r8_c2_rr0 + t3_r8_c2_rr1;

  assign c_8_2 = t4_r8_c2_rr0;
  assign t0_r8_c3_rr0 = a_8_0 * b_0_3;
  assign t0_r8_c3_rr1 = a_8_1 * b_1_3;
  assign t0_r8_c3_rr2 = a_8_2 * b_2_3;
  assign t0_r8_c3_rr3 = a_8_3 * b_3_3;
  assign t0_r8_c3_rr4 = a_8_4 * b_4_3;
  assign t0_r8_c3_rr5 = a_8_5 * b_5_3;
  assign t0_r8_c3_rr6 = a_8_6 * b_6_3;
  assign t0_r8_c3_rr7 = a_8_7 * b_7_3;
  assign t0_r8_c3_rr8 = a_8_8 * b_8_3;
  assign t0_r8_c3_rr9 = a_8_9 * b_9_3;
  assign t0_r8_c3_rr10 = a_8_10 * b_10_3;
  assign t0_r8_c3_rr11 = a_8_11 * b_11_3;
  assign t0_r8_c3_rr12 = a_8_12 * b_12_3;
  assign t0_r8_c3_rr13 = a_8_13 * b_13_3;
  assign t0_r8_c3_rr14 = a_8_14 * b_14_3;
  assign t1_r8_c3_rr0 = t0_r8_c3_rr0 + t0_r8_c3_rr1;
  assign t1_r8_c3_rr1 = t0_r8_c3_rr2 + t0_r8_c3_rr3;
  assign t1_r8_c3_rr2 = t0_r8_c3_rr4 + t0_r8_c3_rr5;
  assign t1_r8_c3_rr3 = t0_r8_c3_rr6 + t0_r8_c3_rr7;
  assign t1_r8_c3_rr4 = t0_r8_c3_rr8 + t0_r8_c3_rr9;
  assign t1_r8_c3_rr5 = t0_r8_c3_rr10 + t0_r8_c3_rr11;
  assign t1_r8_c3_rr6 = t0_r8_c3_rr12 + t0_r8_c3_rr13;
  assign t1_r8_c3_rr7 = t0_r8_c3_rr14;

  assign t2_r8_c3_rr0 = t1_r8_c3_rr0 + t1_r8_c3_rr1;
  assign t2_r8_c3_rr1 = t1_r8_c3_rr2 + t1_r8_c3_rr3;
  assign t2_r8_c3_rr2 = t1_r8_c3_rr4 + t1_r8_c3_rr5;
  assign t2_r8_c3_rr3 = t1_r8_c3_rr6 + t1_r8_c3_rr7;

  assign t3_r8_c3_rr0 = t2_r8_c3_rr0 + t2_r8_c3_rr1;
  assign t3_r8_c3_rr1 = t2_r8_c3_rr2 + t2_r8_c3_rr3;

  assign t4_r8_c3_rr0 = t3_r8_c3_rr0 + t3_r8_c3_rr1;

  assign c_8_3 = t4_r8_c3_rr0;
  assign t0_r8_c4_rr0 = a_8_0 * b_0_4;
  assign t0_r8_c4_rr1 = a_8_1 * b_1_4;
  assign t0_r8_c4_rr2 = a_8_2 * b_2_4;
  assign t0_r8_c4_rr3 = a_8_3 * b_3_4;
  assign t0_r8_c4_rr4 = a_8_4 * b_4_4;
  assign t0_r8_c4_rr5 = a_8_5 * b_5_4;
  assign t0_r8_c4_rr6 = a_8_6 * b_6_4;
  assign t0_r8_c4_rr7 = a_8_7 * b_7_4;
  assign t0_r8_c4_rr8 = a_8_8 * b_8_4;
  assign t0_r8_c4_rr9 = a_8_9 * b_9_4;
  assign t0_r8_c4_rr10 = a_8_10 * b_10_4;
  assign t0_r8_c4_rr11 = a_8_11 * b_11_4;
  assign t0_r8_c4_rr12 = a_8_12 * b_12_4;
  assign t0_r8_c4_rr13 = a_8_13 * b_13_4;
  assign t0_r8_c4_rr14 = a_8_14 * b_14_4;
  assign t1_r8_c4_rr0 = t0_r8_c4_rr0 + t0_r8_c4_rr1;
  assign t1_r8_c4_rr1 = t0_r8_c4_rr2 + t0_r8_c4_rr3;
  assign t1_r8_c4_rr2 = t0_r8_c4_rr4 + t0_r8_c4_rr5;
  assign t1_r8_c4_rr3 = t0_r8_c4_rr6 + t0_r8_c4_rr7;
  assign t1_r8_c4_rr4 = t0_r8_c4_rr8 + t0_r8_c4_rr9;
  assign t1_r8_c4_rr5 = t0_r8_c4_rr10 + t0_r8_c4_rr11;
  assign t1_r8_c4_rr6 = t0_r8_c4_rr12 + t0_r8_c4_rr13;
  assign t1_r8_c4_rr7 = t0_r8_c4_rr14;

  assign t2_r8_c4_rr0 = t1_r8_c4_rr0 + t1_r8_c4_rr1;
  assign t2_r8_c4_rr1 = t1_r8_c4_rr2 + t1_r8_c4_rr3;
  assign t2_r8_c4_rr2 = t1_r8_c4_rr4 + t1_r8_c4_rr5;
  assign t2_r8_c4_rr3 = t1_r8_c4_rr6 + t1_r8_c4_rr7;

  assign t3_r8_c4_rr0 = t2_r8_c4_rr0 + t2_r8_c4_rr1;
  assign t3_r8_c4_rr1 = t2_r8_c4_rr2 + t2_r8_c4_rr3;

  assign t4_r8_c4_rr0 = t3_r8_c4_rr0 + t3_r8_c4_rr1;

  assign c_8_4 = t4_r8_c4_rr0;
  assign t0_r8_c5_rr0 = a_8_0 * b_0_5;
  assign t0_r8_c5_rr1 = a_8_1 * b_1_5;
  assign t0_r8_c5_rr2 = a_8_2 * b_2_5;
  assign t0_r8_c5_rr3 = a_8_3 * b_3_5;
  assign t0_r8_c5_rr4 = a_8_4 * b_4_5;
  assign t0_r8_c5_rr5 = a_8_5 * b_5_5;
  assign t0_r8_c5_rr6 = a_8_6 * b_6_5;
  assign t0_r8_c5_rr7 = a_8_7 * b_7_5;
  assign t0_r8_c5_rr8 = a_8_8 * b_8_5;
  assign t0_r8_c5_rr9 = a_8_9 * b_9_5;
  assign t0_r8_c5_rr10 = a_8_10 * b_10_5;
  assign t0_r8_c5_rr11 = a_8_11 * b_11_5;
  assign t0_r8_c5_rr12 = a_8_12 * b_12_5;
  assign t0_r8_c5_rr13 = a_8_13 * b_13_5;
  assign t0_r8_c5_rr14 = a_8_14 * b_14_5;
  assign t1_r8_c5_rr0 = t0_r8_c5_rr0 + t0_r8_c5_rr1;
  assign t1_r8_c5_rr1 = t0_r8_c5_rr2 + t0_r8_c5_rr3;
  assign t1_r8_c5_rr2 = t0_r8_c5_rr4 + t0_r8_c5_rr5;
  assign t1_r8_c5_rr3 = t0_r8_c5_rr6 + t0_r8_c5_rr7;
  assign t1_r8_c5_rr4 = t0_r8_c5_rr8 + t0_r8_c5_rr9;
  assign t1_r8_c5_rr5 = t0_r8_c5_rr10 + t0_r8_c5_rr11;
  assign t1_r8_c5_rr6 = t0_r8_c5_rr12 + t0_r8_c5_rr13;
  assign t1_r8_c5_rr7 = t0_r8_c5_rr14;

  assign t2_r8_c5_rr0 = t1_r8_c5_rr0 + t1_r8_c5_rr1;
  assign t2_r8_c5_rr1 = t1_r8_c5_rr2 + t1_r8_c5_rr3;
  assign t2_r8_c5_rr2 = t1_r8_c5_rr4 + t1_r8_c5_rr5;
  assign t2_r8_c5_rr3 = t1_r8_c5_rr6 + t1_r8_c5_rr7;

  assign t3_r8_c5_rr0 = t2_r8_c5_rr0 + t2_r8_c5_rr1;
  assign t3_r8_c5_rr1 = t2_r8_c5_rr2 + t2_r8_c5_rr3;

  assign t4_r8_c5_rr0 = t3_r8_c5_rr0 + t3_r8_c5_rr1;

  assign c_8_5 = t4_r8_c5_rr0;
  assign t0_r8_c6_rr0 = a_8_0 * b_0_6;
  assign t0_r8_c6_rr1 = a_8_1 * b_1_6;
  assign t0_r8_c6_rr2 = a_8_2 * b_2_6;
  assign t0_r8_c6_rr3 = a_8_3 * b_3_6;
  assign t0_r8_c6_rr4 = a_8_4 * b_4_6;
  assign t0_r8_c6_rr5 = a_8_5 * b_5_6;
  assign t0_r8_c6_rr6 = a_8_6 * b_6_6;
  assign t0_r8_c6_rr7 = a_8_7 * b_7_6;
  assign t0_r8_c6_rr8 = a_8_8 * b_8_6;
  assign t0_r8_c6_rr9 = a_8_9 * b_9_6;
  assign t0_r8_c6_rr10 = a_8_10 * b_10_6;
  assign t0_r8_c6_rr11 = a_8_11 * b_11_6;
  assign t0_r8_c6_rr12 = a_8_12 * b_12_6;
  assign t0_r8_c6_rr13 = a_8_13 * b_13_6;
  assign t0_r8_c6_rr14 = a_8_14 * b_14_6;
  assign t1_r8_c6_rr0 = t0_r8_c6_rr0 + t0_r8_c6_rr1;
  assign t1_r8_c6_rr1 = t0_r8_c6_rr2 + t0_r8_c6_rr3;
  assign t1_r8_c6_rr2 = t0_r8_c6_rr4 + t0_r8_c6_rr5;
  assign t1_r8_c6_rr3 = t0_r8_c6_rr6 + t0_r8_c6_rr7;
  assign t1_r8_c6_rr4 = t0_r8_c6_rr8 + t0_r8_c6_rr9;
  assign t1_r8_c6_rr5 = t0_r8_c6_rr10 + t0_r8_c6_rr11;
  assign t1_r8_c6_rr6 = t0_r8_c6_rr12 + t0_r8_c6_rr13;
  assign t1_r8_c6_rr7 = t0_r8_c6_rr14;

  assign t2_r8_c6_rr0 = t1_r8_c6_rr0 + t1_r8_c6_rr1;
  assign t2_r8_c6_rr1 = t1_r8_c6_rr2 + t1_r8_c6_rr3;
  assign t2_r8_c6_rr2 = t1_r8_c6_rr4 + t1_r8_c6_rr5;
  assign t2_r8_c6_rr3 = t1_r8_c6_rr6 + t1_r8_c6_rr7;

  assign t3_r8_c6_rr0 = t2_r8_c6_rr0 + t2_r8_c6_rr1;
  assign t3_r8_c6_rr1 = t2_r8_c6_rr2 + t2_r8_c6_rr3;

  assign t4_r8_c6_rr0 = t3_r8_c6_rr0 + t3_r8_c6_rr1;

  assign c_8_6 = t4_r8_c6_rr0;
  assign t0_r8_c7_rr0 = a_8_0 * b_0_7;
  assign t0_r8_c7_rr1 = a_8_1 * b_1_7;
  assign t0_r8_c7_rr2 = a_8_2 * b_2_7;
  assign t0_r8_c7_rr3 = a_8_3 * b_3_7;
  assign t0_r8_c7_rr4 = a_8_4 * b_4_7;
  assign t0_r8_c7_rr5 = a_8_5 * b_5_7;
  assign t0_r8_c7_rr6 = a_8_6 * b_6_7;
  assign t0_r8_c7_rr7 = a_8_7 * b_7_7;
  assign t0_r8_c7_rr8 = a_8_8 * b_8_7;
  assign t0_r8_c7_rr9 = a_8_9 * b_9_7;
  assign t0_r8_c7_rr10 = a_8_10 * b_10_7;
  assign t0_r8_c7_rr11 = a_8_11 * b_11_7;
  assign t0_r8_c7_rr12 = a_8_12 * b_12_7;
  assign t0_r8_c7_rr13 = a_8_13 * b_13_7;
  assign t0_r8_c7_rr14 = a_8_14 * b_14_7;
  assign t1_r8_c7_rr0 = t0_r8_c7_rr0 + t0_r8_c7_rr1;
  assign t1_r8_c7_rr1 = t0_r8_c7_rr2 + t0_r8_c7_rr3;
  assign t1_r8_c7_rr2 = t0_r8_c7_rr4 + t0_r8_c7_rr5;
  assign t1_r8_c7_rr3 = t0_r8_c7_rr6 + t0_r8_c7_rr7;
  assign t1_r8_c7_rr4 = t0_r8_c7_rr8 + t0_r8_c7_rr9;
  assign t1_r8_c7_rr5 = t0_r8_c7_rr10 + t0_r8_c7_rr11;
  assign t1_r8_c7_rr6 = t0_r8_c7_rr12 + t0_r8_c7_rr13;
  assign t1_r8_c7_rr7 = t0_r8_c7_rr14;

  assign t2_r8_c7_rr0 = t1_r8_c7_rr0 + t1_r8_c7_rr1;
  assign t2_r8_c7_rr1 = t1_r8_c7_rr2 + t1_r8_c7_rr3;
  assign t2_r8_c7_rr2 = t1_r8_c7_rr4 + t1_r8_c7_rr5;
  assign t2_r8_c7_rr3 = t1_r8_c7_rr6 + t1_r8_c7_rr7;

  assign t3_r8_c7_rr0 = t2_r8_c7_rr0 + t2_r8_c7_rr1;
  assign t3_r8_c7_rr1 = t2_r8_c7_rr2 + t2_r8_c7_rr3;

  assign t4_r8_c7_rr0 = t3_r8_c7_rr0 + t3_r8_c7_rr1;

  assign c_8_7 = t4_r8_c7_rr0;
  assign t0_r8_c8_rr0 = a_8_0 * b_0_8;
  assign t0_r8_c8_rr1 = a_8_1 * b_1_8;
  assign t0_r8_c8_rr2 = a_8_2 * b_2_8;
  assign t0_r8_c8_rr3 = a_8_3 * b_3_8;
  assign t0_r8_c8_rr4 = a_8_4 * b_4_8;
  assign t0_r8_c8_rr5 = a_8_5 * b_5_8;
  assign t0_r8_c8_rr6 = a_8_6 * b_6_8;
  assign t0_r8_c8_rr7 = a_8_7 * b_7_8;
  assign t0_r8_c8_rr8 = a_8_8 * b_8_8;
  assign t0_r8_c8_rr9 = a_8_9 * b_9_8;
  assign t0_r8_c8_rr10 = a_8_10 * b_10_8;
  assign t0_r8_c8_rr11 = a_8_11 * b_11_8;
  assign t0_r8_c8_rr12 = a_8_12 * b_12_8;
  assign t0_r8_c8_rr13 = a_8_13 * b_13_8;
  assign t0_r8_c8_rr14 = a_8_14 * b_14_8;
  assign t1_r8_c8_rr0 = t0_r8_c8_rr0 + t0_r8_c8_rr1;
  assign t1_r8_c8_rr1 = t0_r8_c8_rr2 + t0_r8_c8_rr3;
  assign t1_r8_c8_rr2 = t0_r8_c8_rr4 + t0_r8_c8_rr5;
  assign t1_r8_c8_rr3 = t0_r8_c8_rr6 + t0_r8_c8_rr7;
  assign t1_r8_c8_rr4 = t0_r8_c8_rr8 + t0_r8_c8_rr9;
  assign t1_r8_c8_rr5 = t0_r8_c8_rr10 + t0_r8_c8_rr11;
  assign t1_r8_c8_rr6 = t0_r8_c8_rr12 + t0_r8_c8_rr13;
  assign t1_r8_c8_rr7 = t0_r8_c8_rr14;

  assign t2_r8_c8_rr0 = t1_r8_c8_rr0 + t1_r8_c8_rr1;
  assign t2_r8_c8_rr1 = t1_r8_c8_rr2 + t1_r8_c8_rr3;
  assign t2_r8_c8_rr2 = t1_r8_c8_rr4 + t1_r8_c8_rr5;
  assign t2_r8_c8_rr3 = t1_r8_c8_rr6 + t1_r8_c8_rr7;

  assign t3_r8_c8_rr0 = t2_r8_c8_rr0 + t2_r8_c8_rr1;
  assign t3_r8_c8_rr1 = t2_r8_c8_rr2 + t2_r8_c8_rr3;

  assign t4_r8_c8_rr0 = t3_r8_c8_rr0 + t3_r8_c8_rr1;

  assign c_8_8 = t4_r8_c8_rr0;
  assign t0_r8_c9_rr0 = a_8_0 * b_0_9;
  assign t0_r8_c9_rr1 = a_8_1 * b_1_9;
  assign t0_r8_c9_rr2 = a_8_2 * b_2_9;
  assign t0_r8_c9_rr3 = a_8_3 * b_3_9;
  assign t0_r8_c9_rr4 = a_8_4 * b_4_9;
  assign t0_r8_c9_rr5 = a_8_5 * b_5_9;
  assign t0_r8_c9_rr6 = a_8_6 * b_6_9;
  assign t0_r8_c9_rr7 = a_8_7 * b_7_9;
  assign t0_r8_c9_rr8 = a_8_8 * b_8_9;
  assign t0_r8_c9_rr9 = a_8_9 * b_9_9;
  assign t0_r8_c9_rr10 = a_8_10 * b_10_9;
  assign t0_r8_c9_rr11 = a_8_11 * b_11_9;
  assign t0_r8_c9_rr12 = a_8_12 * b_12_9;
  assign t0_r8_c9_rr13 = a_8_13 * b_13_9;
  assign t0_r8_c9_rr14 = a_8_14 * b_14_9;
  assign t1_r8_c9_rr0 = t0_r8_c9_rr0 + t0_r8_c9_rr1;
  assign t1_r8_c9_rr1 = t0_r8_c9_rr2 + t0_r8_c9_rr3;
  assign t1_r8_c9_rr2 = t0_r8_c9_rr4 + t0_r8_c9_rr5;
  assign t1_r8_c9_rr3 = t0_r8_c9_rr6 + t0_r8_c9_rr7;
  assign t1_r8_c9_rr4 = t0_r8_c9_rr8 + t0_r8_c9_rr9;
  assign t1_r8_c9_rr5 = t0_r8_c9_rr10 + t0_r8_c9_rr11;
  assign t1_r8_c9_rr6 = t0_r8_c9_rr12 + t0_r8_c9_rr13;
  assign t1_r8_c9_rr7 = t0_r8_c9_rr14;

  assign t2_r8_c9_rr0 = t1_r8_c9_rr0 + t1_r8_c9_rr1;
  assign t2_r8_c9_rr1 = t1_r8_c9_rr2 + t1_r8_c9_rr3;
  assign t2_r8_c9_rr2 = t1_r8_c9_rr4 + t1_r8_c9_rr5;
  assign t2_r8_c9_rr3 = t1_r8_c9_rr6 + t1_r8_c9_rr7;

  assign t3_r8_c9_rr0 = t2_r8_c9_rr0 + t2_r8_c9_rr1;
  assign t3_r8_c9_rr1 = t2_r8_c9_rr2 + t2_r8_c9_rr3;

  assign t4_r8_c9_rr0 = t3_r8_c9_rr0 + t3_r8_c9_rr1;

  assign c_8_9 = t4_r8_c9_rr0;
  assign t0_r8_c10_rr0 = a_8_0 * b_0_10;
  assign t0_r8_c10_rr1 = a_8_1 * b_1_10;
  assign t0_r8_c10_rr2 = a_8_2 * b_2_10;
  assign t0_r8_c10_rr3 = a_8_3 * b_3_10;
  assign t0_r8_c10_rr4 = a_8_4 * b_4_10;
  assign t0_r8_c10_rr5 = a_8_5 * b_5_10;
  assign t0_r8_c10_rr6 = a_8_6 * b_6_10;
  assign t0_r8_c10_rr7 = a_8_7 * b_7_10;
  assign t0_r8_c10_rr8 = a_8_8 * b_8_10;
  assign t0_r8_c10_rr9 = a_8_9 * b_9_10;
  assign t0_r8_c10_rr10 = a_8_10 * b_10_10;
  assign t0_r8_c10_rr11 = a_8_11 * b_11_10;
  assign t0_r8_c10_rr12 = a_8_12 * b_12_10;
  assign t0_r8_c10_rr13 = a_8_13 * b_13_10;
  assign t0_r8_c10_rr14 = a_8_14 * b_14_10;
  assign t1_r8_c10_rr0 = t0_r8_c10_rr0 + t0_r8_c10_rr1;
  assign t1_r8_c10_rr1 = t0_r8_c10_rr2 + t0_r8_c10_rr3;
  assign t1_r8_c10_rr2 = t0_r8_c10_rr4 + t0_r8_c10_rr5;
  assign t1_r8_c10_rr3 = t0_r8_c10_rr6 + t0_r8_c10_rr7;
  assign t1_r8_c10_rr4 = t0_r8_c10_rr8 + t0_r8_c10_rr9;
  assign t1_r8_c10_rr5 = t0_r8_c10_rr10 + t0_r8_c10_rr11;
  assign t1_r8_c10_rr6 = t0_r8_c10_rr12 + t0_r8_c10_rr13;
  assign t1_r8_c10_rr7 = t0_r8_c10_rr14;

  assign t2_r8_c10_rr0 = t1_r8_c10_rr0 + t1_r8_c10_rr1;
  assign t2_r8_c10_rr1 = t1_r8_c10_rr2 + t1_r8_c10_rr3;
  assign t2_r8_c10_rr2 = t1_r8_c10_rr4 + t1_r8_c10_rr5;
  assign t2_r8_c10_rr3 = t1_r8_c10_rr6 + t1_r8_c10_rr7;

  assign t3_r8_c10_rr0 = t2_r8_c10_rr0 + t2_r8_c10_rr1;
  assign t3_r8_c10_rr1 = t2_r8_c10_rr2 + t2_r8_c10_rr3;

  assign t4_r8_c10_rr0 = t3_r8_c10_rr0 + t3_r8_c10_rr1;

  assign c_8_10 = t4_r8_c10_rr0;
  assign t0_r8_c11_rr0 = a_8_0 * b_0_11;
  assign t0_r8_c11_rr1 = a_8_1 * b_1_11;
  assign t0_r8_c11_rr2 = a_8_2 * b_2_11;
  assign t0_r8_c11_rr3 = a_8_3 * b_3_11;
  assign t0_r8_c11_rr4 = a_8_4 * b_4_11;
  assign t0_r8_c11_rr5 = a_8_5 * b_5_11;
  assign t0_r8_c11_rr6 = a_8_6 * b_6_11;
  assign t0_r8_c11_rr7 = a_8_7 * b_7_11;
  assign t0_r8_c11_rr8 = a_8_8 * b_8_11;
  assign t0_r8_c11_rr9 = a_8_9 * b_9_11;
  assign t0_r8_c11_rr10 = a_8_10 * b_10_11;
  assign t0_r8_c11_rr11 = a_8_11 * b_11_11;
  assign t0_r8_c11_rr12 = a_8_12 * b_12_11;
  assign t0_r8_c11_rr13 = a_8_13 * b_13_11;
  assign t0_r8_c11_rr14 = a_8_14 * b_14_11;
  assign t1_r8_c11_rr0 = t0_r8_c11_rr0 + t0_r8_c11_rr1;
  assign t1_r8_c11_rr1 = t0_r8_c11_rr2 + t0_r8_c11_rr3;
  assign t1_r8_c11_rr2 = t0_r8_c11_rr4 + t0_r8_c11_rr5;
  assign t1_r8_c11_rr3 = t0_r8_c11_rr6 + t0_r8_c11_rr7;
  assign t1_r8_c11_rr4 = t0_r8_c11_rr8 + t0_r8_c11_rr9;
  assign t1_r8_c11_rr5 = t0_r8_c11_rr10 + t0_r8_c11_rr11;
  assign t1_r8_c11_rr6 = t0_r8_c11_rr12 + t0_r8_c11_rr13;
  assign t1_r8_c11_rr7 = t0_r8_c11_rr14;

  assign t2_r8_c11_rr0 = t1_r8_c11_rr0 + t1_r8_c11_rr1;
  assign t2_r8_c11_rr1 = t1_r8_c11_rr2 + t1_r8_c11_rr3;
  assign t2_r8_c11_rr2 = t1_r8_c11_rr4 + t1_r8_c11_rr5;
  assign t2_r8_c11_rr3 = t1_r8_c11_rr6 + t1_r8_c11_rr7;

  assign t3_r8_c11_rr0 = t2_r8_c11_rr0 + t2_r8_c11_rr1;
  assign t3_r8_c11_rr1 = t2_r8_c11_rr2 + t2_r8_c11_rr3;

  assign t4_r8_c11_rr0 = t3_r8_c11_rr0 + t3_r8_c11_rr1;

  assign c_8_11 = t4_r8_c11_rr0;
  assign t0_r8_c12_rr0 = a_8_0 * b_0_12;
  assign t0_r8_c12_rr1 = a_8_1 * b_1_12;
  assign t0_r8_c12_rr2 = a_8_2 * b_2_12;
  assign t0_r8_c12_rr3 = a_8_3 * b_3_12;
  assign t0_r8_c12_rr4 = a_8_4 * b_4_12;
  assign t0_r8_c12_rr5 = a_8_5 * b_5_12;
  assign t0_r8_c12_rr6 = a_8_6 * b_6_12;
  assign t0_r8_c12_rr7 = a_8_7 * b_7_12;
  assign t0_r8_c12_rr8 = a_8_8 * b_8_12;
  assign t0_r8_c12_rr9 = a_8_9 * b_9_12;
  assign t0_r8_c12_rr10 = a_8_10 * b_10_12;
  assign t0_r8_c12_rr11 = a_8_11 * b_11_12;
  assign t0_r8_c12_rr12 = a_8_12 * b_12_12;
  assign t0_r8_c12_rr13 = a_8_13 * b_13_12;
  assign t0_r8_c12_rr14 = a_8_14 * b_14_12;
  assign t1_r8_c12_rr0 = t0_r8_c12_rr0 + t0_r8_c12_rr1;
  assign t1_r8_c12_rr1 = t0_r8_c12_rr2 + t0_r8_c12_rr3;
  assign t1_r8_c12_rr2 = t0_r8_c12_rr4 + t0_r8_c12_rr5;
  assign t1_r8_c12_rr3 = t0_r8_c12_rr6 + t0_r8_c12_rr7;
  assign t1_r8_c12_rr4 = t0_r8_c12_rr8 + t0_r8_c12_rr9;
  assign t1_r8_c12_rr5 = t0_r8_c12_rr10 + t0_r8_c12_rr11;
  assign t1_r8_c12_rr6 = t0_r8_c12_rr12 + t0_r8_c12_rr13;
  assign t1_r8_c12_rr7 = t0_r8_c12_rr14;

  assign t2_r8_c12_rr0 = t1_r8_c12_rr0 + t1_r8_c12_rr1;
  assign t2_r8_c12_rr1 = t1_r8_c12_rr2 + t1_r8_c12_rr3;
  assign t2_r8_c12_rr2 = t1_r8_c12_rr4 + t1_r8_c12_rr5;
  assign t2_r8_c12_rr3 = t1_r8_c12_rr6 + t1_r8_c12_rr7;

  assign t3_r8_c12_rr0 = t2_r8_c12_rr0 + t2_r8_c12_rr1;
  assign t3_r8_c12_rr1 = t2_r8_c12_rr2 + t2_r8_c12_rr3;

  assign t4_r8_c12_rr0 = t3_r8_c12_rr0 + t3_r8_c12_rr1;

  assign c_8_12 = t4_r8_c12_rr0;
  assign t0_r8_c13_rr0 = a_8_0 * b_0_13;
  assign t0_r8_c13_rr1 = a_8_1 * b_1_13;
  assign t0_r8_c13_rr2 = a_8_2 * b_2_13;
  assign t0_r8_c13_rr3 = a_8_3 * b_3_13;
  assign t0_r8_c13_rr4 = a_8_4 * b_4_13;
  assign t0_r8_c13_rr5 = a_8_5 * b_5_13;
  assign t0_r8_c13_rr6 = a_8_6 * b_6_13;
  assign t0_r8_c13_rr7 = a_8_7 * b_7_13;
  assign t0_r8_c13_rr8 = a_8_8 * b_8_13;
  assign t0_r8_c13_rr9 = a_8_9 * b_9_13;
  assign t0_r8_c13_rr10 = a_8_10 * b_10_13;
  assign t0_r8_c13_rr11 = a_8_11 * b_11_13;
  assign t0_r8_c13_rr12 = a_8_12 * b_12_13;
  assign t0_r8_c13_rr13 = a_8_13 * b_13_13;
  assign t0_r8_c13_rr14 = a_8_14 * b_14_13;
  assign t1_r8_c13_rr0 = t0_r8_c13_rr0 + t0_r8_c13_rr1;
  assign t1_r8_c13_rr1 = t0_r8_c13_rr2 + t0_r8_c13_rr3;
  assign t1_r8_c13_rr2 = t0_r8_c13_rr4 + t0_r8_c13_rr5;
  assign t1_r8_c13_rr3 = t0_r8_c13_rr6 + t0_r8_c13_rr7;
  assign t1_r8_c13_rr4 = t0_r8_c13_rr8 + t0_r8_c13_rr9;
  assign t1_r8_c13_rr5 = t0_r8_c13_rr10 + t0_r8_c13_rr11;
  assign t1_r8_c13_rr6 = t0_r8_c13_rr12 + t0_r8_c13_rr13;
  assign t1_r8_c13_rr7 = t0_r8_c13_rr14;

  assign t2_r8_c13_rr0 = t1_r8_c13_rr0 + t1_r8_c13_rr1;
  assign t2_r8_c13_rr1 = t1_r8_c13_rr2 + t1_r8_c13_rr3;
  assign t2_r8_c13_rr2 = t1_r8_c13_rr4 + t1_r8_c13_rr5;
  assign t2_r8_c13_rr3 = t1_r8_c13_rr6 + t1_r8_c13_rr7;

  assign t3_r8_c13_rr0 = t2_r8_c13_rr0 + t2_r8_c13_rr1;
  assign t3_r8_c13_rr1 = t2_r8_c13_rr2 + t2_r8_c13_rr3;

  assign t4_r8_c13_rr0 = t3_r8_c13_rr0 + t3_r8_c13_rr1;

  assign c_8_13 = t4_r8_c13_rr0;
  assign t0_r8_c14_rr0 = a_8_0 * b_0_14;
  assign t0_r8_c14_rr1 = a_8_1 * b_1_14;
  assign t0_r8_c14_rr2 = a_8_2 * b_2_14;
  assign t0_r8_c14_rr3 = a_8_3 * b_3_14;
  assign t0_r8_c14_rr4 = a_8_4 * b_4_14;
  assign t0_r8_c14_rr5 = a_8_5 * b_5_14;
  assign t0_r8_c14_rr6 = a_8_6 * b_6_14;
  assign t0_r8_c14_rr7 = a_8_7 * b_7_14;
  assign t0_r8_c14_rr8 = a_8_8 * b_8_14;
  assign t0_r8_c14_rr9 = a_8_9 * b_9_14;
  assign t0_r8_c14_rr10 = a_8_10 * b_10_14;
  assign t0_r8_c14_rr11 = a_8_11 * b_11_14;
  assign t0_r8_c14_rr12 = a_8_12 * b_12_14;
  assign t0_r8_c14_rr13 = a_8_13 * b_13_14;
  assign t0_r8_c14_rr14 = a_8_14 * b_14_14;
  assign t1_r8_c14_rr0 = t0_r8_c14_rr0 + t0_r8_c14_rr1;
  assign t1_r8_c14_rr1 = t0_r8_c14_rr2 + t0_r8_c14_rr3;
  assign t1_r8_c14_rr2 = t0_r8_c14_rr4 + t0_r8_c14_rr5;
  assign t1_r8_c14_rr3 = t0_r8_c14_rr6 + t0_r8_c14_rr7;
  assign t1_r8_c14_rr4 = t0_r8_c14_rr8 + t0_r8_c14_rr9;
  assign t1_r8_c14_rr5 = t0_r8_c14_rr10 + t0_r8_c14_rr11;
  assign t1_r8_c14_rr6 = t0_r8_c14_rr12 + t0_r8_c14_rr13;
  assign t1_r8_c14_rr7 = t0_r8_c14_rr14;

  assign t2_r8_c14_rr0 = t1_r8_c14_rr0 + t1_r8_c14_rr1;
  assign t2_r8_c14_rr1 = t1_r8_c14_rr2 + t1_r8_c14_rr3;
  assign t2_r8_c14_rr2 = t1_r8_c14_rr4 + t1_r8_c14_rr5;
  assign t2_r8_c14_rr3 = t1_r8_c14_rr6 + t1_r8_c14_rr7;

  assign t3_r8_c14_rr0 = t2_r8_c14_rr0 + t2_r8_c14_rr1;
  assign t3_r8_c14_rr1 = t2_r8_c14_rr2 + t2_r8_c14_rr3;

  assign t4_r8_c14_rr0 = t3_r8_c14_rr0 + t3_r8_c14_rr1;

  assign c_8_14 = t4_r8_c14_rr0;
  assign t0_r9_c0_rr0 = a_9_0 * b_0_0;
  assign t0_r9_c0_rr1 = a_9_1 * b_1_0;
  assign t0_r9_c0_rr2 = a_9_2 * b_2_0;
  assign t0_r9_c0_rr3 = a_9_3 * b_3_0;
  assign t0_r9_c0_rr4 = a_9_4 * b_4_0;
  assign t0_r9_c0_rr5 = a_9_5 * b_5_0;
  assign t0_r9_c0_rr6 = a_9_6 * b_6_0;
  assign t0_r9_c0_rr7 = a_9_7 * b_7_0;
  assign t0_r9_c0_rr8 = a_9_8 * b_8_0;
  assign t0_r9_c0_rr9 = a_9_9 * b_9_0;
  assign t0_r9_c0_rr10 = a_9_10 * b_10_0;
  assign t0_r9_c0_rr11 = a_9_11 * b_11_0;
  assign t0_r9_c0_rr12 = a_9_12 * b_12_0;
  assign t0_r9_c0_rr13 = a_9_13 * b_13_0;
  assign t0_r9_c0_rr14 = a_9_14 * b_14_0;
  assign t1_r9_c0_rr0 = t0_r9_c0_rr0 + t0_r9_c0_rr1;
  assign t1_r9_c0_rr1 = t0_r9_c0_rr2 + t0_r9_c0_rr3;
  assign t1_r9_c0_rr2 = t0_r9_c0_rr4 + t0_r9_c0_rr5;
  assign t1_r9_c0_rr3 = t0_r9_c0_rr6 + t0_r9_c0_rr7;
  assign t1_r9_c0_rr4 = t0_r9_c0_rr8 + t0_r9_c0_rr9;
  assign t1_r9_c0_rr5 = t0_r9_c0_rr10 + t0_r9_c0_rr11;
  assign t1_r9_c0_rr6 = t0_r9_c0_rr12 + t0_r9_c0_rr13;
  assign t1_r9_c0_rr7 = t0_r9_c0_rr14;

  assign t2_r9_c0_rr0 = t1_r9_c0_rr0 + t1_r9_c0_rr1;
  assign t2_r9_c0_rr1 = t1_r9_c0_rr2 + t1_r9_c0_rr3;
  assign t2_r9_c0_rr2 = t1_r9_c0_rr4 + t1_r9_c0_rr5;
  assign t2_r9_c0_rr3 = t1_r9_c0_rr6 + t1_r9_c0_rr7;

  assign t3_r9_c0_rr0 = t2_r9_c0_rr0 + t2_r9_c0_rr1;
  assign t3_r9_c0_rr1 = t2_r9_c0_rr2 + t2_r9_c0_rr3;

  assign t4_r9_c0_rr0 = t3_r9_c0_rr0 + t3_r9_c0_rr1;

  assign c_9_0 = t4_r9_c0_rr0;
  assign t0_r9_c1_rr0 = a_9_0 * b_0_1;
  assign t0_r9_c1_rr1 = a_9_1 * b_1_1;
  assign t0_r9_c1_rr2 = a_9_2 * b_2_1;
  assign t0_r9_c1_rr3 = a_9_3 * b_3_1;
  assign t0_r9_c1_rr4 = a_9_4 * b_4_1;
  assign t0_r9_c1_rr5 = a_9_5 * b_5_1;
  assign t0_r9_c1_rr6 = a_9_6 * b_6_1;
  assign t0_r9_c1_rr7 = a_9_7 * b_7_1;
  assign t0_r9_c1_rr8 = a_9_8 * b_8_1;
  assign t0_r9_c1_rr9 = a_9_9 * b_9_1;
  assign t0_r9_c1_rr10 = a_9_10 * b_10_1;
  assign t0_r9_c1_rr11 = a_9_11 * b_11_1;
  assign t0_r9_c1_rr12 = a_9_12 * b_12_1;
  assign t0_r9_c1_rr13 = a_9_13 * b_13_1;
  assign t0_r9_c1_rr14 = a_9_14 * b_14_1;
  assign t1_r9_c1_rr0 = t0_r9_c1_rr0 + t0_r9_c1_rr1;
  assign t1_r9_c1_rr1 = t0_r9_c1_rr2 + t0_r9_c1_rr3;
  assign t1_r9_c1_rr2 = t0_r9_c1_rr4 + t0_r9_c1_rr5;
  assign t1_r9_c1_rr3 = t0_r9_c1_rr6 + t0_r9_c1_rr7;
  assign t1_r9_c1_rr4 = t0_r9_c1_rr8 + t0_r9_c1_rr9;
  assign t1_r9_c1_rr5 = t0_r9_c1_rr10 + t0_r9_c1_rr11;
  assign t1_r9_c1_rr6 = t0_r9_c1_rr12 + t0_r9_c1_rr13;
  assign t1_r9_c1_rr7 = t0_r9_c1_rr14;

  assign t2_r9_c1_rr0 = t1_r9_c1_rr0 + t1_r9_c1_rr1;
  assign t2_r9_c1_rr1 = t1_r9_c1_rr2 + t1_r9_c1_rr3;
  assign t2_r9_c1_rr2 = t1_r9_c1_rr4 + t1_r9_c1_rr5;
  assign t2_r9_c1_rr3 = t1_r9_c1_rr6 + t1_r9_c1_rr7;

  assign t3_r9_c1_rr0 = t2_r9_c1_rr0 + t2_r9_c1_rr1;
  assign t3_r9_c1_rr1 = t2_r9_c1_rr2 + t2_r9_c1_rr3;

  assign t4_r9_c1_rr0 = t3_r9_c1_rr0 + t3_r9_c1_rr1;

  assign c_9_1 = t4_r9_c1_rr0;
  assign t0_r9_c2_rr0 = a_9_0 * b_0_2;
  assign t0_r9_c2_rr1 = a_9_1 * b_1_2;
  assign t0_r9_c2_rr2 = a_9_2 * b_2_2;
  assign t0_r9_c2_rr3 = a_9_3 * b_3_2;
  assign t0_r9_c2_rr4 = a_9_4 * b_4_2;
  assign t0_r9_c2_rr5 = a_9_5 * b_5_2;
  assign t0_r9_c2_rr6 = a_9_6 * b_6_2;
  assign t0_r9_c2_rr7 = a_9_7 * b_7_2;
  assign t0_r9_c2_rr8 = a_9_8 * b_8_2;
  assign t0_r9_c2_rr9 = a_9_9 * b_9_2;
  assign t0_r9_c2_rr10 = a_9_10 * b_10_2;
  assign t0_r9_c2_rr11 = a_9_11 * b_11_2;
  assign t0_r9_c2_rr12 = a_9_12 * b_12_2;
  assign t0_r9_c2_rr13 = a_9_13 * b_13_2;
  assign t0_r9_c2_rr14 = a_9_14 * b_14_2;
  assign t1_r9_c2_rr0 = t0_r9_c2_rr0 + t0_r9_c2_rr1;
  assign t1_r9_c2_rr1 = t0_r9_c2_rr2 + t0_r9_c2_rr3;
  assign t1_r9_c2_rr2 = t0_r9_c2_rr4 + t0_r9_c2_rr5;
  assign t1_r9_c2_rr3 = t0_r9_c2_rr6 + t0_r9_c2_rr7;
  assign t1_r9_c2_rr4 = t0_r9_c2_rr8 + t0_r9_c2_rr9;
  assign t1_r9_c2_rr5 = t0_r9_c2_rr10 + t0_r9_c2_rr11;
  assign t1_r9_c2_rr6 = t0_r9_c2_rr12 + t0_r9_c2_rr13;
  assign t1_r9_c2_rr7 = t0_r9_c2_rr14;

  assign t2_r9_c2_rr0 = t1_r9_c2_rr0 + t1_r9_c2_rr1;
  assign t2_r9_c2_rr1 = t1_r9_c2_rr2 + t1_r9_c2_rr3;
  assign t2_r9_c2_rr2 = t1_r9_c2_rr4 + t1_r9_c2_rr5;
  assign t2_r9_c2_rr3 = t1_r9_c2_rr6 + t1_r9_c2_rr7;

  assign t3_r9_c2_rr0 = t2_r9_c2_rr0 + t2_r9_c2_rr1;
  assign t3_r9_c2_rr1 = t2_r9_c2_rr2 + t2_r9_c2_rr3;

  assign t4_r9_c2_rr0 = t3_r9_c2_rr0 + t3_r9_c2_rr1;

  assign c_9_2 = t4_r9_c2_rr0;
  assign t0_r9_c3_rr0 = a_9_0 * b_0_3;
  assign t0_r9_c3_rr1 = a_9_1 * b_1_3;
  assign t0_r9_c3_rr2 = a_9_2 * b_2_3;
  assign t0_r9_c3_rr3 = a_9_3 * b_3_3;
  assign t0_r9_c3_rr4 = a_9_4 * b_4_3;
  assign t0_r9_c3_rr5 = a_9_5 * b_5_3;
  assign t0_r9_c3_rr6 = a_9_6 * b_6_3;
  assign t0_r9_c3_rr7 = a_9_7 * b_7_3;
  assign t0_r9_c3_rr8 = a_9_8 * b_8_3;
  assign t0_r9_c3_rr9 = a_9_9 * b_9_3;
  assign t0_r9_c3_rr10 = a_9_10 * b_10_3;
  assign t0_r9_c3_rr11 = a_9_11 * b_11_3;
  assign t0_r9_c3_rr12 = a_9_12 * b_12_3;
  assign t0_r9_c3_rr13 = a_9_13 * b_13_3;
  assign t0_r9_c3_rr14 = a_9_14 * b_14_3;
  assign t1_r9_c3_rr0 = t0_r9_c3_rr0 + t0_r9_c3_rr1;
  assign t1_r9_c3_rr1 = t0_r9_c3_rr2 + t0_r9_c3_rr3;
  assign t1_r9_c3_rr2 = t0_r9_c3_rr4 + t0_r9_c3_rr5;
  assign t1_r9_c3_rr3 = t0_r9_c3_rr6 + t0_r9_c3_rr7;
  assign t1_r9_c3_rr4 = t0_r9_c3_rr8 + t0_r9_c3_rr9;
  assign t1_r9_c3_rr5 = t0_r9_c3_rr10 + t0_r9_c3_rr11;
  assign t1_r9_c3_rr6 = t0_r9_c3_rr12 + t0_r9_c3_rr13;
  assign t1_r9_c3_rr7 = t0_r9_c3_rr14;

  assign t2_r9_c3_rr0 = t1_r9_c3_rr0 + t1_r9_c3_rr1;
  assign t2_r9_c3_rr1 = t1_r9_c3_rr2 + t1_r9_c3_rr3;
  assign t2_r9_c3_rr2 = t1_r9_c3_rr4 + t1_r9_c3_rr5;
  assign t2_r9_c3_rr3 = t1_r9_c3_rr6 + t1_r9_c3_rr7;

  assign t3_r9_c3_rr0 = t2_r9_c3_rr0 + t2_r9_c3_rr1;
  assign t3_r9_c3_rr1 = t2_r9_c3_rr2 + t2_r9_c3_rr3;

  assign t4_r9_c3_rr0 = t3_r9_c3_rr0 + t3_r9_c3_rr1;

  assign c_9_3 = t4_r9_c3_rr0;
  assign t0_r9_c4_rr0 = a_9_0 * b_0_4;
  assign t0_r9_c4_rr1 = a_9_1 * b_1_4;
  assign t0_r9_c4_rr2 = a_9_2 * b_2_4;
  assign t0_r9_c4_rr3 = a_9_3 * b_3_4;
  assign t0_r9_c4_rr4 = a_9_4 * b_4_4;
  assign t0_r9_c4_rr5 = a_9_5 * b_5_4;
  assign t0_r9_c4_rr6 = a_9_6 * b_6_4;
  assign t0_r9_c4_rr7 = a_9_7 * b_7_4;
  assign t0_r9_c4_rr8 = a_9_8 * b_8_4;
  assign t0_r9_c4_rr9 = a_9_9 * b_9_4;
  assign t0_r9_c4_rr10 = a_9_10 * b_10_4;
  assign t0_r9_c4_rr11 = a_9_11 * b_11_4;
  assign t0_r9_c4_rr12 = a_9_12 * b_12_4;
  assign t0_r9_c4_rr13 = a_9_13 * b_13_4;
  assign t0_r9_c4_rr14 = a_9_14 * b_14_4;
  assign t1_r9_c4_rr0 = t0_r9_c4_rr0 + t0_r9_c4_rr1;
  assign t1_r9_c4_rr1 = t0_r9_c4_rr2 + t0_r9_c4_rr3;
  assign t1_r9_c4_rr2 = t0_r9_c4_rr4 + t0_r9_c4_rr5;
  assign t1_r9_c4_rr3 = t0_r9_c4_rr6 + t0_r9_c4_rr7;
  assign t1_r9_c4_rr4 = t0_r9_c4_rr8 + t0_r9_c4_rr9;
  assign t1_r9_c4_rr5 = t0_r9_c4_rr10 + t0_r9_c4_rr11;
  assign t1_r9_c4_rr6 = t0_r9_c4_rr12 + t0_r9_c4_rr13;
  assign t1_r9_c4_rr7 = t0_r9_c4_rr14;

  assign t2_r9_c4_rr0 = t1_r9_c4_rr0 + t1_r9_c4_rr1;
  assign t2_r9_c4_rr1 = t1_r9_c4_rr2 + t1_r9_c4_rr3;
  assign t2_r9_c4_rr2 = t1_r9_c4_rr4 + t1_r9_c4_rr5;
  assign t2_r9_c4_rr3 = t1_r9_c4_rr6 + t1_r9_c4_rr7;

  assign t3_r9_c4_rr0 = t2_r9_c4_rr0 + t2_r9_c4_rr1;
  assign t3_r9_c4_rr1 = t2_r9_c4_rr2 + t2_r9_c4_rr3;

  assign t4_r9_c4_rr0 = t3_r9_c4_rr0 + t3_r9_c4_rr1;

  assign c_9_4 = t4_r9_c4_rr0;
  assign t0_r9_c5_rr0 = a_9_0 * b_0_5;
  assign t0_r9_c5_rr1 = a_9_1 * b_1_5;
  assign t0_r9_c5_rr2 = a_9_2 * b_2_5;
  assign t0_r9_c5_rr3 = a_9_3 * b_3_5;
  assign t0_r9_c5_rr4 = a_9_4 * b_4_5;
  assign t0_r9_c5_rr5 = a_9_5 * b_5_5;
  assign t0_r9_c5_rr6 = a_9_6 * b_6_5;
  assign t0_r9_c5_rr7 = a_9_7 * b_7_5;
  assign t0_r9_c5_rr8 = a_9_8 * b_8_5;
  assign t0_r9_c5_rr9 = a_9_9 * b_9_5;
  assign t0_r9_c5_rr10 = a_9_10 * b_10_5;
  assign t0_r9_c5_rr11 = a_9_11 * b_11_5;
  assign t0_r9_c5_rr12 = a_9_12 * b_12_5;
  assign t0_r9_c5_rr13 = a_9_13 * b_13_5;
  assign t0_r9_c5_rr14 = a_9_14 * b_14_5;
  assign t1_r9_c5_rr0 = t0_r9_c5_rr0 + t0_r9_c5_rr1;
  assign t1_r9_c5_rr1 = t0_r9_c5_rr2 + t0_r9_c5_rr3;
  assign t1_r9_c5_rr2 = t0_r9_c5_rr4 + t0_r9_c5_rr5;
  assign t1_r9_c5_rr3 = t0_r9_c5_rr6 + t0_r9_c5_rr7;
  assign t1_r9_c5_rr4 = t0_r9_c5_rr8 + t0_r9_c5_rr9;
  assign t1_r9_c5_rr5 = t0_r9_c5_rr10 + t0_r9_c5_rr11;
  assign t1_r9_c5_rr6 = t0_r9_c5_rr12 + t0_r9_c5_rr13;
  assign t1_r9_c5_rr7 = t0_r9_c5_rr14;

  assign t2_r9_c5_rr0 = t1_r9_c5_rr0 + t1_r9_c5_rr1;
  assign t2_r9_c5_rr1 = t1_r9_c5_rr2 + t1_r9_c5_rr3;
  assign t2_r9_c5_rr2 = t1_r9_c5_rr4 + t1_r9_c5_rr5;
  assign t2_r9_c5_rr3 = t1_r9_c5_rr6 + t1_r9_c5_rr7;

  assign t3_r9_c5_rr0 = t2_r9_c5_rr0 + t2_r9_c5_rr1;
  assign t3_r9_c5_rr1 = t2_r9_c5_rr2 + t2_r9_c5_rr3;

  assign t4_r9_c5_rr0 = t3_r9_c5_rr0 + t3_r9_c5_rr1;

  assign c_9_5 = t4_r9_c5_rr0;
  assign t0_r9_c6_rr0 = a_9_0 * b_0_6;
  assign t0_r9_c6_rr1 = a_9_1 * b_1_6;
  assign t0_r9_c6_rr2 = a_9_2 * b_2_6;
  assign t0_r9_c6_rr3 = a_9_3 * b_3_6;
  assign t0_r9_c6_rr4 = a_9_4 * b_4_6;
  assign t0_r9_c6_rr5 = a_9_5 * b_5_6;
  assign t0_r9_c6_rr6 = a_9_6 * b_6_6;
  assign t0_r9_c6_rr7 = a_9_7 * b_7_6;
  assign t0_r9_c6_rr8 = a_9_8 * b_8_6;
  assign t0_r9_c6_rr9 = a_9_9 * b_9_6;
  assign t0_r9_c6_rr10 = a_9_10 * b_10_6;
  assign t0_r9_c6_rr11 = a_9_11 * b_11_6;
  assign t0_r9_c6_rr12 = a_9_12 * b_12_6;
  assign t0_r9_c6_rr13 = a_9_13 * b_13_6;
  assign t0_r9_c6_rr14 = a_9_14 * b_14_6;
  assign t1_r9_c6_rr0 = t0_r9_c6_rr0 + t0_r9_c6_rr1;
  assign t1_r9_c6_rr1 = t0_r9_c6_rr2 + t0_r9_c6_rr3;
  assign t1_r9_c6_rr2 = t0_r9_c6_rr4 + t0_r9_c6_rr5;
  assign t1_r9_c6_rr3 = t0_r9_c6_rr6 + t0_r9_c6_rr7;
  assign t1_r9_c6_rr4 = t0_r9_c6_rr8 + t0_r9_c6_rr9;
  assign t1_r9_c6_rr5 = t0_r9_c6_rr10 + t0_r9_c6_rr11;
  assign t1_r9_c6_rr6 = t0_r9_c6_rr12 + t0_r9_c6_rr13;
  assign t1_r9_c6_rr7 = t0_r9_c6_rr14;

  assign t2_r9_c6_rr0 = t1_r9_c6_rr0 + t1_r9_c6_rr1;
  assign t2_r9_c6_rr1 = t1_r9_c6_rr2 + t1_r9_c6_rr3;
  assign t2_r9_c6_rr2 = t1_r9_c6_rr4 + t1_r9_c6_rr5;
  assign t2_r9_c6_rr3 = t1_r9_c6_rr6 + t1_r9_c6_rr7;

  assign t3_r9_c6_rr0 = t2_r9_c6_rr0 + t2_r9_c6_rr1;
  assign t3_r9_c6_rr1 = t2_r9_c6_rr2 + t2_r9_c6_rr3;

  assign t4_r9_c6_rr0 = t3_r9_c6_rr0 + t3_r9_c6_rr1;

  assign c_9_6 = t4_r9_c6_rr0;
  assign t0_r9_c7_rr0 = a_9_0 * b_0_7;
  assign t0_r9_c7_rr1 = a_9_1 * b_1_7;
  assign t0_r9_c7_rr2 = a_9_2 * b_2_7;
  assign t0_r9_c7_rr3 = a_9_3 * b_3_7;
  assign t0_r9_c7_rr4 = a_9_4 * b_4_7;
  assign t0_r9_c7_rr5 = a_9_5 * b_5_7;
  assign t0_r9_c7_rr6 = a_9_6 * b_6_7;
  assign t0_r9_c7_rr7 = a_9_7 * b_7_7;
  assign t0_r9_c7_rr8 = a_9_8 * b_8_7;
  assign t0_r9_c7_rr9 = a_9_9 * b_9_7;
  assign t0_r9_c7_rr10 = a_9_10 * b_10_7;
  assign t0_r9_c7_rr11 = a_9_11 * b_11_7;
  assign t0_r9_c7_rr12 = a_9_12 * b_12_7;
  assign t0_r9_c7_rr13 = a_9_13 * b_13_7;
  assign t0_r9_c7_rr14 = a_9_14 * b_14_7;
  assign t1_r9_c7_rr0 = t0_r9_c7_rr0 + t0_r9_c7_rr1;
  assign t1_r9_c7_rr1 = t0_r9_c7_rr2 + t0_r9_c7_rr3;
  assign t1_r9_c7_rr2 = t0_r9_c7_rr4 + t0_r9_c7_rr5;
  assign t1_r9_c7_rr3 = t0_r9_c7_rr6 + t0_r9_c7_rr7;
  assign t1_r9_c7_rr4 = t0_r9_c7_rr8 + t0_r9_c7_rr9;
  assign t1_r9_c7_rr5 = t0_r9_c7_rr10 + t0_r9_c7_rr11;
  assign t1_r9_c7_rr6 = t0_r9_c7_rr12 + t0_r9_c7_rr13;
  assign t1_r9_c7_rr7 = t0_r9_c7_rr14;

  assign t2_r9_c7_rr0 = t1_r9_c7_rr0 + t1_r9_c7_rr1;
  assign t2_r9_c7_rr1 = t1_r9_c7_rr2 + t1_r9_c7_rr3;
  assign t2_r9_c7_rr2 = t1_r9_c7_rr4 + t1_r9_c7_rr5;
  assign t2_r9_c7_rr3 = t1_r9_c7_rr6 + t1_r9_c7_rr7;

  assign t3_r9_c7_rr0 = t2_r9_c7_rr0 + t2_r9_c7_rr1;
  assign t3_r9_c7_rr1 = t2_r9_c7_rr2 + t2_r9_c7_rr3;

  assign t4_r9_c7_rr0 = t3_r9_c7_rr0 + t3_r9_c7_rr1;

  assign c_9_7 = t4_r9_c7_rr0;
  assign t0_r9_c8_rr0 = a_9_0 * b_0_8;
  assign t0_r9_c8_rr1 = a_9_1 * b_1_8;
  assign t0_r9_c8_rr2 = a_9_2 * b_2_8;
  assign t0_r9_c8_rr3 = a_9_3 * b_3_8;
  assign t0_r9_c8_rr4 = a_9_4 * b_4_8;
  assign t0_r9_c8_rr5 = a_9_5 * b_5_8;
  assign t0_r9_c8_rr6 = a_9_6 * b_6_8;
  assign t0_r9_c8_rr7 = a_9_7 * b_7_8;
  assign t0_r9_c8_rr8 = a_9_8 * b_8_8;
  assign t0_r9_c8_rr9 = a_9_9 * b_9_8;
  assign t0_r9_c8_rr10 = a_9_10 * b_10_8;
  assign t0_r9_c8_rr11 = a_9_11 * b_11_8;
  assign t0_r9_c8_rr12 = a_9_12 * b_12_8;
  assign t0_r9_c8_rr13 = a_9_13 * b_13_8;
  assign t0_r9_c8_rr14 = a_9_14 * b_14_8;
  assign t1_r9_c8_rr0 = t0_r9_c8_rr0 + t0_r9_c8_rr1;
  assign t1_r9_c8_rr1 = t0_r9_c8_rr2 + t0_r9_c8_rr3;
  assign t1_r9_c8_rr2 = t0_r9_c8_rr4 + t0_r9_c8_rr5;
  assign t1_r9_c8_rr3 = t0_r9_c8_rr6 + t0_r9_c8_rr7;
  assign t1_r9_c8_rr4 = t0_r9_c8_rr8 + t0_r9_c8_rr9;
  assign t1_r9_c8_rr5 = t0_r9_c8_rr10 + t0_r9_c8_rr11;
  assign t1_r9_c8_rr6 = t0_r9_c8_rr12 + t0_r9_c8_rr13;
  assign t1_r9_c8_rr7 = t0_r9_c8_rr14;

  assign t2_r9_c8_rr0 = t1_r9_c8_rr0 + t1_r9_c8_rr1;
  assign t2_r9_c8_rr1 = t1_r9_c8_rr2 + t1_r9_c8_rr3;
  assign t2_r9_c8_rr2 = t1_r9_c8_rr4 + t1_r9_c8_rr5;
  assign t2_r9_c8_rr3 = t1_r9_c8_rr6 + t1_r9_c8_rr7;

  assign t3_r9_c8_rr0 = t2_r9_c8_rr0 + t2_r9_c8_rr1;
  assign t3_r9_c8_rr1 = t2_r9_c8_rr2 + t2_r9_c8_rr3;

  assign t4_r9_c8_rr0 = t3_r9_c8_rr0 + t3_r9_c8_rr1;

  assign c_9_8 = t4_r9_c8_rr0;
  assign t0_r9_c9_rr0 = a_9_0 * b_0_9;
  assign t0_r9_c9_rr1 = a_9_1 * b_1_9;
  assign t0_r9_c9_rr2 = a_9_2 * b_2_9;
  assign t0_r9_c9_rr3 = a_9_3 * b_3_9;
  assign t0_r9_c9_rr4 = a_9_4 * b_4_9;
  assign t0_r9_c9_rr5 = a_9_5 * b_5_9;
  assign t0_r9_c9_rr6 = a_9_6 * b_6_9;
  assign t0_r9_c9_rr7 = a_9_7 * b_7_9;
  assign t0_r9_c9_rr8 = a_9_8 * b_8_9;
  assign t0_r9_c9_rr9 = a_9_9 * b_9_9;
  assign t0_r9_c9_rr10 = a_9_10 * b_10_9;
  assign t0_r9_c9_rr11 = a_9_11 * b_11_9;
  assign t0_r9_c9_rr12 = a_9_12 * b_12_9;
  assign t0_r9_c9_rr13 = a_9_13 * b_13_9;
  assign t0_r9_c9_rr14 = a_9_14 * b_14_9;
  assign t1_r9_c9_rr0 = t0_r9_c9_rr0 + t0_r9_c9_rr1;
  assign t1_r9_c9_rr1 = t0_r9_c9_rr2 + t0_r9_c9_rr3;
  assign t1_r9_c9_rr2 = t0_r9_c9_rr4 + t0_r9_c9_rr5;
  assign t1_r9_c9_rr3 = t0_r9_c9_rr6 + t0_r9_c9_rr7;
  assign t1_r9_c9_rr4 = t0_r9_c9_rr8 + t0_r9_c9_rr9;
  assign t1_r9_c9_rr5 = t0_r9_c9_rr10 + t0_r9_c9_rr11;
  assign t1_r9_c9_rr6 = t0_r9_c9_rr12 + t0_r9_c9_rr13;
  assign t1_r9_c9_rr7 = t0_r9_c9_rr14;

  assign t2_r9_c9_rr0 = t1_r9_c9_rr0 + t1_r9_c9_rr1;
  assign t2_r9_c9_rr1 = t1_r9_c9_rr2 + t1_r9_c9_rr3;
  assign t2_r9_c9_rr2 = t1_r9_c9_rr4 + t1_r9_c9_rr5;
  assign t2_r9_c9_rr3 = t1_r9_c9_rr6 + t1_r9_c9_rr7;

  assign t3_r9_c9_rr0 = t2_r9_c9_rr0 + t2_r9_c9_rr1;
  assign t3_r9_c9_rr1 = t2_r9_c9_rr2 + t2_r9_c9_rr3;

  assign t4_r9_c9_rr0 = t3_r9_c9_rr0 + t3_r9_c9_rr1;

  assign c_9_9 = t4_r9_c9_rr0;
  assign t0_r9_c10_rr0 = a_9_0 * b_0_10;
  assign t0_r9_c10_rr1 = a_9_1 * b_1_10;
  assign t0_r9_c10_rr2 = a_9_2 * b_2_10;
  assign t0_r9_c10_rr3 = a_9_3 * b_3_10;
  assign t0_r9_c10_rr4 = a_9_4 * b_4_10;
  assign t0_r9_c10_rr5 = a_9_5 * b_5_10;
  assign t0_r9_c10_rr6 = a_9_6 * b_6_10;
  assign t0_r9_c10_rr7 = a_9_7 * b_7_10;
  assign t0_r9_c10_rr8 = a_9_8 * b_8_10;
  assign t0_r9_c10_rr9 = a_9_9 * b_9_10;
  assign t0_r9_c10_rr10 = a_9_10 * b_10_10;
  assign t0_r9_c10_rr11 = a_9_11 * b_11_10;
  assign t0_r9_c10_rr12 = a_9_12 * b_12_10;
  assign t0_r9_c10_rr13 = a_9_13 * b_13_10;
  assign t0_r9_c10_rr14 = a_9_14 * b_14_10;
  assign t1_r9_c10_rr0 = t0_r9_c10_rr0 + t0_r9_c10_rr1;
  assign t1_r9_c10_rr1 = t0_r9_c10_rr2 + t0_r9_c10_rr3;
  assign t1_r9_c10_rr2 = t0_r9_c10_rr4 + t0_r9_c10_rr5;
  assign t1_r9_c10_rr3 = t0_r9_c10_rr6 + t0_r9_c10_rr7;
  assign t1_r9_c10_rr4 = t0_r9_c10_rr8 + t0_r9_c10_rr9;
  assign t1_r9_c10_rr5 = t0_r9_c10_rr10 + t0_r9_c10_rr11;
  assign t1_r9_c10_rr6 = t0_r9_c10_rr12 + t0_r9_c10_rr13;
  assign t1_r9_c10_rr7 = t0_r9_c10_rr14;

  assign t2_r9_c10_rr0 = t1_r9_c10_rr0 + t1_r9_c10_rr1;
  assign t2_r9_c10_rr1 = t1_r9_c10_rr2 + t1_r9_c10_rr3;
  assign t2_r9_c10_rr2 = t1_r9_c10_rr4 + t1_r9_c10_rr5;
  assign t2_r9_c10_rr3 = t1_r9_c10_rr6 + t1_r9_c10_rr7;

  assign t3_r9_c10_rr0 = t2_r9_c10_rr0 + t2_r9_c10_rr1;
  assign t3_r9_c10_rr1 = t2_r9_c10_rr2 + t2_r9_c10_rr3;

  assign t4_r9_c10_rr0 = t3_r9_c10_rr0 + t3_r9_c10_rr1;

  assign c_9_10 = t4_r9_c10_rr0;
  assign t0_r9_c11_rr0 = a_9_0 * b_0_11;
  assign t0_r9_c11_rr1 = a_9_1 * b_1_11;
  assign t0_r9_c11_rr2 = a_9_2 * b_2_11;
  assign t0_r9_c11_rr3 = a_9_3 * b_3_11;
  assign t0_r9_c11_rr4 = a_9_4 * b_4_11;
  assign t0_r9_c11_rr5 = a_9_5 * b_5_11;
  assign t0_r9_c11_rr6 = a_9_6 * b_6_11;
  assign t0_r9_c11_rr7 = a_9_7 * b_7_11;
  assign t0_r9_c11_rr8 = a_9_8 * b_8_11;
  assign t0_r9_c11_rr9 = a_9_9 * b_9_11;
  assign t0_r9_c11_rr10 = a_9_10 * b_10_11;
  assign t0_r9_c11_rr11 = a_9_11 * b_11_11;
  assign t0_r9_c11_rr12 = a_9_12 * b_12_11;
  assign t0_r9_c11_rr13 = a_9_13 * b_13_11;
  assign t0_r9_c11_rr14 = a_9_14 * b_14_11;
  assign t1_r9_c11_rr0 = t0_r9_c11_rr0 + t0_r9_c11_rr1;
  assign t1_r9_c11_rr1 = t0_r9_c11_rr2 + t0_r9_c11_rr3;
  assign t1_r9_c11_rr2 = t0_r9_c11_rr4 + t0_r9_c11_rr5;
  assign t1_r9_c11_rr3 = t0_r9_c11_rr6 + t0_r9_c11_rr7;
  assign t1_r9_c11_rr4 = t0_r9_c11_rr8 + t0_r9_c11_rr9;
  assign t1_r9_c11_rr5 = t0_r9_c11_rr10 + t0_r9_c11_rr11;
  assign t1_r9_c11_rr6 = t0_r9_c11_rr12 + t0_r9_c11_rr13;
  assign t1_r9_c11_rr7 = t0_r9_c11_rr14;

  assign t2_r9_c11_rr0 = t1_r9_c11_rr0 + t1_r9_c11_rr1;
  assign t2_r9_c11_rr1 = t1_r9_c11_rr2 + t1_r9_c11_rr3;
  assign t2_r9_c11_rr2 = t1_r9_c11_rr4 + t1_r9_c11_rr5;
  assign t2_r9_c11_rr3 = t1_r9_c11_rr6 + t1_r9_c11_rr7;

  assign t3_r9_c11_rr0 = t2_r9_c11_rr0 + t2_r9_c11_rr1;
  assign t3_r9_c11_rr1 = t2_r9_c11_rr2 + t2_r9_c11_rr3;

  assign t4_r9_c11_rr0 = t3_r9_c11_rr0 + t3_r9_c11_rr1;

  assign c_9_11 = t4_r9_c11_rr0;
  assign t0_r9_c12_rr0 = a_9_0 * b_0_12;
  assign t0_r9_c12_rr1 = a_9_1 * b_1_12;
  assign t0_r9_c12_rr2 = a_9_2 * b_2_12;
  assign t0_r9_c12_rr3 = a_9_3 * b_3_12;
  assign t0_r9_c12_rr4 = a_9_4 * b_4_12;
  assign t0_r9_c12_rr5 = a_9_5 * b_5_12;
  assign t0_r9_c12_rr6 = a_9_6 * b_6_12;
  assign t0_r9_c12_rr7 = a_9_7 * b_7_12;
  assign t0_r9_c12_rr8 = a_9_8 * b_8_12;
  assign t0_r9_c12_rr9 = a_9_9 * b_9_12;
  assign t0_r9_c12_rr10 = a_9_10 * b_10_12;
  assign t0_r9_c12_rr11 = a_9_11 * b_11_12;
  assign t0_r9_c12_rr12 = a_9_12 * b_12_12;
  assign t0_r9_c12_rr13 = a_9_13 * b_13_12;
  assign t0_r9_c12_rr14 = a_9_14 * b_14_12;
  assign t1_r9_c12_rr0 = t0_r9_c12_rr0 + t0_r9_c12_rr1;
  assign t1_r9_c12_rr1 = t0_r9_c12_rr2 + t0_r9_c12_rr3;
  assign t1_r9_c12_rr2 = t0_r9_c12_rr4 + t0_r9_c12_rr5;
  assign t1_r9_c12_rr3 = t0_r9_c12_rr6 + t0_r9_c12_rr7;
  assign t1_r9_c12_rr4 = t0_r9_c12_rr8 + t0_r9_c12_rr9;
  assign t1_r9_c12_rr5 = t0_r9_c12_rr10 + t0_r9_c12_rr11;
  assign t1_r9_c12_rr6 = t0_r9_c12_rr12 + t0_r9_c12_rr13;
  assign t1_r9_c12_rr7 = t0_r9_c12_rr14;

  assign t2_r9_c12_rr0 = t1_r9_c12_rr0 + t1_r9_c12_rr1;
  assign t2_r9_c12_rr1 = t1_r9_c12_rr2 + t1_r9_c12_rr3;
  assign t2_r9_c12_rr2 = t1_r9_c12_rr4 + t1_r9_c12_rr5;
  assign t2_r9_c12_rr3 = t1_r9_c12_rr6 + t1_r9_c12_rr7;

  assign t3_r9_c12_rr0 = t2_r9_c12_rr0 + t2_r9_c12_rr1;
  assign t3_r9_c12_rr1 = t2_r9_c12_rr2 + t2_r9_c12_rr3;

  assign t4_r9_c12_rr0 = t3_r9_c12_rr0 + t3_r9_c12_rr1;

  assign c_9_12 = t4_r9_c12_rr0;
  assign t0_r9_c13_rr0 = a_9_0 * b_0_13;
  assign t0_r9_c13_rr1 = a_9_1 * b_1_13;
  assign t0_r9_c13_rr2 = a_9_2 * b_2_13;
  assign t0_r9_c13_rr3 = a_9_3 * b_3_13;
  assign t0_r9_c13_rr4 = a_9_4 * b_4_13;
  assign t0_r9_c13_rr5 = a_9_5 * b_5_13;
  assign t0_r9_c13_rr6 = a_9_6 * b_6_13;
  assign t0_r9_c13_rr7 = a_9_7 * b_7_13;
  assign t0_r9_c13_rr8 = a_9_8 * b_8_13;
  assign t0_r9_c13_rr9 = a_9_9 * b_9_13;
  assign t0_r9_c13_rr10 = a_9_10 * b_10_13;
  assign t0_r9_c13_rr11 = a_9_11 * b_11_13;
  assign t0_r9_c13_rr12 = a_9_12 * b_12_13;
  assign t0_r9_c13_rr13 = a_9_13 * b_13_13;
  assign t0_r9_c13_rr14 = a_9_14 * b_14_13;
  assign t1_r9_c13_rr0 = t0_r9_c13_rr0 + t0_r9_c13_rr1;
  assign t1_r9_c13_rr1 = t0_r9_c13_rr2 + t0_r9_c13_rr3;
  assign t1_r9_c13_rr2 = t0_r9_c13_rr4 + t0_r9_c13_rr5;
  assign t1_r9_c13_rr3 = t0_r9_c13_rr6 + t0_r9_c13_rr7;
  assign t1_r9_c13_rr4 = t0_r9_c13_rr8 + t0_r9_c13_rr9;
  assign t1_r9_c13_rr5 = t0_r9_c13_rr10 + t0_r9_c13_rr11;
  assign t1_r9_c13_rr6 = t0_r9_c13_rr12 + t0_r9_c13_rr13;
  assign t1_r9_c13_rr7 = t0_r9_c13_rr14;

  assign t2_r9_c13_rr0 = t1_r9_c13_rr0 + t1_r9_c13_rr1;
  assign t2_r9_c13_rr1 = t1_r9_c13_rr2 + t1_r9_c13_rr3;
  assign t2_r9_c13_rr2 = t1_r9_c13_rr4 + t1_r9_c13_rr5;
  assign t2_r9_c13_rr3 = t1_r9_c13_rr6 + t1_r9_c13_rr7;

  assign t3_r9_c13_rr0 = t2_r9_c13_rr0 + t2_r9_c13_rr1;
  assign t3_r9_c13_rr1 = t2_r9_c13_rr2 + t2_r9_c13_rr3;

  assign t4_r9_c13_rr0 = t3_r9_c13_rr0 + t3_r9_c13_rr1;

  assign c_9_13 = t4_r9_c13_rr0;
  assign t0_r9_c14_rr0 = a_9_0 * b_0_14;
  assign t0_r9_c14_rr1 = a_9_1 * b_1_14;
  assign t0_r9_c14_rr2 = a_9_2 * b_2_14;
  assign t0_r9_c14_rr3 = a_9_3 * b_3_14;
  assign t0_r9_c14_rr4 = a_9_4 * b_4_14;
  assign t0_r9_c14_rr5 = a_9_5 * b_5_14;
  assign t0_r9_c14_rr6 = a_9_6 * b_6_14;
  assign t0_r9_c14_rr7 = a_9_7 * b_7_14;
  assign t0_r9_c14_rr8 = a_9_8 * b_8_14;
  assign t0_r9_c14_rr9 = a_9_9 * b_9_14;
  assign t0_r9_c14_rr10 = a_9_10 * b_10_14;
  assign t0_r9_c14_rr11 = a_9_11 * b_11_14;
  assign t0_r9_c14_rr12 = a_9_12 * b_12_14;
  assign t0_r9_c14_rr13 = a_9_13 * b_13_14;
  assign t0_r9_c14_rr14 = a_9_14 * b_14_14;
  assign t1_r9_c14_rr0 = t0_r9_c14_rr0 + t0_r9_c14_rr1;
  assign t1_r9_c14_rr1 = t0_r9_c14_rr2 + t0_r9_c14_rr3;
  assign t1_r9_c14_rr2 = t0_r9_c14_rr4 + t0_r9_c14_rr5;
  assign t1_r9_c14_rr3 = t0_r9_c14_rr6 + t0_r9_c14_rr7;
  assign t1_r9_c14_rr4 = t0_r9_c14_rr8 + t0_r9_c14_rr9;
  assign t1_r9_c14_rr5 = t0_r9_c14_rr10 + t0_r9_c14_rr11;
  assign t1_r9_c14_rr6 = t0_r9_c14_rr12 + t0_r9_c14_rr13;
  assign t1_r9_c14_rr7 = t0_r9_c14_rr14;

  assign t2_r9_c14_rr0 = t1_r9_c14_rr0 + t1_r9_c14_rr1;
  assign t2_r9_c14_rr1 = t1_r9_c14_rr2 + t1_r9_c14_rr3;
  assign t2_r9_c14_rr2 = t1_r9_c14_rr4 + t1_r9_c14_rr5;
  assign t2_r9_c14_rr3 = t1_r9_c14_rr6 + t1_r9_c14_rr7;

  assign t3_r9_c14_rr0 = t2_r9_c14_rr0 + t2_r9_c14_rr1;
  assign t3_r9_c14_rr1 = t2_r9_c14_rr2 + t2_r9_c14_rr3;

  assign t4_r9_c14_rr0 = t3_r9_c14_rr0 + t3_r9_c14_rr1;

  assign c_9_14 = t4_r9_c14_rr0;
  assign t0_r10_c0_rr0 = a_10_0 * b_0_0;
  assign t0_r10_c0_rr1 = a_10_1 * b_1_0;
  assign t0_r10_c0_rr2 = a_10_2 * b_2_0;
  assign t0_r10_c0_rr3 = a_10_3 * b_3_0;
  assign t0_r10_c0_rr4 = a_10_4 * b_4_0;
  assign t0_r10_c0_rr5 = a_10_5 * b_5_0;
  assign t0_r10_c0_rr6 = a_10_6 * b_6_0;
  assign t0_r10_c0_rr7 = a_10_7 * b_7_0;
  assign t0_r10_c0_rr8 = a_10_8 * b_8_0;
  assign t0_r10_c0_rr9 = a_10_9 * b_9_0;
  assign t0_r10_c0_rr10 = a_10_10 * b_10_0;
  assign t0_r10_c0_rr11 = a_10_11 * b_11_0;
  assign t0_r10_c0_rr12 = a_10_12 * b_12_0;
  assign t0_r10_c0_rr13 = a_10_13 * b_13_0;
  assign t0_r10_c0_rr14 = a_10_14 * b_14_0;
  assign t1_r10_c0_rr0 = t0_r10_c0_rr0 + t0_r10_c0_rr1;
  assign t1_r10_c0_rr1 = t0_r10_c0_rr2 + t0_r10_c0_rr3;
  assign t1_r10_c0_rr2 = t0_r10_c0_rr4 + t0_r10_c0_rr5;
  assign t1_r10_c0_rr3 = t0_r10_c0_rr6 + t0_r10_c0_rr7;
  assign t1_r10_c0_rr4 = t0_r10_c0_rr8 + t0_r10_c0_rr9;
  assign t1_r10_c0_rr5 = t0_r10_c0_rr10 + t0_r10_c0_rr11;
  assign t1_r10_c0_rr6 = t0_r10_c0_rr12 + t0_r10_c0_rr13;
  assign t1_r10_c0_rr7 = t0_r10_c0_rr14;

  assign t2_r10_c0_rr0 = t1_r10_c0_rr0 + t1_r10_c0_rr1;
  assign t2_r10_c0_rr1 = t1_r10_c0_rr2 + t1_r10_c0_rr3;
  assign t2_r10_c0_rr2 = t1_r10_c0_rr4 + t1_r10_c0_rr5;
  assign t2_r10_c0_rr3 = t1_r10_c0_rr6 + t1_r10_c0_rr7;

  assign t3_r10_c0_rr0 = t2_r10_c0_rr0 + t2_r10_c0_rr1;
  assign t3_r10_c0_rr1 = t2_r10_c0_rr2 + t2_r10_c0_rr3;

  assign t4_r10_c0_rr0 = t3_r10_c0_rr0 + t3_r10_c0_rr1;

  assign c_10_0 = t4_r10_c0_rr0;
  assign t0_r10_c1_rr0 = a_10_0 * b_0_1;
  assign t0_r10_c1_rr1 = a_10_1 * b_1_1;
  assign t0_r10_c1_rr2 = a_10_2 * b_2_1;
  assign t0_r10_c1_rr3 = a_10_3 * b_3_1;
  assign t0_r10_c1_rr4 = a_10_4 * b_4_1;
  assign t0_r10_c1_rr5 = a_10_5 * b_5_1;
  assign t0_r10_c1_rr6 = a_10_6 * b_6_1;
  assign t0_r10_c1_rr7 = a_10_7 * b_7_1;
  assign t0_r10_c1_rr8 = a_10_8 * b_8_1;
  assign t0_r10_c1_rr9 = a_10_9 * b_9_1;
  assign t0_r10_c1_rr10 = a_10_10 * b_10_1;
  assign t0_r10_c1_rr11 = a_10_11 * b_11_1;
  assign t0_r10_c1_rr12 = a_10_12 * b_12_1;
  assign t0_r10_c1_rr13 = a_10_13 * b_13_1;
  assign t0_r10_c1_rr14 = a_10_14 * b_14_1;
  assign t1_r10_c1_rr0 = t0_r10_c1_rr0 + t0_r10_c1_rr1;
  assign t1_r10_c1_rr1 = t0_r10_c1_rr2 + t0_r10_c1_rr3;
  assign t1_r10_c1_rr2 = t0_r10_c1_rr4 + t0_r10_c1_rr5;
  assign t1_r10_c1_rr3 = t0_r10_c1_rr6 + t0_r10_c1_rr7;
  assign t1_r10_c1_rr4 = t0_r10_c1_rr8 + t0_r10_c1_rr9;
  assign t1_r10_c1_rr5 = t0_r10_c1_rr10 + t0_r10_c1_rr11;
  assign t1_r10_c1_rr6 = t0_r10_c1_rr12 + t0_r10_c1_rr13;
  assign t1_r10_c1_rr7 = t0_r10_c1_rr14;

  assign t2_r10_c1_rr0 = t1_r10_c1_rr0 + t1_r10_c1_rr1;
  assign t2_r10_c1_rr1 = t1_r10_c1_rr2 + t1_r10_c1_rr3;
  assign t2_r10_c1_rr2 = t1_r10_c1_rr4 + t1_r10_c1_rr5;
  assign t2_r10_c1_rr3 = t1_r10_c1_rr6 + t1_r10_c1_rr7;

  assign t3_r10_c1_rr0 = t2_r10_c1_rr0 + t2_r10_c1_rr1;
  assign t3_r10_c1_rr1 = t2_r10_c1_rr2 + t2_r10_c1_rr3;

  assign t4_r10_c1_rr0 = t3_r10_c1_rr0 + t3_r10_c1_rr1;

  assign c_10_1 = t4_r10_c1_rr0;
  assign t0_r10_c2_rr0 = a_10_0 * b_0_2;
  assign t0_r10_c2_rr1 = a_10_1 * b_1_2;
  assign t0_r10_c2_rr2 = a_10_2 * b_2_2;
  assign t0_r10_c2_rr3 = a_10_3 * b_3_2;
  assign t0_r10_c2_rr4 = a_10_4 * b_4_2;
  assign t0_r10_c2_rr5 = a_10_5 * b_5_2;
  assign t0_r10_c2_rr6 = a_10_6 * b_6_2;
  assign t0_r10_c2_rr7 = a_10_7 * b_7_2;
  assign t0_r10_c2_rr8 = a_10_8 * b_8_2;
  assign t0_r10_c2_rr9 = a_10_9 * b_9_2;
  assign t0_r10_c2_rr10 = a_10_10 * b_10_2;
  assign t0_r10_c2_rr11 = a_10_11 * b_11_2;
  assign t0_r10_c2_rr12 = a_10_12 * b_12_2;
  assign t0_r10_c2_rr13 = a_10_13 * b_13_2;
  assign t0_r10_c2_rr14 = a_10_14 * b_14_2;
  assign t1_r10_c2_rr0 = t0_r10_c2_rr0 + t0_r10_c2_rr1;
  assign t1_r10_c2_rr1 = t0_r10_c2_rr2 + t0_r10_c2_rr3;
  assign t1_r10_c2_rr2 = t0_r10_c2_rr4 + t0_r10_c2_rr5;
  assign t1_r10_c2_rr3 = t0_r10_c2_rr6 + t0_r10_c2_rr7;
  assign t1_r10_c2_rr4 = t0_r10_c2_rr8 + t0_r10_c2_rr9;
  assign t1_r10_c2_rr5 = t0_r10_c2_rr10 + t0_r10_c2_rr11;
  assign t1_r10_c2_rr6 = t0_r10_c2_rr12 + t0_r10_c2_rr13;
  assign t1_r10_c2_rr7 = t0_r10_c2_rr14;

  assign t2_r10_c2_rr0 = t1_r10_c2_rr0 + t1_r10_c2_rr1;
  assign t2_r10_c2_rr1 = t1_r10_c2_rr2 + t1_r10_c2_rr3;
  assign t2_r10_c2_rr2 = t1_r10_c2_rr4 + t1_r10_c2_rr5;
  assign t2_r10_c2_rr3 = t1_r10_c2_rr6 + t1_r10_c2_rr7;

  assign t3_r10_c2_rr0 = t2_r10_c2_rr0 + t2_r10_c2_rr1;
  assign t3_r10_c2_rr1 = t2_r10_c2_rr2 + t2_r10_c2_rr3;

  assign t4_r10_c2_rr0 = t3_r10_c2_rr0 + t3_r10_c2_rr1;

  assign c_10_2 = t4_r10_c2_rr0;
  assign t0_r10_c3_rr0 = a_10_0 * b_0_3;
  assign t0_r10_c3_rr1 = a_10_1 * b_1_3;
  assign t0_r10_c3_rr2 = a_10_2 * b_2_3;
  assign t0_r10_c3_rr3 = a_10_3 * b_3_3;
  assign t0_r10_c3_rr4 = a_10_4 * b_4_3;
  assign t0_r10_c3_rr5 = a_10_5 * b_5_3;
  assign t0_r10_c3_rr6 = a_10_6 * b_6_3;
  assign t0_r10_c3_rr7 = a_10_7 * b_7_3;
  assign t0_r10_c3_rr8 = a_10_8 * b_8_3;
  assign t0_r10_c3_rr9 = a_10_9 * b_9_3;
  assign t0_r10_c3_rr10 = a_10_10 * b_10_3;
  assign t0_r10_c3_rr11 = a_10_11 * b_11_3;
  assign t0_r10_c3_rr12 = a_10_12 * b_12_3;
  assign t0_r10_c3_rr13 = a_10_13 * b_13_3;
  assign t0_r10_c3_rr14 = a_10_14 * b_14_3;
  assign t1_r10_c3_rr0 = t0_r10_c3_rr0 + t0_r10_c3_rr1;
  assign t1_r10_c3_rr1 = t0_r10_c3_rr2 + t0_r10_c3_rr3;
  assign t1_r10_c3_rr2 = t0_r10_c3_rr4 + t0_r10_c3_rr5;
  assign t1_r10_c3_rr3 = t0_r10_c3_rr6 + t0_r10_c3_rr7;
  assign t1_r10_c3_rr4 = t0_r10_c3_rr8 + t0_r10_c3_rr9;
  assign t1_r10_c3_rr5 = t0_r10_c3_rr10 + t0_r10_c3_rr11;
  assign t1_r10_c3_rr6 = t0_r10_c3_rr12 + t0_r10_c3_rr13;
  assign t1_r10_c3_rr7 = t0_r10_c3_rr14;

  assign t2_r10_c3_rr0 = t1_r10_c3_rr0 + t1_r10_c3_rr1;
  assign t2_r10_c3_rr1 = t1_r10_c3_rr2 + t1_r10_c3_rr3;
  assign t2_r10_c3_rr2 = t1_r10_c3_rr4 + t1_r10_c3_rr5;
  assign t2_r10_c3_rr3 = t1_r10_c3_rr6 + t1_r10_c3_rr7;

  assign t3_r10_c3_rr0 = t2_r10_c3_rr0 + t2_r10_c3_rr1;
  assign t3_r10_c3_rr1 = t2_r10_c3_rr2 + t2_r10_c3_rr3;

  assign t4_r10_c3_rr0 = t3_r10_c3_rr0 + t3_r10_c3_rr1;

  assign c_10_3 = t4_r10_c3_rr0;
  assign t0_r10_c4_rr0 = a_10_0 * b_0_4;
  assign t0_r10_c4_rr1 = a_10_1 * b_1_4;
  assign t0_r10_c4_rr2 = a_10_2 * b_2_4;
  assign t0_r10_c4_rr3 = a_10_3 * b_3_4;
  assign t0_r10_c4_rr4 = a_10_4 * b_4_4;
  assign t0_r10_c4_rr5 = a_10_5 * b_5_4;
  assign t0_r10_c4_rr6 = a_10_6 * b_6_4;
  assign t0_r10_c4_rr7 = a_10_7 * b_7_4;
  assign t0_r10_c4_rr8 = a_10_8 * b_8_4;
  assign t0_r10_c4_rr9 = a_10_9 * b_9_4;
  assign t0_r10_c4_rr10 = a_10_10 * b_10_4;
  assign t0_r10_c4_rr11 = a_10_11 * b_11_4;
  assign t0_r10_c4_rr12 = a_10_12 * b_12_4;
  assign t0_r10_c4_rr13 = a_10_13 * b_13_4;
  assign t0_r10_c4_rr14 = a_10_14 * b_14_4;
  assign t1_r10_c4_rr0 = t0_r10_c4_rr0 + t0_r10_c4_rr1;
  assign t1_r10_c4_rr1 = t0_r10_c4_rr2 + t0_r10_c4_rr3;
  assign t1_r10_c4_rr2 = t0_r10_c4_rr4 + t0_r10_c4_rr5;
  assign t1_r10_c4_rr3 = t0_r10_c4_rr6 + t0_r10_c4_rr7;
  assign t1_r10_c4_rr4 = t0_r10_c4_rr8 + t0_r10_c4_rr9;
  assign t1_r10_c4_rr5 = t0_r10_c4_rr10 + t0_r10_c4_rr11;
  assign t1_r10_c4_rr6 = t0_r10_c4_rr12 + t0_r10_c4_rr13;
  assign t1_r10_c4_rr7 = t0_r10_c4_rr14;

  assign t2_r10_c4_rr0 = t1_r10_c4_rr0 + t1_r10_c4_rr1;
  assign t2_r10_c4_rr1 = t1_r10_c4_rr2 + t1_r10_c4_rr3;
  assign t2_r10_c4_rr2 = t1_r10_c4_rr4 + t1_r10_c4_rr5;
  assign t2_r10_c4_rr3 = t1_r10_c4_rr6 + t1_r10_c4_rr7;

  assign t3_r10_c4_rr0 = t2_r10_c4_rr0 + t2_r10_c4_rr1;
  assign t3_r10_c4_rr1 = t2_r10_c4_rr2 + t2_r10_c4_rr3;

  assign t4_r10_c4_rr0 = t3_r10_c4_rr0 + t3_r10_c4_rr1;

  assign c_10_4 = t4_r10_c4_rr0;
  assign t0_r10_c5_rr0 = a_10_0 * b_0_5;
  assign t0_r10_c5_rr1 = a_10_1 * b_1_5;
  assign t0_r10_c5_rr2 = a_10_2 * b_2_5;
  assign t0_r10_c5_rr3 = a_10_3 * b_3_5;
  assign t0_r10_c5_rr4 = a_10_4 * b_4_5;
  assign t0_r10_c5_rr5 = a_10_5 * b_5_5;
  assign t0_r10_c5_rr6 = a_10_6 * b_6_5;
  assign t0_r10_c5_rr7 = a_10_7 * b_7_5;
  assign t0_r10_c5_rr8 = a_10_8 * b_8_5;
  assign t0_r10_c5_rr9 = a_10_9 * b_9_5;
  assign t0_r10_c5_rr10 = a_10_10 * b_10_5;
  assign t0_r10_c5_rr11 = a_10_11 * b_11_5;
  assign t0_r10_c5_rr12 = a_10_12 * b_12_5;
  assign t0_r10_c5_rr13 = a_10_13 * b_13_5;
  assign t0_r10_c5_rr14 = a_10_14 * b_14_5;
  assign t1_r10_c5_rr0 = t0_r10_c5_rr0 + t0_r10_c5_rr1;
  assign t1_r10_c5_rr1 = t0_r10_c5_rr2 + t0_r10_c5_rr3;
  assign t1_r10_c5_rr2 = t0_r10_c5_rr4 + t0_r10_c5_rr5;
  assign t1_r10_c5_rr3 = t0_r10_c5_rr6 + t0_r10_c5_rr7;
  assign t1_r10_c5_rr4 = t0_r10_c5_rr8 + t0_r10_c5_rr9;
  assign t1_r10_c5_rr5 = t0_r10_c5_rr10 + t0_r10_c5_rr11;
  assign t1_r10_c5_rr6 = t0_r10_c5_rr12 + t0_r10_c5_rr13;
  assign t1_r10_c5_rr7 = t0_r10_c5_rr14;

  assign t2_r10_c5_rr0 = t1_r10_c5_rr0 + t1_r10_c5_rr1;
  assign t2_r10_c5_rr1 = t1_r10_c5_rr2 + t1_r10_c5_rr3;
  assign t2_r10_c5_rr2 = t1_r10_c5_rr4 + t1_r10_c5_rr5;
  assign t2_r10_c5_rr3 = t1_r10_c5_rr6 + t1_r10_c5_rr7;

  assign t3_r10_c5_rr0 = t2_r10_c5_rr0 + t2_r10_c5_rr1;
  assign t3_r10_c5_rr1 = t2_r10_c5_rr2 + t2_r10_c5_rr3;

  assign t4_r10_c5_rr0 = t3_r10_c5_rr0 + t3_r10_c5_rr1;

  assign c_10_5 = t4_r10_c5_rr0;
  assign t0_r10_c6_rr0 = a_10_0 * b_0_6;
  assign t0_r10_c6_rr1 = a_10_1 * b_1_6;
  assign t0_r10_c6_rr2 = a_10_2 * b_2_6;
  assign t0_r10_c6_rr3 = a_10_3 * b_3_6;
  assign t0_r10_c6_rr4 = a_10_4 * b_4_6;
  assign t0_r10_c6_rr5 = a_10_5 * b_5_6;
  assign t0_r10_c6_rr6 = a_10_6 * b_6_6;
  assign t0_r10_c6_rr7 = a_10_7 * b_7_6;
  assign t0_r10_c6_rr8 = a_10_8 * b_8_6;
  assign t0_r10_c6_rr9 = a_10_9 * b_9_6;
  assign t0_r10_c6_rr10 = a_10_10 * b_10_6;
  assign t0_r10_c6_rr11 = a_10_11 * b_11_6;
  assign t0_r10_c6_rr12 = a_10_12 * b_12_6;
  assign t0_r10_c6_rr13 = a_10_13 * b_13_6;
  assign t0_r10_c6_rr14 = a_10_14 * b_14_6;
  assign t1_r10_c6_rr0 = t0_r10_c6_rr0 + t0_r10_c6_rr1;
  assign t1_r10_c6_rr1 = t0_r10_c6_rr2 + t0_r10_c6_rr3;
  assign t1_r10_c6_rr2 = t0_r10_c6_rr4 + t0_r10_c6_rr5;
  assign t1_r10_c6_rr3 = t0_r10_c6_rr6 + t0_r10_c6_rr7;
  assign t1_r10_c6_rr4 = t0_r10_c6_rr8 + t0_r10_c6_rr9;
  assign t1_r10_c6_rr5 = t0_r10_c6_rr10 + t0_r10_c6_rr11;
  assign t1_r10_c6_rr6 = t0_r10_c6_rr12 + t0_r10_c6_rr13;
  assign t1_r10_c6_rr7 = t0_r10_c6_rr14;

  assign t2_r10_c6_rr0 = t1_r10_c6_rr0 + t1_r10_c6_rr1;
  assign t2_r10_c6_rr1 = t1_r10_c6_rr2 + t1_r10_c6_rr3;
  assign t2_r10_c6_rr2 = t1_r10_c6_rr4 + t1_r10_c6_rr5;
  assign t2_r10_c6_rr3 = t1_r10_c6_rr6 + t1_r10_c6_rr7;

  assign t3_r10_c6_rr0 = t2_r10_c6_rr0 + t2_r10_c6_rr1;
  assign t3_r10_c6_rr1 = t2_r10_c6_rr2 + t2_r10_c6_rr3;

  assign t4_r10_c6_rr0 = t3_r10_c6_rr0 + t3_r10_c6_rr1;

  assign c_10_6 = t4_r10_c6_rr0;
  assign t0_r10_c7_rr0 = a_10_0 * b_0_7;
  assign t0_r10_c7_rr1 = a_10_1 * b_1_7;
  assign t0_r10_c7_rr2 = a_10_2 * b_2_7;
  assign t0_r10_c7_rr3 = a_10_3 * b_3_7;
  assign t0_r10_c7_rr4 = a_10_4 * b_4_7;
  assign t0_r10_c7_rr5 = a_10_5 * b_5_7;
  assign t0_r10_c7_rr6 = a_10_6 * b_6_7;
  assign t0_r10_c7_rr7 = a_10_7 * b_7_7;
  assign t0_r10_c7_rr8 = a_10_8 * b_8_7;
  assign t0_r10_c7_rr9 = a_10_9 * b_9_7;
  assign t0_r10_c7_rr10 = a_10_10 * b_10_7;
  assign t0_r10_c7_rr11 = a_10_11 * b_11_7;
  assign t0_r10_c7_rr12 = a_10_12 * b_12_7;
  assign t0_r10_c7_rr13 = a_10_13 * b_13_7;
  assign t0_r10_c7_rr14 = a_10_14 * b_14_7;
  assign t1_r10_c7_rr0 = t0_r10_c7_rr0 + t0_r10_c7_rr1;
  assign t1_r10_c7_rr1 = t0_r10_c7_rr2 + t0_r10_c7_rr3;
  assign t1_r10_c7_rr2 = t0_r10_c7_rr4 + t0_r10_c7_rr5;
  assign t1_r10_c7_rr3 = t0_r10_c7_rr6 + t0_r10_c7_rr7;
  assign t1_r10_c7_rr4 = t0_r10_c7_rr8 + t0_r10_c7_rr9;
  assign t1_r10_c7_rr5 = t0_r10_c7_rr10 + t0_r10_c7_rr11;
  assign t1_r10_c7_rr6 = t0_r10_c7_rr12 + t0_r10_c7_rr13;
  assign t1_r10_c7_rr7 = t0_r10_c7_rr14;

  assign t2_r10_c7_rr0 = t1_r10_c7_rr0 + t1_r10_c7_rr1;
  assign t2_r10_c7_rr1 = t1_r10_c7_rr2 + t1_r10_c7_rr3;
  assign t2_r10_c7_rr2 = t1_r10_c7_rr4 + t1_r10_c7_rr5;
  assign t2_r10_c7_rr3 = t1_r10_c7_rr6 + t1_r10_c7_rr7;

  assign t3_r10_c7_rr0 = t2_r10_c7_rr0 + t2_r10_c7_rr1;
  assign t3_r10_c7_rr1 = t2_r10_c7_rr2 + t2_r10_c7_rr3;

  assign t4_r10_c7_rr0 = t3_r10_c7_rr0 + t3_r10_c7_rr1;

  assign c_10_7 = t4_r10_c7_rr0;
  assign t0_r10_c8_rr0 = a_10_0 * b_0_8;
  assign t0_r10_c8_rr1 = a_10_1 * b_1_8;
  assign t0_r10_c8_rr2 = a_10_2 * b_2_8;
  assign t0_r10_c8_rr3 = a_10_3 * b_3_8;
  assign t0_r10_c8_rr4 = a_10_4 * b_4_8;
  assign t0_r10_c8_rr5 = a_10_5 * b_5_8;
  assign t0_r10_c8_rr6 = a_10_6 * b_6_8;
  assign t0_r10_c8_rr7 = a_10_7 * b_7_8;
  assign t0_r10_c8_rr8 = a_10_8 * b_8_8;
  assign t0_r10_c8_rr9 = a_10_9 * b_9_8;
  assign t0_r10_c8_rr10 = a_10_10 * b_10_8;
  assign t0_r10_c8_rr11 = a_10_11 * b_11_8;
  assign t0_r10_c8_rr12 = a_10_12 * b_12_8;
  assign t0_r10_c8_rr13 = a_10_13 * b_13_8;
  assign t0_r10_c8_rr14 = a_10_14 * b_14_8;
  assign t1_r10_c8_rr0 = t0_r10_c8_rr0 + t0_r10_c8_rr1;
  assign t1_r10_c8_rr1 = t0_r10_c8_rr2 + t0_r10_c8_rr3;
  assign t1_r10_c8_rr2 = t0_r10_c8_rr4 + t0_r10_c8_rr5;
  assign t1_r10_c8_rr3 = t0_r10_c8_rr6 + t0_r10_c8_rr7;
  assign t1_r10_c8_rr4 = t0_r10_c8_rr8 + t0_r10_c8_rr9;
  assign t1_r10_c8_rr5 = t0_r10_c8_rr10 + t0_r10_c8_rr11;
  assign t1_r10_c8_rr6 = t0_r10_c8_rr12 + t0_r10_c8_rr13;
  assign t1_r10_c8_rr7 = t0_r10_c8_rr14;

  assign t2_r10_c8_rr0 = t1_r10_c8_rr0 + t1_r10_c8_rr1;
  assign t2_r10_c8_rr1 = t1_r10_c8_rr2 + t1_r10_c8_rr3;
  assign t2_r10_c8_rr2 = t1_r10_c8_rr4 + t1_r10_c8_rr5;
  assign t2_r10_c8_rr3 = t1_r10_c8_rr6 + t1_r10_c8_rr7;

  assign t3_r10_c8_rr0 = t2_r10_c8_rr0 + t2_r10_c8_rr1;
  assign t3_r10_c8_rr1 = t2_r10_c8_rr2 + t2_r10_c8_rr3;

  assign t4_r10_c8_rr0 = t3_r10_c8_rr0 + t3_r10_c8_rr1;

  assign c_10_8 = t4_r10_c8_rr0;
  assign t0_r10_c9_rr0 = a_10_0 * b_0_9;
  assign t0_r10_c9_rr1 = a_10_1 * b_1_9;
  assign t0_r10_c9_rr2 = a_10_2 * b_2_9;
  assign t0_r10_c9_rr3 = a_10_3 * b_3_9;
  assign t0_r10_c9_rr4 = a_10_4 * b_4_9;
  assign t0_r10_c9_rr5 = a_10_5 * b_5_9;
  assign t0_r10_c9_rr6 = a_10_6 * b_6_9;
  assign t0_r10_c9_rr7 = a_10_7 * b_7_9;
  assign t0_r10_c9_rr8 = a_10_8 * b_8_9;
  assign t0_r10_c9_rr9 = a_10_9 * b_9_9;
  assign t0_r10_c9_rr10 = a_10_10 * b_10_9;
  assign t0_r10_c9_rr11 = a_10_11 * b_11_9;
  assign t0_r10_c9_rr12 = a_10_12 * b_12_9;
  assign t0_r10_c9_rr13 = a_10_13 * b_13_9;
  assign t0_r10_c9_rr14 = a_10_14 * b_14_9;
  assign t1_r10_c9_rr0 = t0_r10_c9_rr0 + t0_r10_c9_rr1;
  assign t1_r10_c9_rr1 = t0_r10_c9_rr2 + t0_r10_c9_rr3;
  assign t1_r10_c9_rr2 = t0_r10_c9_rr4 + t0_r10_c9_rr5;
  assign t1_r10_c9_rr3 = t0_r10_c9_rr6 + t0_r10_c9_rr7;
  assign t1_r10_c9_rr4 = t0_r10_c9_rr8 + t0_r10_c9_rr9;
  assign t1_r10_c9_rr5 = t0_r10_c9_rr10 + t0_r10_c9_rr11;
  assign t1_r10_c9_rr6 = t0_r10_c9_rr12 + t0_r10_c9_rr13;
  assign t1_r10_c9_rr7 = t0_r10_c9_rr14;

  assign t2_r10_c9_rr0 = t1_r10_c9_rr0 + t1_r10_c9_rr1;
  assign t2_r10_c9_rr1 = t1_r10_c9_rr2 + t1_r10_c9_rr3;
  assign t2_r10_c9_rr2 = t1_r10_c9_rr4 + t1_r10_c9_rr5;
  assign t2_r10_c9_rr3 = t1_r10_c9_rr6 + t1_r10_c9_rr7;

  assign t3_r10_c9_rr0 = t2_r10_c9_rr0 + t2_r10_c9_rr1;
  assign t3_r10_c9_rr1 = t2_r10_c9_rr2 + t2_r10_c9_rr3;

  assign t4_r10_c9_rr0 = t3_r10_c9_rr0 + t3_r10_c9_rr1;

  assign c_10_9 = t4_r10_c9_rr0;
  assign t0_r10_c10_rr0 = a_10_0 * b_0_10;
  assign t0_r10_c10_rr1 = a_10_1 * b_1_10;
  assign t0_r10_c10_rr2 = a_10_2 * b_2_10;
  assign t0_r10_c10_rr3 = a_10_3 * b_3_10;
  assign t0_r10_c10_rr4 = a_10_4 * b_4_10;
  assign t0_r10_c10_rr5 = a_10_5 * b_5_10;
  assign t0_r10_c10_rr6 = a_10_6 * b_6_10;
  assign t0_r10_c10_rr7 = a_10_7 * b_7_10;
  assign t0_r10_c10_rr8 = a_10_8 * b_8_10;
  assign t0_r10_c10_rr9 = a_10_9 * b_9_10;
  assign t0_r10_c10_rr10 = a_10_10 * b_10_10;
  assign t0_r10_c10_rr11 = a_10_11 * b_11_10;
  assign t0_r10_c10_rr12 = a_10_12 * b_12_10;
  assign t0_r10_c10_rr13 = a_10_13 * b_13_10;
  assign t0_r10_c10_rr14 = a_10_14 * b_14_10;
  assign t1_r10_c10_rr0 = t0_r10_c10_rr0 + t0_r10_c10_rr1;
  assign t1_r10_c10_rr1 = t0_r10_c10_rr2 + t0_r10_c10_rr3;
  assign t1_r10_c10_rr2 = t0_r10_c10_rr4 + t0_r10_c10_rr5;
  assign t1_r10_c10_rr3 = t0_r10_c10_rr6 + t0_r10_c10_rr7;
  assign t1_r10_c10_rr4 = t0_r10_c10_rr8 + t0_r10_c10_rr9;
  assign t1_r10_c10_rr5 = t0_r10_c10_rr10 + t0_r10_c10_rr11;
  assign t1_r10_c10_rr6 = t0_r10_c10_rr12 + t0_r10_c10_rr13;
  assign t1_r10_c10_rr7 = t0_r10_c10_rr14;

  assign t2_r10_c10_rr0 = t1_r10_c10_rr0 + t1_r10_c10_rr1;
  assign t2_r10_c10_rr1 = t1_r10_c10_rr2 + t1_r10_c10_rr3;
  assign t2_r10_c10_rr2 = t1_r10_c10_rr4 + t1_r10_c10_rr5;
  assign t2_r10_c10_rr3 = t1_r10_c10_rr6 + t1_r10_c10_rr7;

  assign t3_r10_c10_rr0 = t2_r10_c10_rr0 + t2_r10_c10_rr1;
  assign t3_r10_c10_rr1 = t2_r10_c10_rr2 + t2_r10_c10_rr3;

  assign t4_r10_c10_rr0 = t3_r10_c10_rr0 + t3_r10_c10_rr1;

  assign c_10_10 = t4_r10_c10_rr0;
  assign t0_r10_c11_rr0 = a_10_0 * b_0_11;
  assign t0_r10_c11_rr1 = a_10_1 * b_1_11;
  assign t0_r10_c11_rr2 = a_10_2 * b_2_11;
  assign t0_r10_c11_rr3 = a_10_3 * b_3_11;
  assign t0_r10_c11_rr4 = a_10_4 * b_4_11;
  assign t0_r10_c11_rr5 = a_10_5 * b_5_11;
  assign t0_r10_c11_rr6 = a_10_6 * b_6_11;
  assign t0_r10_c11_rr7 = a_10_7 * b_7_11;
  assign t0_r10_c11_rr8 = a_10_8 * b_8_11;
  assign t0_r10_c11_rr9 = a_10_9 * b_9_11;
  assign t0_r10_c11_rr10 = a_10_10 * b_10_11;
  assign t0_r10_c11_rr11 = a_10_11 * b_11_11;
  assign t0_r10_c11_rr12 = a_10_12 * b_12_11;
  assign t0_r10_c11_rr13 = a_10_13 * b_13_11;
  assign t0_r10_c11_rr14 = a_10_14 * b_14_11;
  assign t1_r10_c11_rr0 = t0_r10_c11_rr0 + t0_r10_c11_rr1;
  assign t1_r10_c11_rr1 = t0_r10_c11_rr2 + t0_r10_c11_rr3;
  assign t1_r10_c11_rr2 = t0_r10_c11_rr4 + t0_r10_c11_rr5;
  assign t1_r10_c11_rr3 = t0_r10_c11_rr6 + t0_r10_c11_rr7;
  assign t1_r10_c11_rr4 = t0_r10_c11_rr8 + t0_r10_c11_rr9;
  assign t1_r10_c11_rr5 = t0_r10_c11_rr10 + t0_r10_c11_rr11;
  assign t1_r10_c11_rr6 = t0_r10_c11_rr12 + t0_r10_c11_rr13;
  assign t1_r10_c11_rr7 = t0_r10_c11_rr14;

  assign t2_r10_c11_rr0 = t1_r10_c11_rr0 + t1_r10_c11_rr1;
  assign t2_r10_c11_rr1 = t1_r10_c11_rr2 + t1_r10_c11_rr3;
  assign t2_r10_c11_rr2 = t1_r10_c11_rr4 + t1_r10_c11_rr5;
  assign t2_r10_c11_rr3 = t1_r10_c11_rr6 + t1_r10_c11_rr7;

  assign t3_r10_c11_rr0 = t2_r10_c11_rr0 + t2_r10_c11_rr1;
  assign t3_r10_c11_rr1 = t2_r10_c11_rr2 + t2_r10_c11_rr3;

  assign t4_r10_c11_rr0 = t3_r10_c11_rr0 + t3_r10_c11_rr1;

  assign c_10_11 = t4_r10_c11_rr0;
  assign t0_r10_c12_rr0 = a_10_0 * b_0_12;
  assign t0_r10_c12_rr1 = a_10_1 * b_1_12;
  assign t0_r10_c12_rr2 = a_10_2 * b_2_12;
  assign t0_r10_c12_rr3 = a_10_3 * b_3_12;
  assign t0_r10_c12_rr4 = a_10_4 * b_4_12;
  assign t0_r10_c12_rr5 = a_10_5 * b_5_12;
  assign t0_r10_c12_rr6 = a_10_6 * b_6_12;
  assign t0_r10_c12_rr7 = a_10_7 * b_7_12;
  assign t0_r10_c12_rr8 = a_10_8 * b_8_12;
  assign t0_r10_c12_rr9 = a_10_9 * b_9_12;
  assign t0_r10_c12_rr10 = a_10_10 * b_10_12;
  assign t0_r10_c12_rr11 = a_10_11 * b_11_12;
  assign t0_r10_c12_rr12 = a_10_12 * b_12_12;
  assign t0_r10_c12_rr13 = a_10_13 * b_13_12;
  assign t0_r10_c12_rr14 = a_10_14 * b_14_12;
  assign t1_r10_c12_rr0 = t0_r10_c12_rr0 + t0_r10_c12_rr1;
  assign t1_r10_c12_rr1 = t0_r10_c12_rr2 + t0_r10_c12_rr3;
  assign t1_r10_c12_rr2 = t0_r10_c12_rr4 + t0_r10_c12_rr5;
  assign t1_r10_c12_rr3 = t0_r10_c12_rr6 + t0_r10_c12_rr7;
  assign t1_r10_c12_rr4 = t0_r10_c12_rr8 + t0_r10_c12_rr9;
  assign t1_r10_c12_rr5 = t0_r10_c12_rr10 + t0_r10_c12_rr11;
  assign t1_r10_c12_rr6 = t0_r10_c12_rr12 + t0_r10_c12_rr13;
  assign t1_r10_c12_rr7 = t0_r10_c12_rr14;

  assign t2_r10_c12_rr0 = t1_r10_c12_rr0 + t1_r10_c12_rr1;
  assign t2_r10_c12_rr1 = t1_r10_c12_rr2 + t1_r10_c12_rr3;
  assign t2_r10_c12_rr2 = t1_r10_c12_rr4 + t1_r10_c12_rr5;
  assign t2_r10_c12_rr3 = t1_r10_c12_rr6 + t1_r10_c12_rr7;

  assign t3_r10_c12_rr0 = t2_r10_c12_rr0 + t2_r10_c12_rr1;
  assign t3_r10_c12_rr1 = t2_r10_c12_rr2 + t2_r10_c12_rr3;

  assign t4_r10_c12_rr0 = t3_r10_c12_rr0 + t3_r10_c12_rr1;

  assign c_10_12 = t4_r10_c12_rr0;
  assign t0_r10_c13_rr0 = a_10_0 * b_0_13;
  assign t0_r10_c13_rr1 = a_10_1 * b_1_13;
  assign t0_r10_c13_rr2 = a_10_2 * b_2_13;
  assign t0_r10_c13_rr3 = a_10_3 * b_3_13;
  assign t0_r10_c13_rr4 = a_10_4 * b_4_13;
  assign t0_r10_c13_rr5 = a_10_5 * b_5_13;
  assign t0_r10_c13_rr6 = a_10_6 * b_6_13;
  assign t0_r10_c13_rr7 = a_10_7 * b_7_13;
  assign t0_r10_c13_rr8 = a_10_8 * b_8_13;
  assign t0_r10_c13_rr9 = a_10_9 * b_9_13;
  assign t0_r10_c13_rr10 = a_10_10 * b_10_13;
  assign t0_r10_c13_rr11 = a_10_11 * b_11_13;
  assign t0_r10_c13_rr12 = a_10_12 * b_12_13;
  assign t0_r10_c13_rr13 = a_10_13 * b_13_13;
  assign t0_r10_c13_rr14 = a_10_14 * b_14_13;
  assign t1_r10_c13_rr0 = t0_r10_c13_rr0 + t0_r10_c13_rr1;
  assign t1_r10_c13_rr1 = t0_r10_c13_rr2 + t0_r10_c13_rr3;
  assign t1_r10_c13_rr2 = t0_r10_c13_rr4 + t0_r10_c13_rr5;
  assign t1_r10_c13_rr3 = t0_r10_c13_rr6 + t0_r10_c13_rr7;
  assign t1_r10_c13_rr4 = t0_r10_c13_rr8 + t0_r10_c13_rr9;
  assign t1_r10_c13_rr5 = t0_r10_c13_rr10 + t0_r10_c13_rr11;
  assign t1_r10_c13_rr6 = t0_r10_c13_rr12 + t0_r10_c13_rr13;
  assign t1_r10_c13_rr7 = t0_r10_c13_rr14;

  assign t2_r10_c13_rr0 = t1_r10_c13_rr0 + t1_r10_c13_rr1;
  assign t2_r10_c13_rr1 = t1_r10_c13_rr2 + t1_r10_c13_rr3;
  assign t2_r10_c13_rr2 = t1_r10_c13_rr4 + t1_r10_c13_rr5;
  assign t2_r10_c13_rr3 = t1_r10_c13_rr6 + t1_r10_c13_rr7;

  assign t3_r10_c13_rr0 = t2_r10_c13_rr0 + t2_r10_c13_rr1;
  assign t3_r10_c13_rr1 = t2_r10_c13_rr2 + t2_r10_c13_rr3;

  assign t4_r10_c13_rr0 = t3_r10_c13_rr0 + t3_r10_c13_rr1;

  assign c_10_13 = t4_r10_c13_rr0;
  assign t0_r10_c14_rr0 = a_10_0 * b_0_14;
  assign t0_r10_c14_rr1 = a_10_1 * b_1_14;
  assign t0_r10_c14_rr2 = a_10_2 * b_2_14;
  assign t0_r10_c14_rr3 = a_10_3 * b_3_14;
  assign t0_r10_c14_rr4 = a_10_4 * b_4_14;
  assign t0_r10_c14_rr5 = a_10_5 * b_5_14;
  assign t0_r10_c14_rr6 = a_10_6 * b_6_14;
  assign t0_r10_c14_rr7 = a_10_7 * b_7_14;
  assign t0_r10_c14_rr8 = a_10_8 * b_8_14;
  assign t0_r10_c14_rr9 = a_10_9 * b_9_14;
  assign t0_r10_c14_rr10 = a_10_10 * b_10_14;
  assign t0_r10_c14_rr11 = a_10_11 * b_11_14;
  assign t0_r10_c14_rr12 = a_10_12 * b_12_14;
  assign t0_r10_c14_rr13 = a_10_13 * b_13_14;
  assign t0_r10_c14_rr14 = a_10_14 * b_14_14;
  assign t1_r10_c14_rr0 = t0_r10_c14_rr0 + t0_r10_c14_rr1;
  assign t1_r10_c14_rr1 = t0_r10_c14_rr2 + t0_r10_c14_rr3;
  assign t1_r10_c14_rr2 = t0_r10_c14_rr4 + t0_r10_c14_rr5;
  assign t1_r10_c14_rr3 = t0_r10_c14_rr6 + t0_r10_c14_rr7;
  assign t1_r10_c14_rr4 = t0_r10_c14_rr8 + t0_r10_c14_rr9;
  assign t1_r10_c14_rr5 = t0_r10_c14_rr10 + t0_r10_c14_rr11;
  assign t1_r10_c14_rr6 = t0_r10_c14_rr12 + t0_r10_c14_rr13;
  assign t1_r10_c14_rr7 = t0_r10_c14_rr14;

  assign t2_r10_c14_rr0 = t1_r10_c14_rr0 + t1_r10_c14_rr1;
  assign t2_r10_c14_rr1 = t1_r10_c14_rr2 + t1_r10_c14_rr3;
  assign t2_r10_c14_rr2 = t1_r10_c14_rr4 + t1_r10_c14_rr5;
  assign t2_r10_c14_rr3 = t1_r10_c14_rr6 + t1_r10_c14_rr7;

  assign t3_r10_c14_rr0 = t2_r10_c14_rr0 + t2_r10_c14_rr1;
  assign t3_r10_c14_rr1 = t2_r10_c14_rr2 + t2_r10_c14_rr3;

  assign t4_r10_c14_rr0 = t3_r10_c14_rr0 + t3_r10_c14_rr1;

  assign c_10_14 = t4_r10_c14_rr0;
  assign t0_r11_c0_rr0 = a_11_0 * b_0_0;
  assign t0_r11_c0_rr1 = a_11_1 * b_1_0;
  assign t0_r11_c0_rr2 = a_11_2 * b_2_0;
  assign t0_r11_c0_rr3 = a_11_3 * b_3_0;
  assign t0_r11_c0_rr4 = a_11_4 * b_4_0;
  assign t0_r11_c0_rr5 = a_11_5 * b_5_0;
  assign t0_r11_c0_rr6 = a_11_6 * b_6_0;
  assign t0_r11_c0_rr7 = a_11_7 * b_7_0;
  assign t0_r11_c0_rr8 = a_11_8 * b_8_0;
  assign t0_r11_c0_rr9 = a_11_9 * b_9_0;
  assign t0_r11_c0_rr10 = a_11_10 * b_10_0;
  assign t0_r11_c0_rr11 = a_11_11 * b_11_0;
  assign t0_r11_c0_rr12 = a_11_12 * b_12_0;
  assign t0_r11_c0_rr13 = a_11_13 * b_13_0;
  assign t0_r11_c0_rr14 = a_11_14 * b_14_0;
  assign t1_r11_c0_rr0 = t0_r11_c0_rr0 + t0_r11_c0_rr1;
  assign t1_r11_c0_rr1 = t0_r11_c0_rr2 + t0_r11_c0_rr3;
  assign t1_r11_c0_rr2 = t0_r11_c0_rr4 + t0_r11_c0_rr5;
  assign t1_r11_c0_rr3 = t0_r11_c0_rr6 + t0_r11_c0_rr7;
  assign t1_r11_c0_rr4 = t0_r11_c0_rr8 + t0_r11_c0_rr9;
  assign t1_r11_c0_rr5 = t0_r11_c0_rr10 + t0_r11_c0_rr11;
  assign t1_r11_c0_rr6 = t0_r11_c0_rr12 + t0_r11_c0_rr13;
  assign t1_r11_c0_rr7 = t0_r11_c0_rr14;

  assign t2_r11_c0_rr0 = t1_r11_c0_rr0 + t1_r11_c0_rr1;
  assign t2_r11_c0_rr1 = t1_r11_c0_rr2 + t1_r11_c0_rr3;
  assign t2_r11_c0_rr2 = t1_r11_c0_rr4 + t1_r11_c0_rr5;
  assign t2_r11_c0_rr3 = t1_r11_c0_rr6 + t1_r11_c0_rr7;

  assign t3_r11_c0_rr0 = t2_r11_c0_rr0 + t2_r11_c0_rr1;
  assign t3_r11_c0_rr1 = t2_r11_c0_rr2 + t2_r11_c0_rr3;

  assign t4_r11_c0_rr0 = t3_r11_c0_rr0 + t3_r11_c0_rr1;

  assign c_11_0 = t4_r11_c0_rr0;
  assign t0_r11_c1_rr0 = a_11_0 * b_0_1;
  assign t0_r11_c1_rr1 = a_11_1 * b_1_1;
  assign t0_r11_c1_rr2 = a_11_2 * b_2_1;
  assign t0_r11_c1_rr3 = a_11_3 * b_3_1;
  assign t0_r11_c1_rr4 = a_11_4 * b_4_1;
  assign t0_r11_c1_rr5 = a_11_5 * b_5_1;
  assign t0_r11_c1_rr6 = a_11_6 * b_6_1;
  assign t0_r11_c1_rr7 = a_11_7 * b_7_1;
  assign t0_r11_c1_rr8 = a_11_8 * b_8_1;
  assign t0_r11_c1_rr9 = a_11_9 * b_9_1;
  assign t0_r11_c1_rr10 = a_11_10 * b_10_1;
  assign t0_r11_c1_rr11 = a_11_11 * b_11_1;
  assign t0_r11_c1_rr12 = a_11_12 * b_12_1;
  assign t0_r11_c1_rr13 = a_11_13 * b_13_1;
  assign t0_r11_c1_rr14 = a_11_14 * b_14_1;
  assign t1_r11_c1_rr0 = t0_r11_c1_rr0 + t0_r11_c1_rr1;
  assign t1_r11_c1_rr1 = t0_r11_c1_rr2 + t0_r11_c1_rr3;
  assign t1_r11_c1_rr2 = t0_r11_c1_rr4 + t0_r11_c1_rr5;
  assign t1_r11_c1_rr3 = t0_r11_c1_rr6 + t0_r11_c1_rr7;
  assign t1_r11_c1_rr4 = t0_r11_c1_rr8 + t0_r11_c1_rr9;
  assign t1_r11_c1_rr5 = t0_r11_c1_rr10 + t0_r11_c1_rr11;
  assign t1_r11_c1_rr6 = t0_r11_c1_rr12 + t0_r11_c1_rr13;
  assign t1_r11_c1_rr7 = t0_r11_c1_rr14;

  assign t2_r11_c1_rr0 = t1_r11_c1_rr0 + t1_r11_c1_rr1;
  assign t2_r11_c1_rr1 = t1_r11_c1_rr2 + t1_r11_c1_rr3;
  assign t2_r11_c1_rr2 = t1_r11_c1_rr4 + t1_r11_c1_rr5;
  assign t2_r11_c1_rr3 = t1_r11_c1_rr6 + t1_r11_c1_rr7;

  assign t3_r11_c1_rr0 = t2_r11_c1_rr0 + t2_r11_c1_rr1;
  assign t3_r11_c1_rr1 = t2_r11_c1_rr2 + t2_r11_c1_rr3;

  assign t4_r11_c1_rr0 = t3_r11_c1_rr0 + t3_r11_c1_rr1;

  assign c_11_1 = t4_r11_c1_rr0;
  assign t0_r11_c2_rr0 = a_11_0 * b_0_2;
  assign t0_r11_c2_rr1 = a_11_1 * b_1_2;
  assign t0_r11_c2_rr2 = a_11_2 * b_2_2;
  assign t0_r11_c2_rr3 = a_11_3 * b_3_2;
  assign t0_r11_c2_rr4 = a_11_4 * b_4_2;
  assign t0_r11_c2_rr5 = a_11_5 * b_5_2;
  assign t0_r11_c2_rr6 = a_11_6 * b_6_2;
  assign t0_r11_c2_rr7 = a_11_7 * b_7_2;
  assign t0_r11_c2_rr8 = a_11_8 * b_8_2;
  assign t0_r11_c2_rr9 = a_11_9 * b_9_2;
  assign t0_r11_c2_rr10 = a_11_10 * b_10_2;
  assign t0_r11_c2_rr11 = a_11_11 * b_11_2;
  assign t0_r11_c2_rr12 = a_11_12 * b_12_2;
  assign t0_r11_c2_rr13 = a_11_13 * b_13_2;
  assign t0_r11_c2_rr14 = a_11_14 * b_14_2;
  assign t1_r11_c2_rr0 = t0_r11_c2_rr0 + t0_r11_c2_rr1;
  assign t1_r11_c2_rr1 = t0_r11_c2_rr2 + t0_r11_c2_rr3;
  assign t1_r11_c2_rr2 = t0_r11_c2_rr4 + t0_r11_c2_rr5;
  assign t1_r11_c2_rr3 = t0_r11_c2_rr6 + t0_r11_c2_rr7;
  assign t1_r11_c2_rr4 = t0_r11_c2_rr8 + t0_r11_c2_rr9;
  assign t1_r11_c2_rr5 = t0_r11_c2_rr10 + t0_r11_c2_rr11;
  assign t1_r11_c2_rr6 = t0_r11_c2_rr12 + t0_r11_c2_rr13;
  assign t1_r11_c2_rr7 = t0_r11_c2_rr14;

  assign t2_r11_c2_rr0 = t1_r11_c2_rr0 + t1_r11_c2_rr1;
  assign t2_r11_c2_rr1 = t1_r11_c2_rr2 + t1_r11_c2_rr3;
  assign t2_r11_c2_rr2 = t1_r11_c2_rr4 + t1_r11_c2_rr5;
  assign t2_r11_c2_rr3 = t1_r11_c2_rr6 + t1_r11_c2_rr7;

  assign t3_r11_c2_rr0 = t2_r11_c2_rr0 + t2_r11_c2_rr1;
  assign t3_r11_c2_rr1 = t2_r11_c2_rr2 + t2_r11_c2_rr3;

  assign t4_r11_c2_rr0 = t3_r11_c2_rr0 + t3_r11_c2_rr1;

  assign c_11_2 = t4_r11_c2_rr0;
  assign t0_r11_c3_rr0 = a_11_0 * b_0_3;
  assign t0_r11_c3_rr1 = a_11_1 * b_1_3;
  assign t0_r11_c3_rr2 = a_11_2 * b_2_3;
  assign t0_r11_c3_rr3 = a_11_3 * b_3_3;
  assign t0_r11_c3_rr4 = a_11_4 * b_4_3;
  assign t0_r11_c3_rr5 = a_11_5 * b_5_3;
  assign t0_r11_c3_rr6 = a_11_6 * b_6_3;
  assign t0_r11_c3_rr7 = a_11_7 * b_7_3;
  assign t0_r11_c3_rr8 = a_11_8 * b_8_3;
  assign t0_r11_c3_rr9 = a_11_9 * b_9_3;
  assign t0_r11_c3_rr10 = a_11_10 * b_10_3;
  assign t0_r11_c3_rr11 = a_11_11 * b_11_3;
  assign t0_r11_c3_rr12 = a_11_12 * b_12_3;
  assign t0_r11_c3_rr13 = a_11_13 * b_13_3;
  assign t0_r11_c3_rr14 = a_11_14 * b_14_3;
  assign t1_r11_c3_rr0 = t0_r11_c3_rr0 + t0_r11_c3_rr1;
  assign t1_r11_c3_rr1 = t0_r11_c3_rr2 + t0_r11_c3_rr3;
  assign t1_r11_c3_rr2 = t0_r11_c3_rr4 + t0_r11_c3_rr5;
  assign t1_r11_c3_rr3 = t0_r11_c3_rr6 + t0_r11_c3_rr7;
  assign t1_r11_c3_rr4 = t0_r11_c3_rr8 + t0_r11_c3_rr9;
  assign t1_r11_c3_rr5 = t0_r11_c3_rr10 + t0_r11_c3_rr11;
  assign t1_r11_c3_rr6 = t0_r11_c3_rr12 + t0_r11_c3_rr13;
  assign t1_r11_c3_rr7 = t0_r11_c3_rr14;

  assign t2_r11_c3_rr0 = t1_r11_c3_rr0 + t1_r11_c3_rr1;
  assign t2_r11_c3_rr1 = t1_r11_c3_rr2 + t1_r11_c3_rr3;
  assign t2_r11_c3_rr2 = t1_r11_c3_rr4 + t1_r11_c3_rr5;
  assign t2_r11_c3_rr3 = t1_r11_c3_rr6 + t1_r11_c3_rr7;

  assign t3_r11_c3_rr0 = t2_r11_c3_rr0 + t2_r11_c3_rr1;
  assign t3_r11_c3_rr1 = t2_r11_c3_rr2 + t2_r11_c3_rr3;

  assign t4_r11_c3_rr0 = t3_r11_c3_rr0 + t3_r11_c3_rr1;

  assign c_11_3 = t4_r11_c3_rr0;
  assign t0_r11_c4_rr0 = a_11_0 * b_0_4;
  assign t0_r11_c4_rr1 = a_11_1 * b_1_4;
  assign t0_r11_c4_rr2 = a_11_2 * b_2_4;
  assign t0_r11_c4_rr3 = a_11_3 * b_3_4;
  assign t0_r11_c4_rr4 = a_11_4 * b_4_4;
  assign t0_r11_c4_rr5 = a_11_5 * b_5_4;
  assign t0_r11_c4_rr6 = a_11_6 * b_6_4;
  assign t0_r11_c4_rr7 = a_11_7 * b_7_4;
  assign t0_r11_c4_rr8 = a_11_8 * b_8_4;
  assign t0_r11_c4_rr9 = a_11_9 * b_9_4;
  assign t0_r11_c4_rr10 = a_11_10 * b_10_4;
  assign t0_r11_c4_rr11 = a_11_11 * b_11_4;
  assign t0_r11_c4_rr12 = a_11_12 * b_12_4;
  assign t0_r11_c4_rr13 = a_11_13 * b_13_4;
  assign t0_r11_c4_rr14 = a_11_14 * b_14_4;
  assign t1_r11_c4_rr0 = t0_r11_c4_rr0 + t0_r11_c4_rr1;
  assign t1_r11_c4_rr1 = t0_r11_c4_rr2 + t0_r11_c4_rr3;
  assign t1_r11_c4_rr2 = t0_r11_c4_rr4 + t0_r11_c4_rr5;
  assign t1_r11_c4_rr3 = t0_r11_c4_rr6 + t0_r11_c4_rr7;
  assign t1_r11_c4_rr4 = t0_r11_c4_rr8 + t0_r11_c4_rr9;
  assign t1_r11_c4_rr5 = t0_r11_c4_rr10 + t0_r11_c4_rr11;
  assign t1_r11_c4_rr6 = t0_r11_c4_rr12 + t0_r11_c4_rr13;
  assign t1_r11_c4_rr7 = t0_r11_c4_rr14;

  assign t2_r11_c4_rr0 = t1_r11_c4_rr0 + t1_r11_c4_rr1;
  assign t2_r11_c4_rr1 = t1_r11_c4_rr2 + t1_r11_c4_rr3;
  assign t2_r11_c4_rr2 = t1_r11_c4_rr4 + t1_r11_c4_rr5;
  assign t2_r11_c4_rr3 = t1_r11_c4_rr6 + t1_r11_c4_rr7;

  assign t3_r11_c4_rr0 = t2_r11_c4_rr0 + t2_r11_c4_rr1;
  assign t3_r11_c4_rr1 = t2_r11_c4_rr2 + t2_r11_c4_rr3;

  assign t4_r11_c4_rr0 = t3_r11_c4_rr0 + t3_r11_c4_rr1;

  assign c_11_4 = t4_r11_c4_rr0;
  assign t0_r11_c5_rr0 = a_11_0 * b_0_5;
  assign t0_r11_c5_rr1 = a_11_1 * b_1_5;
  assign t0_r11_c5_rr2 = a_11_2 * b_2_5;
  assign t0_r11_c5_rr3 = a_11_3 * b_3_5;
  assign t0_r11_c5_rr4 = a_11_4 * b_4_5;
  assign t0_r11_c5_rr5 = a_11_5 * b_5_5;
  assign t0_r11_c5_rr6 = a_11_6 * b_6_5;
  assign t0_r11_c5_rr7 = a_11_7 * b_7_5;
  assign t0_r11_c5_rr8 = a_11_8 * b_8_5;
  assign t0_r11_c5_rr9 = a_11_9 * b_9_5;
  assign t0_r11_c5_rr10 = a_11_10 * b_10_5;
  assign t0_r11_c5_rr11 = a_11_11 * b_11_5;
  assign t0_r11_c5_rr12 = a_11_12 * b_12_5;
  assign t0_r11_c5_rr13 = a_11_13 * b_13_5;
  assign t0_r11_c5_rr14 = a_11_14 * b_14_5;
  assign t1_r11_c5_rr0 = t0_r11_c5_rr0 + t0_r11_c5_rr1;
  assign t1_r11_c5_rr1 = t0_r11_c5_rr2 + t0_r11_c5_rr3;
  assign t1_r11_c5_rr2 = t0_r11_c5_rr4 + t0_r11_c5_rr5;
  assign t1_r11_c5_rr3 = t0_r11_c5_rr6 + t0_r11_c5_rr7;
  assign t1_r11_c5_rr4 = t0_r11_c5_rr8 + t0_r11_c5_rr9;
  assign t1_r11_c5_rr5 = t0_r11_c5_rr10 + t0_r11_c5_rr11;
  assign t1_r11_c5_rr6 = t0_r11_c5_rr12 + t0_r11_c5_rr13;
  assign t1_r11_c5_rr7 = t0_r11_c5_rr14;

  assign t2_r11_c5_rr0 = t1_r11_c5_rr0 + t1_r11_c5_rr1;
  assign t2_r11_c5_rr1 = t1_r11_c5_rr2 + t1_r11_c5_rr3;
  assign t2_r11_c5_rr2 = t1_r11_c5_rr4 + t1_r11_c5_rr5;
  assign t2_r11_c5_rr3 = t1_r11_c5_rr6 + t1_r11_c5_rr7;

  assign t3_r11_c5_rr0 = t2_r11_c5_rr0 + t2_r11_c5_rr1;
  assign t3_r11_c5_rr1 = t2_r11_c5_rr2 + t2_r11_c5_rr3;

  assign t4_r11_c5_rr0 = t3_r11_c5_rr0 + t3_r11_c5_rr1;

  assign c_11_5 = t4_r11_c5_rr0;
  assign t0_r11_c6_rr0 = a_11_0 * b_0_6;
  assign t0_r11_c6_rr1 = a_11_1 * b_1_6;
  assign t0_r11_c6_rr2 = a_11_2 * b_2_6;
  assign t0_r11_c6_rr3 = a_11_3 * b_3_6;
  assign t0_r11_c6_rr4 = a_11_4 * b_4_6;
  assign t0_r11_c6_rr5 = a_11_5 * b_5_6;
  assign t0_r11_c6_rr6 = a_11_6 * b_6_6;
  assign t0_r11_c6_rr7 = a_11_7 * b_7_6;
  assign t0_r11_c6_rr8 = a_11_8 * b_8_6;
  assign t0_r11_c6_rr9 = a_11_9 * b_9_6;
  assign t0_r11_c6_rr10 = a_11_10 * b_10_6;
  assign t0_r11_c6_rr11 = a_11_11 * b_11_6;
  assign t0_r11_c6_rr12 = a_11_12 * b_12_6;
  assign t0_r11_c6_rr13 = a_11_13 * b_13_6;
  assign t0_r11_c6_rr14 = a_11_14 * b_14_6;
  assign t1_r11_c6_rr0 = t0_r11_c6_rr0 + t0_r11_c6_rr1;
  assign t1_r11_c6_rr1 = t0_r11_c6_rr2 + t0_r11_c6_rr3;
  assign t1_r11_c6_rr2 = t0_r11_c6_rr4 + t0_r11_c6_rr5;
  assign t1_r11_c6_rr3 = t0_r11_c6_rr6 + t0_r11_c6_rr7;
  assign t1_r11_c6_rr4 = t0_r11_c6_rr8 + t0_r11_c6_rr9;
  assign t1_r11_c6_rr5 = t0_r11_c6_rr10 + t0_r11_c6_rr11;
  assign t1_r11_c6_rr6 = t0_r11_c6_rr12 + t0_r11_c6_rr13;
  assign t1_r11_c6_rr7 = t0_r11_c6_rr14;

  assign t2_r11_c6_rr0 = t1_r11_c6_rr0 + t1_r11_c6_rr1;
  assign t2_r11_c6_rr1 = t1_r11_c6_rr2 + t1_r11_c6_rr3;
  assign t2_r11_c6_rr2 = t1_r11_c6_rr4 + t1_r11_c6_rr5;
  assign t2_r11_c6_rr3 = t1_r11_c6_rr6 + t1_r11_c6_rr7;

  assign t3_r11_c6_rr0 = t2_r11_c6_rr0 + t2_r11_c6_rr1;
  assign t3_r11_c6_rr1 = t2_r11_c6_rr2 + t2_r11_c6_rr3;

  assign t4_r11_c6_rr0 = t3_r11_c6_rr0 + t3_r11_c6_rr1;

  assign c_11_6 = t4_r11_c6_rr0;
  assign t0_r11_c7_rr0 = a_11_0 * b_0_7;
  assign t0_r11_c7_rr1 = a_11_1 * b_1_7;
  assign t0_r11_c7_rr2 = a_11_2 * b_2_7;
  assign t0_r11_c7_rr3 = a_11_3 * b_3_7;
  assign t0_r11_c7_rr4 = a_11_4 * b_4_7;
  assign t0_r11_c7_rr5 = a_11_5 * b_5_7;
  assign t0_r11_c7_rr6 = a_11_6 * b_6_7;
  assign t0_r11_c7_rr7 = a_11_7 * b_7_7;
  assign t0_r11_c7_rr8 = a_11_8 * b_8_7;
  assign t0_r11_c7_rr9 = a_11_9 * b_9_7;
  assign t0_r11_c7_rr10 = a_11_10 * b_10_7;
  assign t0_r11_c7_rr11 = a_11_11 * b_11_7;
  assign t0_r11_c7_rr12 = a_11_12 * b_12_7;
  assign t0_r11_c7_rr13 = a_11_13 * b_13_7;
  assign t0_r11_c7_rr14 = a_11_14 * b_14_7;
  assign t1_r11_c7_rr0 = t0_r11_c7_rr0 + t0_r11_c7_rr1;
  assign t1_r11_c7_rr1 = t0_r11_c7_rr2 + t0_r11_c7_rr3;
  assign t1_r11_c7_rr2 = t0_r11_c7_rr4 + t0_r11_c7_rr5;
  assign t1_r11_c7_rr3 = t0_r11_c7_rr6 + t0_r11_c7_rr7;
  assign t1_r11_c7_rr4 = t0_r11_c7_rr8 + t0_r11_c7_rr9;
  assign t1_r11_c7_rr5 = t0_r11_c7_rr10 + t0_r11_c7_rr11;
  assign t1_r11_c7_rr6 = t0_r11_c7_rr12 + t0_r11_c7_rr13;
  assign t1_r11_c7_rr7 = t0_r11_c7_rr14;

  assign t2_r11_c7_rr0 = t1_r11_c7_rr0 + t1_r11_c7_rr1;
  assign t2_r11_c7_rr1 = t1_r11_c7_rr2 + t1_r11_c7_rr3;
  assign t2_r11_c7_rr2 = t1_r11_c7_rr4 + t1_r11_c7_rr5;
  assign t2_r11_c7_rr3 = t1_r11_c7_rr6 + t1_r11_c7_rr7;

  assign t3_r11_c7_rr0 = t2_r11_c7_rr0 + t2_r11_c7_rr1;
  assign t3_r11_c7_rr1 = t2_r11_c7_rr2 + t2_r11_c7_rr3;

  assign t4_r11_c7_rr0 = t3_r11_c7_rr0 + t3_r11_c7_rr1;

  assign c_11_7 = t4_r11_c7_rr0;
  assign t0_r11_c8_rr0 = a_11_0 * b_0_8;
  assign t0_r11_c8_rr1 = a_11_1 * b_1_8;
  assign t0_r11_c8_rr2 = a_11_2 * b_2_8;
  assign t0_r11_c8_rr3 = a_11_3 * b_3_8;
  assign t0_r11_c8_rr4 = a_11_4 * b_4_8;
  assign t0_r11_c8_rr5 = a_11_5 * b_5_8;
  assign t0_r11_c8_rr6 = a_11_6 * b_6_8;
  assign t0_r11_c8_rr7 = a_11_7 * b_7_8;
  assign t0_r11_c8_rr8 = a_11_8 * b_8_8;
  assign t0_r11_c8_rr9 = a_11_9 * b_9_8;
  assign t0_r11_c8_rr10 = a_11_10 * b_10_8;
  assign t0_r11_c8_rr11 = a_11_11 * b_11_8;
  assign t0_r11_c8_rr12 = a_11_12 * b_12_8;
  assign t0_r11_c8_rr13 = a_11_13 * b_13_8;
  assign t0_r11_c8_rr14 = a_11_14 * b_14_8;
  assign t1_r11_c8_rr0 = t0_r11_c8_rr0 + t0_r11_c8_rr1;
  assign t1_r11_c8_rr1 = t0_r11_c8_rr2 + t0_r11_c8_rr3;
  assign t1_r11_c8_rr2 = t0_r11_c8_rr4 + t0_r11_c8_rr5;
  assign t1_r11_c8_rr3 = t0_r11_c8_rr6 + t0_r11_c8_rr7;
  assign t1_r11_c8_rr4 = t0_r11_c8_rr8 + t0_r11_c8_rr9;
  assign t1_r11_c8_rr5 = t0_r11_c8_rr10 + t0_r11_c8_rr11;
  assign t1_r11_c8_rr6 = t0_r11_c8_rr12 + t0_r11_c8_rr13;
  assign t1_r11_c8_rr7 = t0_r11_c8_rr14;

  assign t2_r11_c8_rr0 = t1_r11_c8_rr0 + t1_r11_c8_rr1;
  assign t2_r11_c8_rr1 = t1_r11_c8_rr2 + t1_r11_c8_rr3;
  assign t2_r11_c8_rr2 = t1_r11_c8_rr4 + t1_r11_c8_rr5;
  assign t2_r11_c8_rr3 = t1_r11_c8_rr6 + t1_r11_c8_rr7;

  assign t3_r11_c8_rr0 = t2_r11_c8_rr0 + t2_r11_c8_rr1;
  assign t3_r11_c8_rr1 = t2_r11_c8_rr2 + t2_r11_c8_rr3;

  assign t4_r11_c8_rr0 = t3_r11_c8_rr0 + t3_r11_c8_rr1;

  assign c_11_8 = t4_r11_c8_rr0;
  assign t0_r11_c9_rr0 = a_11_0 * b_0_9;
  assign t0_r11_c9_rr1 = a_11_1 * b_1_9;
  assign t0_r11_c9_rr2 = a_11_2 * b_2_9;
  assign t0_r11_c9_rr3 = a_11_3 * b_3_9;
  assign t0_r11_c9_rr4 = a_11_4 * b_4_9;
  assign t0_r11_c9_rr5 = a_11_5 * b_5_9;
  assign t0_r11_c9_rr6 = a_11_6 * b_6_9;
  assign t0_r11_c9_rr7 = a_11_7 * b_7_9;
  assign t0_r11_c9_rr8 = a_11_8 * b_8_9;
  assign t0_r11_c9_rr9 = a_11_9 * b_9_9;
  assign t0_r11_c9_rr10 = a_11_10 * b_10_9;
  assign t0_r11_c9_rr11 = a_11_11 * b_11_9;
  assign t0_r11_c9_rr12 = a_11_12 * b_12_9;
  assign t0_r11_c9_rr13 = a_11_13 * b_13_9;
  assign t0_r11_c9_rr14 = a_11_14 * b_14_9;
  assign t1_r11_c9_rr0 = t0_r11_c9_rr0 + t0_r11_c9_rr1;
  assign t1_r11_c9_rr1 = t0_r11_c9_rr2 + t0_r11_c9_rr3;
  assign t1_r11_c9_rr2 = t0_r11_c9_rr4 + t0_r11_c9_rr5;
  assign t1_r11_c9_rr3 = t0_r11_c9_rr6 + t0_r11_c9_rr7;
  assign t1_r11_c9_rr4 = t0_r11_c9_rr8 + t0_r11_c9_rr9;
  assign t1_r11_c9_rr5 = t0_r11_c9_rr10 + t0_r11_c9_rr11;
  assign t1_r11_c9_rr6 = t0_r11_c9_rr12 + t0_r11_c9_rr13;
  assign t1_r11_c9_rr7 = t0_r11_c9_rr14;

  assign t2_r11_c9_rr0 = t1_r11_c9_rr0 + t1_r11_c9_rr1;
  assign t2_r11_c9_rr1 = t1_r11_c9_rr2 + t1_r11_c9_rr3;
  assign t2_r11_c9_rr2 = t1_r11_c9_rr4 + t1_r11_c9_rr5;
  assign t2_r11_c9_rr3 = t1_r11_c9_rr6 + t1_r11_c9_rr7;

  assign t3_r11_c9_rr0 = t2_r11_c9_rr0 + t2_r11_c9_rr1;
  assign t3_r11_c9_rr1 = t2_r11_c9_rr2 + t2_r11_c9_rr3;

  assign t4_r11_c9_rr0 = t3_r11_c9_rr0 + t3_r11_c9_rr1;

  assign c_11_9 = t4_r11_c9_rr0;
  assign t0_r11_c10_rr0 = a_11_0 * b_0_10;
  assign t0_r11_c10_rr1 = a_11_1 * b_1_10;
  assign t0_r11_c10_rr2 = a_11_2 * b_2_10;
  assign t0_r11_c10_rr3 = a_11_3 * b_3_10;
  assign t0_r11_c10_rr4 = a_11_4 * b_4_10;
  assign t0_r11_c10_rr5 = a_11_5 * b_5_10;
  assign t0_r11_c10_rr6 = a_11_6 * b_6_10;
  assign t0_r11_c10_rr7 = a_11_7 * b_7_10;
  assign t0_r11_c10_rr8 = a_11_8 * b_8_10;
  assign t0_r11_c10_rr9 = a_11_9 * b_9_10;
  assign t0_r11_c10_rr10 = a_11_10 * b_10_10;
  assign t0_r11_c10_rr11 = a_11_11 * b_11_10;
  assign t0_r11_c10_rr12 = a_11_12 * b_12_10;
  assign t0_r11_c10_rr13 = a_11_13 * b_13_10;
  assign t0_r11_c10_rr14 = a_11_14 * b_14_10;
  assign t1_r11_c10_rr0 = t0_r11_c10_rr0 + t0_r11_c10_rr1;
  assign t1_r11_c10_rr1 = t0_r11_c10_rr2 + t0_r11_c10_rr3;
  assign t1_r11_c10_rr2 = t0_r11_c10_rr4 + t0_r11_c10_rr5;
  assign t1_r11_c10_rr3 = t0_r11_c10_rr6 + t0_r11_c10_rr7;
  assign t1_r11_c10_rr4 = t0_r11_c10_rr8 + t0_r11_c10_rr9;
  assign t1_r11_c10_rr5 = t0_r11_c10_rr10 + t0_r11_c10_rr11;
  assign t1_r11_c10_rr6 = t0_r11_c10_rr12 + t0_r11_c10_rr13;
  assign t1_r11_c10_rr7 = t0_r11_c10_rr14;

  assign t2_r11_c10_rr0 = t1_r11_c10_rr0 + t1_r11_c10_rr1;
  assign t2_r11_c10_rr1 = t1_r11_c10_rr2 + t1_r11_c10_rr3;
  assign t2_r11_c10_rr2 = t1_r11_c10_rr4 + t1_r11_c10_rr5;
  assign t2_r11_c10_rr3 = t1_r11_c10_rr6 + t1_r11_c10_rr7;

  assign t3_r11_c10_rr0 = t2_r11_c10_rr0 + t2_r11_c10_rr1;
  assign t3_r11_c10_rr1 = t2_r11_c10_rr2 + t2_r11_c10_rr3;

  assign t4_r11_c10_rr0 = t3_r11_c10_rr0 + t3_r11_c10_rr1;

  assign c_11_10 = t4_r11_c10_rr0;
  assign t0_r11_c11_rr0 = a_11_0 * b_0_11;
  assign t0_r11_c11_rr1 = a_11_1 * b_1_11;
  assign t0_r11_c11_rr2 = a_11_2 * b_2_11;
  assign t0_r11_c11_rr3 = a_11_3 * b_3_11;
  assign t0_r11_c11_rr4 = a_11_4 * b_4_11;
  assign t0_r11_c11_rr5 = a_11_5 * b_5_11;
  assign t0_r11_c11_rr6 = a_11_6 * b_6_11;
  assign t0_r11_c11_rr7 = a_11_7 * b_7_11;
  assign t0_r11_c11_rr8 = a_11_8 * b_8_11;
  assign t0_r11_c11_rr9 = a_11_9 * b_9_11;
  assign t0_r11_c11_rr10 = a_11_10 * b_10_11;
  assign t0_r11_c11_rr11 = a_11_11 * b_11_11;
  assign t0_r11_c11_rr12 = a_11_12 * b_12_11;
  assign t0_r11_c11_rr13 = a_11_13 * b_13_11;
  assign t0_r11_c11_rr14 = a_11_14 * b_14_11;
  assign t1_r11_c11_rr0 = t0_r11_c11_rr0 + t0_r11_c11_rr1;
  assign t1_r11_c11_rr1 = t0_r11_c11_rr2 + t0_r11_c11_rr3;
  assign t1_r11_c11_rr2 = t0_r11_c11_rr4 + t0_r11_c11_rr5;
  assign t1_r11_c11_rr3 = t0_r11_c11_rr6 + t0_r11_c11_rr7;
  assign t1_r11_c11_rr4 = t0_r11_c11_rr8 + t0_r11_c11_rr9;
  assign t1_r11_c11_rr5 = t0_r11_c11_rr10 + t0_r11_c11_rr11;
  assign t1_r11_c11_rr6 = t0_r11_c11_rr12 + t0_r11_c11_rr13;
  assign t1_r11_c11_rr7 = t0_r11_c11_rr14;

  assign t2_r11_c11_rr0 = t1_r11_c11_rr0 + t1_r11_c11_rr1;
  assign t2_r11_c11_rr1 = t1_r11_c11_rr2 + t1_r11_c11_rr3;
  assign t2_r11_c11_rr2 = t1_r11_c11_rr4 + t1_r11_c11_rr5;
  assign t2_r11_c11_rr3 = t1_r11_c11_rr6 + t1_r11_c11_rr7;

  assign t3_r11_c11_rr0 = t2_r11_c11_rr0 + t2_r11_c11_rr1;
  assign t3_r11_c11_rr1 = t2_r11_c11_rr2 + t2_r11_c11_rr3;

  assign t4_r11_c11_rr0 = t3_r11_c11_rr0 + t3_r11_c11_rr1;

  assign c_11_11 = t4_r11_c11_rr0;
  assign t0_r11_c12_rr0 = a_11_0 * b_0_12;
  assign t0_r11_c12_rr1 = a_11_1 * b_1_12;
  assign t0_r11_c12_rr2 = a_11_2 * b_2_12;
  assign t0_r11_c12_rr3 = a_11_3 * b_3_12;
  assign t0_r11_c12_rr4 = a_11_4 * b_4_12;
  assign t0_r11_c12_rr5 = a_11_5 * b_5_12;
  assign t0_r11_c12_rr6 = a_11_6 * b_6_12;
  assign t0_r11_c12_rr7 = a_11_7 * b_7_12;
  assign t0_r11_c12_rr8 = a_11_8 * b_8_12;
  assign t0_r11_c12_rr9 = a_11_9 * b_9_12;
  assign t0_r11_c12_rr10 = a_11_10 * b_10_12;
  assign t0_r11_c12_rr11 = a_11_11 * b_11_12;
  assign t0_r11_c12_rr12 = a_11_12 * b_12_12;
  assign t0_r11_c12_rr13 = a_11_13 * b_13_12;
  assign t0_r11_c12_rr14 = a_11_14 * b_14_12;
  assign t1_r11_c12_rr0 = t0_r11_c12_rr0 + t0_r11_c12_rr1;
  assign t1_r11_c12_rr1 = t0_r11_c12_rr2 + t0_r11_c12_rr3;
  assign t1_r11_c12_rr2 = t0_r11_c12_rr4 + t0_r11_c12_rr5;
  assign t1_r11_c12_rr3 = t0_r11_c12_rr6 + t0_r11_c12_rr7;
  assign t1_r11_c12_rr4 = t0_r11_c12_rr8 + t0_r11_c12_rr9;
  assign t1_r11_c12_rr5 = t0_r11_c12_rr10 + t0_r11_c12_rr11;
  assign t1_r11_c12_rr6 = t0_r11_c12_rr12 + t0_r11_c12_rr13;
  assign t1_r11_c12_rr7 = t0_r11_c12_rr14;

  assign t2_r11_c12_rr0 = t1_r11_c12_rr0 + t1_r11_c12_rr1;
  assign t2_r11_c12_rr1 = t1_r11_c12_rr2 + t1_r11_c12_rr3;
  assign t2_r11_c12_rr2 = t1_r11_c12_rr4 + t1_r11_c12_rr5;
  assign t2_r11_c12_rr3 = t1_r11_c12_rr6 + t1_r11_c12_rr7;

  assign t3_r11_c12_rr0 = t2_r11_c12_rr0 + t2_r11_c12_rr1;
  assign t3_r11_c12_rr1 = t2_r11_c12_rr2 + t2_r11_c12_rr3;

  assign t4_r11_c12_rr0 = t3_r11_c12_rr0 + t3_r11_c12_rr1;

  assign c_11_12 = t4_r11_c12_rr0;
  assign t0_r11_c13_rr0 = a_11_0 * b_0_13;
  assign t0_r11_c13_rr1 = a_11_1 * b_1_13;
  assign t0_r11_c13_rr2 = a_11_2 * b_2_13;
  assign t0_r11_c13_rr3 = a_11_3 * b_3_13;
  assign t0_r11_c13_rr4 = a_11_4 * b_4_13;
  assign t0_r11_c13_rr5 = a_11_5 * b_5_13;
  assign t0_r11_c13_rr6 = a_11_6 * b_6_13;
  assign t0_r11_c13_rr7 = a_11_7 * b_7_13;
  assign t0_r11_c13_rr8 = a_11_8 * b_8_13;
  assign t0_r11_c13_rr9 = a_11_9 * b_9_13;
  assign t0_r11_c13_rr10 = a_11_10 * b_10_13;
  assign t0_r11_c13_rr11 = a_11_11 * b_11_13;
  assign t0_r11_c13_rr12 = a_11_12 * b_12_13;
  assign t0_r11_c13_rr13 = a_11_13 * b_13_13;
  assign t0_r11_c13_rr14 = a_11_14 * b_14_13;
  assign t1_r11_c13_rr0 = t0_r11_c13_rr0 + t0_r11_c13_rr1;
  assign t1_r11_c13_rr1 = t0_r11_c13_rr2 + t0_r11_c13_rr3;
  assign t1_r11_c13_rr2 = t0_r11_c13_rr4 + t0_r11_c13_rr5;
  assign t1_r11_c13_rr3 = t0_r11_c13_rr6 + t0_r11_c13_rr7;
  assign t1_r11_c13_rr4 = t0_r11_c13_rr8 + t0_r11_c13_rr9;
  assign t1_r11_c13_rr5 = t0_r11_c13_rr10 + t0_r11_c13_rr11;
  assign t1_r11_c13_rr6 = t0_r11_c13_rr12 + t0_r11_c13_rr13;
  assign t1_r11_c13_rr7 = t0_r11_c13_rr14;

  assign t2_r11_c13_rr0 = t1_r11_c13_rr0 + t1_r11_c13_rr1;
  assign t2_r11_c13_rr1 = t1_r11_c13_rr2 + t1_r11_c13_rr3;
  assign t2_r11_c13_rr2 = t1_r11_c13_rr4 + t1_r11_c13_rr5;
  assign t2_r11_c13_rr3 = t1_r11_c13_rr6 + t1_r11_c13_rr7;

  assign t3_r11_c13_rr0 = t2_r11_c13_rr0 + t2_r11_c13_rr1;
  assign t3_r11_c13_rr1 = t2_r11_c13_rr2 + t2_r11_c13_rr3;

  assign t4_r11_c13_rr0 = t3_r11_c13_rr0 + t3_r11_c13_rr1;

  assign c_11_13 = t4_r11_c13_rr0;
  assign t0_r11_c14_rr0 = a_11_0 * b_0_14;
  assign t0_r11_c14_rr1 = a_11_1 * b_1_14;
  assign t0_r11_c14_rr2 = a_11_2 * b_2_14;
  assign t0_r11_c14_rr3 = a_11_3 * b_3_14;
  assign t0_r11_c14_rr4 = a_11_4 * b_4_14;
  assign t0_r11_c14_rr5 = a_11_5 * b_5_14;
  assign t0_r11_c14_rr6 = a_11_6 * b_6_14;
  assign t0_r11_c14_rr7 = a_11_7 * b_7_14;
  assign t0_r11_c14_rr8 = a_11_8 * b_8_14;
  assign t0_r11_c14_rr9 = a_11_9 * b_9_14;
  assign t0_r11_c14_rr10 = a_11_10 * b_10_14;
  assign t0_r11_c14_rr11 = a_11_11 * b_11_14;
  assign t0_r11_c14_rr12 = a_11_12 * b_12_14;
  assign t0_r11_c14_rr13 = a_11_13 * b_13_14;
  assign t0_r11_c14_rr14 = a_11_14 * b_14_14;
  assign t1_r11_c14_rr0 = t0_r11_c14_rr0 + t0_r11_c14_rr1;
  assign t1_r11_c14_rr1 = t0_r11_c14_rr2 + t0_r11_c14_rr3;
  assign t1_r11_c14_rr2 = t0_r11_c14_rr4 + t0_r11_c14_rr5;
  assign t1_r11_c14_rr3 = t0_r11_c14_rr6 + t0_r11_c14_rr7;
  assign t1_r11_c14_rr4 = t0_r11_c14_rr8 + t0_r11_c14_rr9;
  assign t1_r11_c14_rr5 = t0_r11_c14_rr10 + t0_r11_c14_rr11;
  assign t1_r11_c14_rr6 = t0_r11_c14_rr12 + t0_r11_c14_rr13;
  assign t1_r11_c14_rr7 = t0_r11_c14_rr14;

  assign t2_r11_c14_rr0 = t1_r11_c14_rr0 + t1_r11_c14_rr1;
  assign t2_r11_c14_rr1 = t1_r11_c14_rr2 + t1_r11_c14_rr3;
  assign t2_r11_c14_rr2 = t1_r11_c14_rr4 + t1_r11_c14_rr5;
  assign t2_r11_c14_rr3 = t1_r11_c14_rr6 + t1_r11_c14_rr7;

  assign t3_r11_c14_rr0 = t2_r11_c14_rr0 + t2_r11_c14_rr1;
  assign t3_r11_c14_rr1 = t2_r11_c14_rr2 + t2_r11_c14_rr3;

  assign t4_r11_c14_rr0 = t3_r11_c14_rr0 + t3_r11_c14_rr1;

  assign c_11_14 = t4_r11_c14_rr0;
  assign t0_r12_c0_rr0 = a_12_0 * b_0_0;
  assign t0_r12_c0_rr1 = a_12_1 * b_1_0;
  assign t0_r12_c0_rr2 = a_12_2 * b_2_0;
  assign t0_r12_c0_rr3 = a_12_3 * b_3_0;
  assign t0_r12_c0_rr4 = a_12_4 * b_4_0;
  assign t0_r12_c0_rr5 = a_12_5 * b_5_0;
  assign t0_r12_c0_rr6 = a_12_6 * b_6_0;
  assign t0_r12_c0_rr7 = a_12_7 * b_7_0;
  assign t0_r12_c0_rr8 = a_12_8 * b_8_0;
  assign t0_r12_c0_rr9 = a_12_9 * b_9_0;
  assign t0_r12_c0_rr10 = a_12_10 * b_10_0;
  assign t0_r12_c0_rr11 = a_12_11 * b_11_0;
  assign t0_r12_c0_rr12 = a_12_12 * b_12_0;
  assign t0_r12_c0_rr13 = a_12_13 * b_13_0;
  assign t0_r12_c0_rr14 = a_12_14 * b_14_0;
  assign t1_r12_c0_rr0 = t0_r12_c0_rr0 + t0_r12_c0_rr1;
  assign t1_r12_c0_rr1 = t0_r12_c0_rr2 + t0_r12_c0_rr3;
  assign t1_r12_c0_rr2 = t0_r12_c0_rr4 + t0_r12_c0_rr5;
  assign t1_r12_c0_rr3 = t0_r12_c0_rr6 + t0_r12_c0_rr7;
  assign t1_r12_c0_rr4 = t0_r12_c0_rr8 + t0_r12_c0_rr9;
  assign t1_r12_c0_rr5 = t0_r12_c0_rr10 + t0_r12_c0_rr11;
  assign t1_r12_c0_rr6 = t0_r12_c0_rr12 + t0_r12_c0_rr13;
  assign t1_r12_c0_rr7 = t0_r12_c0_rr14;

  assign t2_r12_c0_rr0 = t1_r12_c0_rr0 + t1_r12_c0_rr1;
  assign t2_r12_c0_rr1 = t1_r12_c0_rr2 + t1_r12_c0_rr3;
  assign t2_r12_c0_rr2 = t1_r12_c0_rr4 + t1_r12_c0_rr5;
  assign t2_r12_c0_rr3 = t1_r12_c0_rr6 + t1_r12_c0_rr7;

  assign t3_r12_c0_rr0 = t2_r12_c0_rr0 + t2_r12_c0_rr1;
  assign t3_r12_c0_rr1 = t2_r12_c0_rr2 + t2_r12_c0_rr3;

  assign t4_r12_c0_rr0 = t3_r12_c0_rr0 + t3_r12_c0_rr1;

  assign c_12_0 = t4_r12_c0_rr0;
  assign t0_r12_c1_rr0 = a_12_0 * b_0_1;
  assign t0_r12_c1_rr1 = a_12_1 * b_1_1;
  assign t0_r12_c1_rr2 = a_12_2 * b_2_1;
  assign t0_r12_c1_rr3 = a_12_3 * b_3_1;
  assign t0_r12_c1_rr4 = a_12_4 * b_4_1;
  assign t0_r12_c1_rr5 = a_12_5 * b_5_1;
  assign t0_r12_c1_rr6 = a_12_6 * b_6_1;
  assign t0_r12_c1_rr7 = a_12_7 * b_7_1;
  assign t0_r12_c1_rr8 = a_12_8 * b_8_1;
  assign t0_r12_c1_rr9 = a_12_9 * b_9_1;
  assign t0_r12_c1_rr10 = a_12_10 * b_10_1;
  assign t0_r12_c1_rr11 = a_12_11 * b_11_1;
  assign t0_r12_c1_rr12 = a_12_12 * b_12_1;
  assign t0_r12_c1_rr13 = a_12_13 * b_13_1;
  assign t0_r12_c1_rr14 = a_12_14 * b_14_1;
  assign t1_r12_c1_rr0 = t0_r12_c1_rr0 + t0_r12_c1_rr1;
  assign t1_r12_c1_rr1 = t0_r12_c1_rr2 + t0_r12_c1_rr3;
  assign t1_r12_c1_rr2 = t0_r12_c1_rr4 + t0_r12_c1_rr5;
  assign t1_r12_c1_rr3 = t0_r12_c1_rr6 + t0_r12_c1_rr7;
  assign t1_r12_c1_rr4 = t0_r12_c1_rr8 + t0_r12_c1_rr9;
  assign t1_r12_c1_rr5 = t0_r12_c1_rr10 + t0_r12_c1_rr11;
  assign t1_r12_c1_rr6 = t0_r12_c1_rr12 + t0_r12_c1_rr13;
  assign t1_r12_c1_rr7 = t0_r12_c1_rr14;

  assign t2_r12_c1_rr0 = t1_r12_c1_rr0 + t1_r12_c1_rr1;
  assign t2_r12_c1_rr1 = t1_r12_c1_rr2 + t1_r12_c1_rr3;
  assign t2_r12_c1_rr2 = t1_r12_c1_rr4 + t1_r12_c1_rr5;
  assign t2_r12_c1_rr3 = t1_r12_c1_rr6 + t1_r12_c1_rr7;

  assign t3_r12_c1_rr0 = t2_r12_c1_rr0 + t2_r12_c1_rr1;
  assign t3_r12_c1_rr1 = t2_r12_c1_rr2 + t2_r12_c1_rr3;

  assign t4_r12_c1_rr0 = t3_r12_c1_rr0 + t3_r12_c1_rr1;

  assign c_12_1 = t4_r12_c1_rr0;
  assign t0_r12_c2_rr0 = a_12_0 * b_0_2;
  assign t0_r12_c2_rr1 = a_12_1 * b_1_2;
  assign t0_r12_c2_rr2 = a_12_2 * b_2_2;
  assign t0_r12_c2_rr3 = a_12_3 * b_3_2;
  assign t0_r12_c2_rr4 = a_12_4 * b_4_2;
  assign t0_r12_c2_rr5 = a_12_5 * b_5_2;
  assign t0_r12_c2_rr6 = a_12_6 * b_6_2;
  assign t0_r12_c2_rr7 = a_12_7 * b_7_2;
  assign t0_r12_c2_rr8 = a_12_8 * b_8_2;
  assign t0_r12_c2_rr9 = a_12_9 * b_9_2;
  assign t0_r12_c2_rr10 = a_12_10 * b_10_2;
  assign t0_r12_c2_rr11 = a_12_11 * b_11_2;
  assign t0_r12_c2_rr12 = a_12_12 * b_12_2;
  assign t0_r12_c2_rr13 = a_12_13 * b_13_2;
  assign t0_r12_c2_rr14 = a_12_14 * b_14_2;
  assign t1_r12_c2_rr0 = t0_r12_c2_rr0 + t0_r12_c2_rr1;
  assign t1_r12_c2_rr1 = t0_r12_c2_rr2 + t0_r12_c2_rr3;
  assign t1_r12_c2_rr2 = t0_r12_c2_rr4 + t0_r12_c2_rr5;
  assign t1_r12_c2_rr3 = t0_r12_c2_rr6 + t0_r12_c2_rr7;
  assign t1_r12_c2_rr4 = t0_r12_c2_rr8 + t0_r12_c2_rr9;
  assign t1_r12_c2_rr5 = t0_r12_c2_rr10 + t0_r12_c2_rr11;
  assign t1_r12_c2_rr6 = t0_r12_c2_rr12 + t0_r12_c2_rr13;
  assign t1_r12_c2_rr7 = t0_r12_c2_rr14;

  assign t2_r12_c2_rr0 = t1_r12_c2_rr0 + t1_r12_c2_rr1;
  assign t2_r12_c2_rr1 = t1_r12_c2_rr2 + t1_r12_c2_rr3;
  assign t2_r12_c2_rr2 = t1_r12_c2_rr4 + t1_r12_c2_rr5;
  assign t2_r12_c2_rr3 = t1_r12_c2_rr6 + t1_r12_c2_rr7;

  assign t3_r12_c2_rr0 = t2_r12_c2_rr0 + t2_r12_c2_rr1;
  assign t3_r12_c2_rr1 = t2_r12_c2_rr2 + t2_r12_c2_rr3;

  assign t4_r12_c2_rr0 = t3_r12_c2_rr0 + t3_r12_c2_rr1;

  assign c_12_2 = t4_r12_c2_rr0;
  assign t0_r12_c3_rr0 = a_12_0 * b_0_3;
  assign t0_r12_c3_rr1 = a_12_1 * b_1_3;
  assign t0_r12_c3_rr2 = a_12_2 * b_2_3;
  assign t0_r12_c3_rr3 = a_12_3 * b_3_3;
  assign t0_r12_c3_rr4 = a_12_4 * b_4_3;
  assign t0_r12_c3_rr5 = a_12_5 * b_5_3;
  assign t0_r12_c3_rr6 = a_12_6 * b_6_3;
  assign t0_r12_c3_rr7 = a_12_7 * b_7_3;
  assign t0_r12_c3_rr8 = a_12_8 * b_8_3;
  assign t0_r12_c3_rr9 = a_12_9 * b_9_3;
  assign t0_r12_c3_rr10 = a_12_10 * b_10_3;
  assign t0_r12_c3_rr11 = a_12_11 * b_11_3;
  assign t0_r12_c3_rr12 = a_12_12 * b_12_3;
  assign t0_r12_c3_rr13 = a_12_13 * b_13_3;
  assign t0_r12_c3_rr14 = a_12_14 * b_14_3;
  assign t1_r12_c3_rr0 = t0_r12_c3_rr0 + t0_r12_c3_rr1;
  assign t1_r12_c3_rr1 = t0_r12_c3_rr2 + t0_r12_c3_rr3;
  assign t1_r12_c3_rr2 = t0_r12_c3_rr4 + t0_r12_c3_rr5;
  assign t1_r12_c3_rr3 = t0_r12_c3_rr6 + t0_r12_c3_rr7;
  assign t1_r12_c3_rr4 = t0_r12_c3_rr8 + t0_r12_c3_rr9;
  assign t1_r12_c3_rr5 = t0_r12_c3_rr10 + t0_r12_c3_rr11;
  assign t1_r12_c3_rr6 = t0_r12_c3_rr12 + t0_r12_c3_rr13;
  assign t1_r12_c3_rr7 = t0_r12_c3_rr14;

  assign t2_r12_c3_rr0 = t1_r12_c3_rr0 + t1_r12_c3_rr1;
  assign t2_r12_c3_rr1 = t1_r12_c3_rr2 + t1_r12_c3_rr3;
  assign t2_r12_c3_rr2 = t1_r12_c3_rr4 + t1_r12_c3_rr5;
  assign t2_r12_c3_rr3 = t1_r12_c3_rr6 + t1_r12_c3_rr7;

  assign t3_r12_c3_rr0 = t2_r12_c3_rr0 + t2_r12_c3_rr1;
  assign t3_r12_c3_rr1 = t2_r12_c3_rr2 + t2_r12_c3_rr3;

  assign t4_r12_c3_rr0 = t3_r12_c3_rr0 + t3_r12_c3_rr1;

  assign c_12_3 = t4_r12_c3_rr0;
  assign t0_r12_c4_rr0 = a_12_0 * b_0_4;
  assign t0_r12_c4_rr1 = a_12_1 * b_1_4;
  assign t0_r12_c4_rr2 = a_12_2 * b_2_4;
  assign t0_r12_c4_rr3 = a_12_3 * b_3_4;
  assign t0_r12_c4_rr4 = a_12_4 * b_4_4;
  assign t0_r12_c4_rr5 = a_12_5 * b_5_4;
  assign t0_r12_c4_rr6 = a_12_6 * b_6_4;
  assign t0_r12_c4_rr7 = a_12_7 * b_7_4;
  assign t0_r12_c4_rr8 = a_12_8 * b_8_4;
  assign t0_r12_c4_rr9 = a_12_9 * b_9_4;
  assign t0_r12_c4_rr10 = a_12_10 * b_10_4;
  assign t0_r12_c4_rr11 = a_12_11 * b_11_4;
  assign t0_r12_c4_rr12 = a_12_12 * b_12_4;
  assign t0_r12_c4_rr13 = a_12_13 * b_13_4;
  assign t0_r12_c4_rr14 = a_12_14 * b_14_4;
  assign t1_r12_c4_rr0 = t0_r12_c4_rr0 + t0_r12_c4_rr1;
  assign t1_r12_c4_rr1 = t0_r12_c4_rr2 + t0_r12_c4_rr3;
  assign t1_r12_c4_rr2 = t0_r12_c4_rr4 + t0_r12_c4_rr5;
  assign t1_r12_c4_rr3 = t0_r12_c4_rr6 + t0_r12_c4_rr7;
  assign t1_r12_c4_rr4 = t0_r12_c4_rr8 + t0_r12_c4_rr9;
  assign t1_r12_c4_rr5 = t0_r12_c4_rr10 + t0_r12_c4_rr11;
  assign t1_r12_c4_rr6 = t0_r12_c4_rr12 + t0_r12_c4_rr13;
  assign t1_r12_c4_rr7 = t0_r12_c4_rr14;

  assign t2_r12_c4_rr0 = t1_r12_c4_rr0 + t1_r12_c4_rr1;
  assign t2_r12_c4_rr1 = t1_r12_c4_rr2 + t1_r12_c4_rr3;
  assign t2_r12_c4_rr2 = t1_r12_c4_rr4 + t1_r12_c4_rr5;
  assign t2_r12_c4_rr3 = t1_r12_c4_rr6 + t1_r12_c4_rr7;

  assign t3_r12_c4_rr0 = t2_r12_c4_rr0 + t2_r12_c4_rr1;
  assign t3_r12_c4_rr1 = t2_r12_c4_rr2 + t2_r12_c4_rr3;

  assign t4_r12_c4_rr0 = t3_r12_c4_rr0 + t3_r12_c4_rr1;

  assign c_12_4 = t4_r12_c4_rr0;
  assign t0_r12_c5_rr0 = a_12_0 * b_0_5;
  assign t0_r12_c5_rr1 = a_12_1 * b_1_5;
  assign t0_r12_c5_rr2 = a_12_2 * b_2_5;
  assign t0_r12_c5_rr3 = a_12_3 * b_3_5;
  assign t0_r12_c5_rr4 = a_12_4 * b_4_5;
  assign t0_r12_c5_rr5 = a_12_5 * b_5_5;
  assign t0_r12_c5_rr6 = a_12_6 * b_6_5;
  assign t0_r12_c5_rr7 = a_12_7 * b_7_5;
  assign t0_r12_c5_rr8 = a_12_8 * b_8_5;
  assign t0_r12_c5_rr9 = a_12_9 * b_9_5;
  assign t0_r12_c5_rr10 = a_12_10 * b_10_5;
  assign t0_r12_c5_rr11 = a_12_11 * b_11_5;
  assign t0_r12_c5_rr12 = a_12_12 * b_12_5;
  assign t0_r12_c5_rr13 = a_12_13 * b_13_5;
  assign t0_r12_c5_rr14 = a_12_14 * b_14_5;
  assign t1_r12_c5_rr0 = t0_r12_c5_rr0 + t0_r12_c5_rr1;
  assign t1_r12_c5_rr1 = t0_r12_c5_rr2 + t0_r12_c5_rr3;
  assign t1_r12_c5_rr2 = t0_r12_c5_rr4 + t0_r12_c5_rr5;
  assign t1_r12_c5_rr3 = t0_r12_c5_rr6 + t0_r12_c5_rr7;
  assign t1_r12_c5_rr4 = t0_r12_c5_rr8 + t0_r12_c5_rr9;
  assign t1_r12_c5_rr5 = t0_r12_c5_rr10 + t0_r12_c5_rr11;
  assign t1_r12_c5_rr6 = t0_r12_c5_rr12 + t0_r12_c5_rr13;
  assign t1_r12_c5_rr7 = t0_r12_c5_rr14;

  assign t2_r12_c5_rr0 = t1_r12_c5_rr0 + t1_r12_c5_rr1;
  assign t2_r12_c5_rr1 = t1_r12_c5_rr2 + t1_r12_c5_rr3;
  assign t2_r12_c5_rr2 = t1_r12_c5_rr4 + t1_r12_c5_rr5;
  assign t2_r12_c5_rr3 = t1_r12_c5_rr6 + t1_r12_c5_rr7;

  assign t3_r12_c5_rr0 = t2_r12_c5_rr0 + t2_r12_c5_rr1;
  assign t3_r12_c5_rr1 = t2_r12_c5_rr2 + t2_r12_c5_rr3;

  assign t4_r12_c5_rr0 = t3_r12_c5_rr0 + t3_r12_c5_rr1;

  assign c_12_5 = t4_r12_c5_rr0;
  assign t0_r12_c6_rr0 = a_12_0 * b_0_6;
  assign t0_r12_c6_rr1 = a_12_1 * b_1_6;
  assign t0_r12_c6_rr2 = a_12_2 * b_2_6;
  assign t0_r12_c6_rr3 = a_12_3 * b_3_6;
  assign t0_r12_c6_rr4 = a_12_4 * b_4_6;
  assign t0_r12_c6_rr5 = a_12_5 * b_5_6;
  assign t0_r12_c6_rr6 = a_12_6 * b_6_6;
  assign t0_r12_c6_rr7 = a_12_7 * b_7_6;
  assign t0_r12_c6_rr8 = a_12_8 * b_8_6;
  assign t0_r12_c6_rr9 = a_12_9 * b_9_6;
  assign t0_r12_c6_rr10 = a_12_10 * b_10_6;
  assign t0_r12_c6_rr11 = a_12_11 * b_11_6;
  assign t0_r12_c6_rr12 = a_12_12 * b_12_6;
  assign t0_r12_c6_rr13 = a_12_13 * b_13_6;
  assign t0_r12_c6_rr14 = a_12_14 * b_14_6;
  assign t1_r12_c6_rr0 = t0_r12_c6_rr0 + t0_r12_c6_rr1;
  assign t1_r12_c6_rr1 = t0_r12_c6_rr2 + t0_r12_c6_rr3;
  assign t1_r12_c6_rr2 = t0_r12_c6_rr4 + t0_r12_c6_rr5;
  assign t1_r12_c6_rr3 = t0_r12_c6_rr6 + t0_r12_c6_rr7;
  assign t1_r12_c6_rr4 = t0_r12_c6_rr8 + t0_r12_c6_rr9;
  assign t1_r12_c6_rr5 = t0_r12_c6_rr10 + t0_r12_c6_rr11;
  assign t1_r12_c6_rr6 = t0_r12_c6_rr12 + t0_r12_c6_rr13;
  assign t1_r12_c6_rr7 = t0_r12_c6_rr14;

  assign t2_r12_c6_rr0 = t1_r12_c6_rr0 + t1_r12_c6_rr1;
  assign t2_r12_c6_rr1 = t1_r12_c6_rr2 + t1_r12_c6_rr3;
  assign t2_r12_c6_rr2 = t1_r12_c6_rr4 + t1_r12_c6_rr5;
  assign t2_r12_c6_rr3 = t1_r12_c6_rr6 + t1_r12_c6_rr7;

  assign t3_r12_c6_rr0 = t2_r12_c6_rr0 + t2_r12_c6_rr1;
  assign t3_r12_c6_rr1 = t2_r12_c6_rr2 + t2_r12_c6_rr3;

  assign t4_r12_c6_rr0 = t3_r12_c6_rr0 + t3_r12_c6_rr1;

  assign c_12_6 = t4_r12_c6_rr0;
  assign t0_r12_c7_rr0 = a_12_0 * b_0_7;
  assign t0_r12_c7_rr1 = a_12_1 * b_1_7;
  assign t0_r12_c7_rr2 = a_12_2 * b_2_7;
  assign t0_r12_c7_rr3 = a_12_3 * b_3_7;
  assign t0_r12_c7_rr4 = a_12_4 * b_4_7;
  assign t0_r12_c7_rr5 = a_12_5 * b_5_7;
  assign t0_r12_c7_rr6 = a_12_6 * b_6_7;
  assign t0_r12_c7_rr7 = a_12_7 * b_7_7;
  assign t0_r12_c7_rr8 = a_12_8 * b_8_7;
  assign t0_r12_c7_rr9 = a_12_9 * b_9_7;
  assign t0_r12_c7_rr10 = a_12_10 * b_10_7;
  assign t0_r12_c7_rr11 = a_12_11 * b_11_7;
  assign t0_r12_c7_rr12 = a_12_12 * b_12_7;
  assign t0_r12_c7_rr13 = a_12_13 * b_13_7;
  assign t0_r12_c7_rr14 = a_12_14 * b_14_7;
  assign t1_r12_c7_rr0 = t0_r12_c7_rr0 + t0_r12_c7_rr1;
  assign t1_r12_c7_rr1 = t0_r12_c7_rr2 + t0_r12_c7_rr3;
  assign t1_r12_c7_rr2 = t0_r12_c7_rr4 + t0_r12_c7_rr5;
  assign t1_r12_c7_rr3 = t0_r12_c7_rr6 + t0_r12_c7_rr7;
  assign t1_r12_c7_rr4 = t0_r12_c7_rr8 + t0_r12_c7_rr9;
  assign t1_r12_c7_rr5 = t0_r12_c7_rr10 + t0_r12_c7_rr11;
  assign t1_r12_c7_rr6 = t0_r12_c7_rr12 + t0_r12_c7_rr13;
  assign t1_r12_c7_rr7 = t0_r12_c7_rr14;

  assign t2_r12_c7_rr0 = t1_r12_c7_rr0 + t1_r12_c7_rr1;
  assign t2_r12_c7_rr1 = t1_r12_c7_rr2 + t1_r12_c7_rr3;
  assign t2_r12_c7_rr2 = t1_r12_c7_rr4 + t1_r12_c7_rr5;
  assign t2_r12_c7_rr3 = t1_r12_c7_rr6 + t1_r12_c7_rr7;

  assign t3_r12_c7_rr0 = t2_r12_c7_rr0 + t2_r12_c7_rr1;
  assign t3_r12_c7_rr1 = t2_r12_c7_rr2 + t2_r12_c7_rr3;

  assign t4_r12_c7_rr0 = t3_r12_c7_rr0 + t3_r12_c7_rr1;

  assign c_12_7 = t4_r12_c7_rr0;
  assign t0_r12_c8_rr0 = a_12_0 * b_0_8;
  assign t0_r12_c8_rr1 = a_12_1 * b_1_8;
  assign t0_r12_c8_rr2 = a_12_2 * b_2_8;
  assign t0_r12_c8_rr3 = a_12_3 * b_3_8;
  assign t0_r12_c8_rr4 = a_12_4 * b_4_8;
  assign t0_r12_c8_rr5 = a_12_5 * b_5_8;
  assign t0_r12_c8_rr6 = a_12_6 * b_6_8;
  assign t0_r12_c8_rr7 = a_12_7 * b_7_8;
  assign t0_r12_c8_rr8 = a_12_8 * b_8_8;
  assign t0_r12_c8_rr9 = a_12_9 * b_9_8;
  assign t0_r12_c8_rr10 = a_12_10 * b_10_8;
  assign t0_r12_c8_rr11 = a_12_11 * b_11_8;
  assign t0_r12_c8_rr12 = a_12_12 * b_12_8;
  assign t0_r12_c8_rr13 = a_12_13 * b_13_8;
  assign t0_r12_c8_rr14 = a_12_14 * b_14_8;
  assign t1_r12_c8_rr0 = t0_r12_c8_rr0 + t0_r12_c8_rr1;
  assign t1_r12_c8_rr1 = t0_r12_c8_rr2 + t0_r12_c8_rr3;
  assign t1_r12_c8_rr2 = t0_r12_c8_rr4 + t0_r12_c8_rr5;
  assign t1_r12_c8_rr3 = t0_r12_c8_rr6 + t0_r12_c8_rr7;
  assign t1_r12_c8_rr4 = t0_r12_c8_rr8 + t0_r12_c8_rr9;
  assign t1_r12_c8_rr5 = t0_r12_c8_rr10 + t0_r12_c8_rr11;
  assign t1_r12_c8_rr6 = t0_r12_c8_rr12 + t0_r12_c8_rr13;
  assign t1_r12_c8_rr7 = t0_r12_c8_rr14;

  assign t2_r12_c8_rr0 = t1_r12_c8_rr0 + t1_r12_c8_rr1;
  assign t2_r12_c8_rr1 = t1_r12_c8_rr2 + t1_r12_c8_rr3;
  assign t2_r12_c8_rr2 = t1_r12_c8_rr4 + t1_r12_c8_rr5;
  assign t2_r12_c8_rr3 = t1_r12_c8_rr6 + t1_r12_c8_rr7;

  assign t3_r12_c8_rr0 = t2_r12_c8_rr0 + t2_r12_c8_rr1;
  assign t3_r12_c8_rr1 = t2_r12_c8_rr2 + t2_r12_c8_rr3;

  assign t4_r12_c8_rr0 = t3_r12_c8_rr0 + t3_r12_c8_rr1;

  assign c_12_8 = t4_r12_c8_rr0;
  assign t0_r12_c9_rr0 = a_12_0 * b_0_9;
  assign t0_r12_c9_rr1 = a_12_1 * b_1_9;
  assign t0_r12_c9_rr2 = a_12_2 * b_2_9;
  assign t0_r12_c9_rr3 = a_12_3 * b_3_9;
  assign t0_r12_c9_rr4 = a_12_4 * b_4_9;
  assign t0_r12_c9_rr5 = a_12_5 * b_5_9;
  assign t0_r12_c9_rr6 = a_12_6 * b_6_9;
  assign t0_r12_c9_rr7 = a_12_7 * b_7_9;
  assign t0_r12_c9_rr8 = a_12_8 * b_8_9;
  assign t0_r12_c9_rr9 = a_12_9 * b_9_9;
  assign t0_r12_c9_rr10 = a_12_10 * b_10_9;
  assign t0_r12_c9_rr11 = a_12_11 * b_11_9;
  assign t0_r12_c9_rr12 = a_12_12 * b_12_9;
  assign t0_r12_c9_rr13 = a_12_13 * b_13_9;
  assign t0_r12_c9_rr14 = a_12_14 * b_14_9;
  assign t1_r12_c9_rr0 = t0_r12_c9_rr0 + t0_r12_c9_rr1;
  assign t1_r12_c9_rr1 = t0_r12_c9_rr2 + t0_r12_c9_rr3;
  assign t1_r12_c9_rr2 = t0_r12_c9_rr4 + t0_r12_c9_rr5;
  assign t1_r12_c9_rr3 = t0_r12_c9_rr6 + t0_r12_c9_rr7;
  assign t1_r12_c9_rr4 = t0_r12_c9_rr8 + t0_r12_c9_rr9;
  assign t1_r12_c9_rr5 = t0_r12_c9_rr10 + t0_r12_c9_rr11;
  assign t1_r12_c9_rr6 = t0_r12_c9_rr12 + t0_r12_c9_rr13;
  assign t1_r12_c9_rr7 = t0_r12_c9_rr14;

  assign t2_r12_c9_rr0 = t1_r12_c9_rr0 + t1_r12_c9_rr1;
  assign t2_r12_c9_rr1 = t1_r12_c9_rr2 + t1_r12_c9_rr3;
  assign t2_r12_c9_rr2 = t1_r12_c9_rr4 + t1_r12_c9_rr5;
  assign t2_r12_c9_rr3 = t1_r12_c9_rr6 + t1_r12_c9_rr7;

  assign t3_r12_c9_rr0 = t2_r12_c9_rr0 + t2_r12_c9_rr1;
  assign t3_r12_c9_rr1 = t2_r12_c9_rr2 + t2_r12_c9_rr3;

  assign t4_r12_c9_rr0 = t3_r12_c9_rr0 + t3_r12_c9_rr1;

  assign c_12_9 = t4_r12_c9_rr0;
  assign t0_r12_c10_rr0 = a_12_0 * b_0_10;
  assign t0_r12_c10_rr1 = a_12_1 * b_1_10;
  assign t0_r12_c10_rr2 = a_12_2 * b_2_10;
  assign t0_r12_c10_rr3 = a_12_3 * b_3_10;
  assign t0_r12_c10_rr4 = a_12_4 * b_4_10;
  assign t0_r12_c10_rr5 = a_12_5 * b_5_10;
  assign t0_r12_c10_rr6 = a_12_6 * b_6_10;
  assign t0_r12_c10_rr7 = a_12_7 * b_7_10;
  assign t0_r12_c10_rr8 = a_12_8 * b_8_10;
  assign t0_r12_c10_rr9 = a_12_9 * b_9_10;
  assign t0_r12_c10_rr10 = a_12_10 * b_10_10;
  assign t0_r12_c10_rr11 = a_12_11 * b_11_10;
  assign t0_r12_c10_rr12 = a_12_12 * b_12_10;
  assign t0_r12_c10_rr13 = a_12_13 * b_13_10;
  assign t0_r12_c10_rr14 = a_12_14 * b_14_10;
  assign t1_r12_c10_rr0 = t0_r12_c10_rr0 + t0_r12_c10_rr1;
  assign t1_r12_c10_rr1 = t0_r12_c10_rr2 + t0_r12_c10_rr3;
  assign t1_r12_c10_rr2 = t0_r12_c10_rr4 + t0_r12_c10_rr5;
  assign t1_r12_c10_rr3 = t0_r12_c10_rr6 + t0_r12_c10_rr7;
  assign t1_r12_c10_rr4 = t0_r12_c10_rr8 + t0_r12_c10_rr9;
  assign t1_r12_c10_rr5 = t0_r12_c10_rr10 + t0_r12_c10_rr11;
  assign t1_r12_c10_rr6 = t0_r12_c10_rr12 + t0_r12_c10_rr13;
  assign t1_r12_c10_rr7 = t0_r12_c10_rr14;

  assign t2_r12_c10_rr0 = t1_r12_c10_rr0 + t1_r12_c10_rr1;
  assign t2_r12_c10_rr1 = t1_r12_c10_rr2 + t1_r12_c10_rr3;
  assign t2_r12_c10_rr2 = t1_r12_c10_rr4 + t1_r12_c10_rr5;
  assign t2_r12_c10_rr3 = t1_r12_c10_rr6 + t1_r12_c10_rr7;

  assign t3_r12_c10_rr0 = t2_r12_c10_rr0 + t2_r12_c10_rr1;
  assign t3_r12_c10_rr1 = t2_r12_c10_rr2 + t2_r12_c10_rr3;

  assign t4_r12_c10_rr0 = t3_r12_c10_rr0 + t3_r12_c10_rr1;

  assign c_12_10 = t4_r12_c10_rr0;
  assign t0_r12_c11_rr0 = a_12_0 * b_0_11;
  assign t0_r12_c11_rr1 = a_12_1 * b_1_11;
  assign t0_r12_c11_rr2 = a_12_2 * b_2_11;
  assign t0_r12_c11_rr3 = a_12_3 * b_3_11;
  assign t0_r12_c11_rr4 = a_12_4 * b_4_11;
  assign t0_r12_c11_rr5 = a_12_5 * b_5_11;
  assign t0_r12_c11_rr6 = a_12_6 * b_6_11;
  assign t0_r12_c11_rr7 = a_12_7 * b_7_11;
  assign t0_r12_c11_rr8 = a_12_8 * b_8_11;
  assign t0_r12_c11_rr9 = a_12_9 * b_9_11;
  assign t0_r12_c11_rr10 = a_12_10 * b_10_11;
  assign t0_r12_c11_rr11 = a_12_11 * b_11_11;
  assign t0_r12_c11_rr12 = a_12_12 * b_12_11;
  assign t0_r12_c11_rr13 = a_12_13 * b_13_11;
  assign t0_r12_c11_rr14 = a_12_14 * b_14_11;
  assign t1_r12_c11_rr0 = t0_r12_c11_rr0 + t0_r12_c11_rr1;
  assign t1_r12_c11_rr1 = t0_r12_c11_rr2 + t0_r12_c11_rr3;
  assign t1_r12_c11_rr2 = t0_r12_c11_rr4 + t0_r12_c11_rr5;
  assign t1_r12_c11_rr3 = t0_r12_c11_rr6 + t0_r12_c11_rr7;
  assign t1_r12_c11_rr4 = t0_r12_c11_rr8 + t0_r12_c11_rr9;
  assign t1_r12_c11_rr5 = t0_r12_c11_rr10 + t0_r12_c11_rr11;
  assign t1_r12_c11_rr6 = t0_r12_c11_rr12 + t0_r12_c11_rr13;
  assign t1_r12_c11_rr7 = t0_r12_c11_rr14;

  assign t2_r12_c11_rr0 = t1_r12_c11_rr0 + t1_r12_c11_rr1;
  assign t2_r12_c11_rr1 = t1_r12_c11_rr2 + t1_r12_c11_rr3;
  assign t2_r12_c11_rr2 = t1_r12_c11_rr4 + t1_r12_c11_rr5;
  assign t2_r12_c11_rr3 = t1_r12_c11_rr6 + t1_r12_c11_rr7;

  assign t3_r12_c11_rr0 = t2_r12_c11_rr0 + t2_r12_c11_rr1;
  assign t3_r12_c11_rr1 = t2_r12_c11_rr2 + t2_r12_c11_rr3;

  assign t4_r12_c11_rr0 = t3_r12_c11_rr0 + t3_r12_c11_rr1;

  assign c_12_11 = t4_r12_c11_rr0;
  assign t0_r12_c12_rr0 = a_12_0 * b_0_12;
  assign t0_r12_c12_rr1 = a_12_1 * b_1_12;
  assign t0_r12_c12_rr2 = a_12_2 * b_2_12;
  assign t0_r12_c12_rr3 = a_12_3 * b_3_12;
  assign t0_r12_c12_rr4 = a_12_4 * b_4_12;
  assign t0_r12_c12_rr5 = a_12_5 * b_5_12;
  assign t0_r12_c12_rr6 = a_12_6 * b_6_12;
  assign t0_r12_c12_rr7 = a_12_7 * b_7_12;
  assign t0_r12_c12_rr8 = a_12_8 * b_8_12;
  assign t0_r12_c12_rr9 = a_12_9 * b_9_12;
  assign t0_r12_c12_rr10 = a_12_10 * b_10_12;
  assign t0_r12_c12_rr11 = a_12_11 * b_11_12;
  assign t0_r12_c12_rr12 = a_12_12 * b_12_12;
  assign t0_r12_c12_rr13 = a_12_13 * b_13_12;
  assign t0_r12_c12_rr14 = a_12_14 * b_14_12;
  assign t1_r12_c12_rr0 = t0_r12_c12_rr0 + t0_r12_c12_rr1;
  assign t1_r12_c12_rr1 = t0_r12_c12_rr2 + t0_r12_c12_rr3;
  assign t1_r12_c12_rr2 = t0_r12_c12_rr4 + t0_r12_c12_rr5;
  assign t1_r12_c12_rr3 = t0_r12_c12_rr6 + t0_r12_c12_rr7;
  assign t1_r12_c12_rr4 = t0_r12_c12_rr8 + t0_r12_c12_rr9;
  assign t1_r12_c12_rr5 = t0_r12_c12_rr10 + t0_r12_c12_rr11;
  assign t1_r12_c12_rr6 = t0_r12_c12_rr12 + t0_r12_c12_rr13;
  assign t1_r12_c12_rr7 = t0_r12_c12_rr14;

  assign t2_r12_c12_rr0 = t1_r12_c12_rr0 + t1_r12_c12_rr1;
  assign t2_r12_c12_rr1 = t1_r12_c12_rr2 + t1_r12_c12_rr3;
  assign t2_r12_c12_rr2 = t1_r12_c12_rr4 + t1_r12_c12_rr5;
  assign t2_r12_c12_rr3 = t1_r12_c12_rr6 + t1_r12_c12_rr7;

  assign t3_r12_c12_rr0 = t2_r12_c12_rr0 + t2_r12_c12_rr1;
  assign t3_r12_c12_rr1 = t2_r12_c12_rr2 + t2_r12_c12_rr3;

  assign t4_r12_c12_rr0 = t3_r12_c12_rr0 + t3_r12_c12_rr1;

  assign c_12_12 = t4_r12_c12_rr0;
  assign t0_r12_c13_rr0 = a_12_0 * b_0_13;
  assign t0_r12_c13_rr1 = a_12_1 * b_1_13;
  assign t0_r12_c13_rr2 = a_12_2 * b_2_13;
  assign t0_r12_c13_rr3 = a_12_3 * b_3_13;
  assign t0_r12_c13_rr4 = a_12_4 * b_4_13;
  assign t0_r12_c13_rr5 = a_12_5 * b_5_13;
  assign t0_r12_c13_rr6 = a_12_6 * b_6_13;
  assign t0_r12_c13_rr7 = a_12_7 * b_7_13;
  assign t0_r12_c13_rr8 = a_12_8 * b_8_13;
  assign t0_r12_c13_rr9 = a_12_9 * b_9_13;
  assign t0_r12_c13_rr10 = a_12_10 * b_10_13;
  assign t0_r12_c13_rr11 = a_12_11 * b_11_13;
  assign t0_r12_c13_rr12 = a_12_12 * b_12_13;
  assign t0_r12_c13_rr13 = a_12_13 * b_13_13;
  assign t0_r12_c13_rr14 = a_12_14 * b_14_13;
  assign t1_r12_c13_rr0 = t0_r12_c13_rr0 + t0_r12_c13_rr1;
  assign t1_r12_c13_rr1 = t0_r12_c13_rr2 + t0_r12_c13_rr3;
  assign t1_r12_c13_rr2 = t0_r12_c13_rr4 + t0_r12_c13_rr5;
  assign t1_r12_c13_rr3 = t0_r12_c13_rr6 + t0_r12_c13_rr7;
  assign t1_r12_c13_rr4 = t0_r12_c13_rr8 + t0_r12_c13_rr9;
  assign t1_r12_c13_rr5 = t0_r12_c13_rr10 + t0_r12_c13_rr11;
  assign t1_r12_c13_rr6 = t0_r12_c13_rr12 + t0_r12_c13_rr13;
  assign t1_r12_c13_rr7 = t0_r12_c13_rr14;

  assign t2_r12_c13_rr0 = t1_r12_c13_rr0 + t1_r12_c13_rr1;
  assign t2_r12_c13_rr1 = t1_r12_c13_rr2 + t1_r12_c13_rr3;
  assign t2_r12_c13_rr2 = t1_r12_c13_rr4 + t1_r12_c13_rr5;
  assign t2_r12_c13_rr3 = t1_r12_c13_rr6 + t1_r12_c13_rr7;

  assign t3_r12_c13_rr0 = t2_r12_c13_rr0 + t2_r12_c13_rr1;
  assign t3_r12_c13_rr1 = t2_r12_c13_rr2 + t2_r12_c13_rr3;

  assign t4_r12_c13_rr0 = t3_r12_c13_rr0 + t3_r12_c13_rr1;

  assign c_12_13 = t4_r12_c13_rr0;
  assign t0_r12_c14_rr0 = a_12_0 * b_0_14;
  assign t0_r12_c14_rr1 = a_12_1 * b_1_14;
  assign t0_r12_c14_rr2 = a_12_2 * b_2_14;
  assign t0_r12_c14_rr3 = a_12_3 * b_3_14;
  assign t0_r12_c14_rr4 = a_12_4 * b_4_14;
  assign t0_r12_c14_rr5 = a_12_5 * b_5_14;
  assign t0_r12_c14_rr6 = a_12_6 * b_6_14;
  assign t0_r12_c14_rr7 = a_12_7 * b_7_14;
  assign t0_r12_c14_rr8 = a_12_8 * b_8_14;
  assign t0_r12_c14_rr9 = a_12_9 * b_9_14;
  assign t0_r12_c14_rr10 = a_12_10 * b_10_14;
  assign t0_r12_c14_rr11 = a_12_11 * b_11_14;
  assign t0_r12_c14_rr12 = a_12_12 * b_12_14;
  assign t0_r12_c14_rr13 = a_12_13 * b_13_14;
  assign t0_r12_c14_rr14 = a_12_14 * b_14_14;
  assign t1_r12_c14_rr0 = t0_r12_c14_rr0 + t0_r12_c14_rr1;
  assign t1_r12_c14_rr1 = t0_r12_c14_rr2 + t0_r12_c14_rr3;
  assign t1_r12_c14_rr2 = t0_r12_c14_rr4 + t0_r12_c14_rr5;
  assign t1_r12_c14_rr3 = t0_r12_c14_rr6 + t0_r12_c14_rr7;
  assign t1_r12_c14_rr4 = t0_r12_c14_rr8 + t0_r12_c14_rr9;
  assign t1_r12_c14_rr5 = t0_r12_c14_rr10 + t0_r12_c14_rr11;
  assign t1_r12_c14_rr6 = t0_r12_c14_rr12 + t0_r12_c14_rr13;
  assign t1_r12_c14_rr7 = t0_r12_c14_rr14;

  assign t2_r12_c14_rr0 = t1_r12_c14_rr0 + t1_r12_c14_rr1;
  assign t2_r12_c14_rr1 = t1_r12_c14_rr2 + t1_r12_c14_rr3;
  assign t2_r12_c14_rr2 = t1_r12_c14_rr4 + t1_r12_c14_rr5;
  assign t2_r12_c14_rr3 = t1_r12_c14_rr6 + t1_r12_c14_rr7;

  assign t3_r12_c14_rr0 = t2_r12_c14_rr0 + t2_r12_c14_rr1;
  assign t3_r12_c14_rr1 = t2_r12_c14_rr2 + t2_r12_c14_rr3;

  assign t4_r12_c14_rr0 = t3_r12_c14_rr0 + t3_r12_c14_rr1;

  assign c_12_14 = t4_r12_c14_rr0;
  assign t0_r13_c0_rr0 = a_13_0 * b_0_0;
  assign t0_r13_c0_rr1 = a_13_1 * b_1_0;
  assign t0_r13_c0_rr2 = a_13_2 * b_2_0;
  assign t0_r13_c0_rr3 = a_13_3 * b_3_0;
  assign t0_r13_c0_rr4 = a_13_4 * b_4_0;
  assign t0_r13_c0_rr5 = a_13_5 * b_5_0;
  assign t0_r13_c0_rr6 = a_13_6 * b_6_0;
  assign t0_r13_c0_rr7 = a_13_7 * b_7_0;
  assign t0_r13_c0_rr8 = a_13_8 * b_8_0;
  assign t0_r13_c0_rr9 = a_13_9 * b_9_0;
  assign t0_r13_c0_rr10 = a_13_10 * b_10_0;
  assign t0_r13_c0_rr11 = a_13_11 * b_11_0;
  assign t0_r13_c0_rr12 = a_13_12 * b_12_0;
  assign t0_r13_c0_rr13 = a_13_13 * b_13_0;
  assign t0_r13_c0_rr14 = a_13_14 * b_14_0;
  assign t1_r13_c0_rr0 = t0_r13_c0_rr0 + t0_r13_c0_rr1;
  assign t1_r13_c0_rr1 = t0_r13_c0_rr2 + t0_r13_c0_rr3;
  assign t1_r13_c0_rr2 = t0_r13_c0_rr4 + t0_r13_c0_rr5;
  assign t1_r13_c0_rr3 = t0_r13_c0_rr6 + t0_r13_c0_rr7;
  assign t1_r13_c0_rr4 = t0_r13_c0_rr8 + t0_r13_c0_rr9;
  assign t1_r13_c0_rr5 = t0_r13_c0_rr10 + t0_r13_c0_rr11;
  assign t1_r13_c0_rr6 = t0_r13_c0_rr12 + t0_r13_c0_rr13;
  assign t1_r13_c0_rr7 = t0_r13_c0_rr14;

  assign t2_r13_c0_rr0 = t1_r13_c0_rr0 + t1_r13_c0_rr1;
  assign t2_r13_c0_rr1 = t1_r13_c0_rr2 + t1_r13_c0_rr3;
  assign t2_r13_c0_rr2 = t1_r13_c0_rr4 + t1_r13_c0_rr5;
  assign t2_r13_c0_rr3 = t1_r13_c0_rr6 + t1_r13_c0_rr7;

  assign t3_r13_c0_rr0 = t2_r13_c0_rr0 + t2_r13_c0_rr1;
  assign t3_r13_c0_rr1 = t2_r13_c0_rr2 + t2_r13_c0_rr3;

  assign t4_r13_c0_rr0 = t3_r13_c0_rr0 + t3_r13_c0_rr1;

  assign c_13_0 = t4_r13_c0_rr0;
  assign t0_r13_c1_rr0 = a_13_0 * b_0_1;
  assign t0_r13_c1_rr1 = a_13_1 * b_1_1;
  assign t0_r13_c1_rr2 = a_13_2 * b_2_1;
  assign t0_r13_c1_rr3 = a_13_3 * b_3_1;
  assign t0_r13_c1_rr4 = a_13_4 * b_4_1;
  assign t0_r13_c1_rr5 = a_13_5 * b_5_1;
  assign t0_r13_c1_rr6 = a_13_6 * b_6_1;
  assign t0_r13_c1_rr7 = a_13_7 * b_7_1;
  assign t0_r13_c1_rr8 = a_13_8 * b_8_1;
  assign t0_r13_c1_rr9 = a_13_9 * b_9_1;
  assign t0_r13_c1_rr10 = a_13_10 * b_10_1;
  assign t0_r13_c1_rr11 = a_13_11 * b_11_1;
  assign t0_r13_c1_rr12 = a_13_12 * b_12_1;
  assign t0_r13_c1_rr13 = a_13_13 * b_13_1;
  assign t0_r13_c1_rr14 = a_13_14 * b_14_1;
  assign t1_r13_c1_rr0 = t0_r13_c1_rr0 + t0_r13_c1_rr1;
  assign t1_r13_c1_rr1 = t0_r13_c1_rr2 + t0_r13_c1_rr3;
  assign t1_r13_c1_rr2 = t0_r13_c1_rr4 + t0_r13_c1_rr5;
  assign t1_r13_c1_rr3 = t0_r13_c1_rr6 + t0_r13_c1_rr7;
  assign t1_r13_c1_rr4 = t0_r13_c1_rr8 + t0_r13_c1_rr9;
  assign t1_r13_c1_rr5 = t0_r13_c1_rr10 + t0_r13_c1_rr11;
  assign t1_r13_c1_rr6 = t0_r13_c1_rr12 + t0_r13_c1_rr13;
  assign t1_r13_c1_rr7 = t0_r13_c1_rr14;

  assign t2_r13_c1_rr0 = t1_r13_c1_rr0 + t1_r13_c1_rr1;
  assign t2_r13_c1_rr1 = t1_r13_c1_rr2 + t1_r13_c1_rr3;
  assign t2_r13_c1_rr2 = t1_r13_c1_rr4 + t1_r13_c1_rr5;
  assign t2_r13_c1_rr3 = t1_r13_c1_rr6 + t1_r13_c1_rr7;

  assign t3_r13_c1_rr0 = t2_r13_c1_rr0 + t2_r13_c1_rr1;
  assign t3_r13_c1_rr1 = t2_r13_c1_rr2 + t2_r13_c1_rr3;

  assign t4_r13_c1_rr0 = t3_r13_c1_rr0 + t3_r13_c1_rr1;

  assign c_13_1 = t4_r13_c1_rr0;
  assign t0_r13_c2_rr0 = a_13_0 * b_0_2;
  assign t0_r13_c2_rr1 = a_13_1 * b_1_2;
  assign t0_r13_c2_rr2 = a_13_2 * b_2_2;
  assign t0_r13_c2_rr3 = a_13_3 * b_3_2;
  assign t0_r13_c2_rr4 = a_13_4 * b_4_2;
  assign t0_r13_c2_rr5 = a_13_5 * b_5_2;
  assign t0_r13_c2_rr6 = a_13_6 * b_6_2;
  assign t0_r13_c2_rr7 = a_13_7 * b_7_2;
  assign t0_r13_c2_rr8 = a_13_8 * b_8_2;
  assign t0_r13_c2_rr9 = a_13_9 * b_9_2;
  assign t0_r13_c2_rr10 = a_13_10 * b_10_2;
  assign t0_r13_c2_rr11 = a_13_11 * b_11_2;
  assign t0_r13_c2_rr12 = a_13_12 * b_12_2;
  assign t0_r13_c2_rr13 = a_13_13 * b_13_2;
  assign t0_r13_c2_rr14 = a_13_14 * b_14_2;
  assign t1_r13_c2_rr0 = t0_r13_c2_rr0 + t0_r13_c2_rr1;
  assign t1_r13_c2_rr1 = t0_r13_c2_rr2 + t0_r13_c2_rr3;
  assign t1_r13_c2_rr2 = t0_r13_c2_rr4 + t0_r13_c2_rr5;
  assign t1_r13_c2_rr3 = t0_r13_c2_rr6 + t0_r13_c2_rr7;
  assign t1_r13_c2_rr4 = t0_r13_c2_rr8 + t0_r13_c2_rr9;
  assign t1_r13_c2_rr5 = t0_r13_c2_rr10 + t0_r13_c2_rr11;
  assign t1_r13_c2_rr6 = t0_r13_c2_rr12 + t0_r13_c2_rr13;
  assign t1_r13_c2_rr7 = t0_r13_c2_rr14;

  assign t2_r13_c2_rr0 = t1_r13_c2_rr0 + t1_r13_c2_rr1;
  assign t2_r13_c2_rr1 = t1_r13_c2_rr2 + t1_r13_c2_rr3;
  assign t2_r13_c2_rr2 = t1_r13_c2_rr4 + t1_r13_c2_rr5;
  assign t2_r13_c2_rr3 = t1_r13_c2_rr6 + t1_r13_c2_rr7;

  assign t3_r13_c2_rr0 = t2_r13_c2_rr0 + t2_r13_c2_rr1;
  assign t3_r13_c2_rr1 = t2_r13_c2_rr2 + t2_r13_c2_rr3;

  assign t4_r13_c2_rr0 = t3_r13_c2_rr0 + t3_r13_c2_rr1;

  assign c_13_2 = t4_r13_c2_rr0;
  assign t0_r13_c3_rr0 = a_13_0 * b_0_3;
  assign t0_r13_c3_rr1 = a_13_1 * b_1_3;
  assign t0_r13_c3_rr2 = a_13_2 * b_2_3;
  assign t0_r13_c3_rr3 = a_13_3 * b_3_3;
  assign t0_r13_c3_rr4 = a_13_4 * b_4_3;
  assign t0_r13_c3_rr5 = a_13_5 * b_5_3;
  assign t0_r13_c3_rr6 = a_13_6 * b_6_3;
  assign t0_r13_c3_rr7 = a_13_7 * b_7_3;
  assign t0_r13_c3_rr8 = a_13_8 * b_8_3;
  assign t0_r13_c3_rr9 = a_13_9 * b_9_3;
  assign t0_r13_c3_rr10 = a_13_10 * b_10_3;
  assign t0_r13_c3_rr11 = a_13_11 * b_11_3;
  assign t0_r13_c3_rr12 = a_13_12 * b_12_3;
  assign t0_r13_c3_rr13 = a_13_13 * b_13_3;
  assign t0_r13_c3_rr14 = a_13_14 * b_14_3;
  assign t1_r13_c3_rr0 = t0_r13_c3_rr0 + t0_r13_c3_rr1;
  assign t1_r13_c3_rr1 = t0_r13_c3_rr2 + t0_r13_c3_rr3;
  assign t1_r13_c3_rr2 = t0_r13_c3_rr4 + t0_r13_c3_rr5;
  assign t1_r13_c3_rr3 = t0_r13_c3_rr6 + t0_r13_c3_rr7;
  assign t1_r13_c3_rr4 = t0_r13_c3_rr8 + t0_r13_c3_rr9;
  assign t1_r13_c3_rr5 = t0_r13_c3_rr10 + t0_r13_c3_rr11;
  assign t1_r13_c3_rr6 = t0_r13_c3_rr12 + t0_r13_c3_rr13;
  assign t1_r13_c3_rr7 = t0_r13_c3_rr14;

  assign t2_r13_c3_rr0 = t1_r13_c3_rr0 + t1_r13_c3_rr1;
  assign t2_r13_c3_rr1 = t1_r13_c3_rr2 + t1_r13_c3_rr3;
  assign t2_r13_c3_rr2 = t1_r13_c3_rr4 + t1_r13_c3_rr5;
  assign t2_r13_c3_rr3 = t1_r13_c3_rr6 + t1_r13_c3_rr7;

  assign t3_r13_c3_rr0 = t2_r13_c3_rr0 + t2_r13_c3_rr1;
  assign t3_r13_c3_rr1 = t2_r13_c3_rr2 + t2_r13_c3_rr3;

  assign t4_r13_c3_rr0 = t3_r13_c3_rr0 + t3_r13_c3_rr1;

  assign c_13_3 = t4_r13_c3_rr0;
  assign t0_r13_c4_rr0 = a_13_0 * b_0_4;
  assign t0_r13_c4_rr1 = a_13_1 * b_1_4;
  assign t0_r13_c4_rr2 = a_13_2 * b_2_4;
  assign t0_r13_c4_rr3 = a_13_3 * b_3_4;
  assign t0_r13_c4_rr4 = a_13_4 * b_4_4;
  assign t0_r13_c4_rr5 = a_13_5 * b_5_4;
  assign t0_r13_c4_rr6 = a_13_6 * b_6_4;
  assign t0_r13_c4_rr7 = a_13_7 * b_7_4;
  assign t0_r13_c4_rr8 = a_13_8 * b_8_4;
  assign t0_r13_c4_rr9 = a_13_9 * b_9_4;
  assign t0_r13_c4_rr10 = a_13_10 * b_10_4;
  assign t0_r13_c4_rr11 = a_13_11 * b_11_4;
  assign t0_r13_c4_rr12 = a_13_12 * b_12_4;
  assign t0_r13_c4_rr13 = a_13_13 * b_13_4;
  assign t0_r13_c4_rr14 = a_13_14 * b_14_4;
  assign t1_r13_c4_rr0 = t0_r13_c4_rr0 + t0_r13_c4_rr1;
  assign t1_r13_c4_rr1 = t0_r13_c4_rr2 + t0_r13_c4_rr3;
  assign t1_r13_c4_rr2 = t0_r13_c4_rr4 + t0_r13_c4_rr5;
  assign t1_r13_c4_rr3 = t0_r13_c4_rr6 + t0_r13_c4_rr7;
  assign t1_r13_c4_rr4 = t0_r13_c4_rr8 + t0_r13_c4_rr9;
  assign t1_r13_c4_rr5 = t0_r13_c4_rr10 + t0_r13_c4_rr11;
  assign t1_r13_c4_rr6 = t0_r13_c4_rr12 + t0_r13_c4_rr13;
  assign t1_r13_c4_rr7 = t0_r13_c4_rr14;

  assign t2_r13_c4_rr0 = t1_r13_c4_rr0 + t1_r13_c4_rr1;
  assign t2_r13_c4_rr1 = t1_r13_c4_rr2 + t1_r13_c4_rr3;
  assign t2_r13_c4_rr2 = t1_r13_c4_rr4 + t1_r13_c4_rr5;
  assign t2_r13_c4_rr3 = t1_r13_c4_rr6 + t1_r13_c4_rr7;

  assign t3_r13_c4_rr0 = t2_r13_c4_rr0 + t2_r13_c4_rr1;
  assign t3_r13_c4_rr1 = t2_r13_c4_rr2 + t2_r13_c4_rr3;

  assign t4_r13_c4_rr0 = t3_r13_c4_rr0 + t3_r13_c4_rr1;

  assign c_13_4 = t4_r13_c4_rr0;
  assign t0_r13_c5_rr0 = a_13_0 * b_0_5;
  assign t0_r13_c5_rr1 = a_13_1 * b_1_5;
  assign t0_r13_c5_rr2 = a_13_2 * b_2_5;
  assign t0_r13_c5_rr3 = a_13_3 * b_3_5;
  assign t0_r13_c5_rr4 = a_13_4 * b_4_5;
  assign t0_r13_c5_rr5 = a_13_5 * b_5_5;
  assign t0_r13_c5_rr6 = a_13_6 * b_6_5;
  assign t0_r13_c5_rr7 = a_13_7 * b_7_5;
  assign t0_r13_c5_rr8 = a_13_8 * b_8_5;
  assign t0_r13_c5_rr9 = a_13_9 * b_9_5;
  assign t0_r13_c5_rr10 = a_13_10 * b_10_5;
  assign t0_r13_c5_rr11 = a_13_11 * b_11_5;
  assign t0_r13_c5_rr12 = a_13_12 * b_12_5;
  assign t0_r13_c5_rr13 = a_13_13 * b_13_5;
  assign t0_r13_c5_rr14 = a_13_14 * b_14_5;
  assign t1_r13_c5_rr0 = t0_r13_c5_rr0 + t0_r13_c5_rr1;
  assign t1_r13_c5_rr1 = t0_r13_c5_rr2 + t0_r13_c5_rr3;
  assign t1_r13_c5_rr2 = t0_r13_c5_rr4 + t0_r13_c5_rr5;
  assign t1_r13_c5_rr3 = t0_r13_c5_rr6 + t0_r13_c5_rr7;
  assign t1_r13_c5_rr4 = t0_r13_c5_rr8 + t0_r13_c5_rr9;
  assign t1_r13_c5_rr5 = t0_r13_c5_rr10 + t0_r13_c5_rr11;
  assign t1_r13_c5_rr6 = t0_r13_c5_rr12 + t0_r13_c5_rr13;
  assign t1_r13_c5_rr7 = t0_r13_c5_rr14;

  assign t2_r13_c5_rr0 = t1_r13_c5_rr0 + t1_r13_c5_rr1;
  assign t2_r13_c5_rr1 = t1_r13_c5_rr2 + t1_r13_c5_rr3;
  assign t2_r13_c5_rr2 = t1_r13_c5_rr4 + t1_r13_c5_rr5;
  assign t2_r13_c5_rr3 = t1_r13_c5_rr6 + t1_r13_c5_rr7;

  assign t3_r13_c5_rr0 = t2_r13_c5_rr0 + t2_r13_c5_rr1;
  assign t3_r13_c5_rr1 = t2_r13_c5_rr2 + t2_r13_c5_rr3;

  assign t4_r13_c5_rr0 = t3_r13_c5_rr0 + t3_r13_c5_rr1;

  assign c_13_5 = t4_r13_c5_rr0;
  assign t0_r13_c6_rr0 = a_13_0 * b_0_6;
  assign t0_r13_c6_rr1 = a_13_1 * b_1_6;
  assign t0_r13_c6_rr2 = a_13_2 * b_2_6;
  assign t0_r13_c6_rr3 = a_13_3 * b_3_6;
  assign t0_r13_c6_rr4 = a_13_4 * b_4_6;
  assign t0_r13_c6_rr5 = a_13_5 * b_5_6;
  assign t0_r13_c6_rr6 = a_13_6 * b_6_6;
  assign t0_r13_c6_rr7 = a_13_7 * b_7_6;
  assign t0_r13_c6_rr8 = a_13_8 * b_8_6;
  assign t0_r13_c6_rr9 = a_13_9 * b_9_6;
  assign t0_r13_c6_rr10 = a_13_10 * b_10_6;
  assign t0_r13_c6_rr11 = a_13_11 * b_11_6;
  assign t0_r13_c6_rr12 = a_13_12 * b_12_6;
  assign t0_r13_c6_rr13 = a_13_13 * b_13_6;
  assign t0_r13_c6_rr14 = a_13_14 * b_14_6;
  assign t1_r13_c6_rr0 = t0_r13_c6_rr0 + t0_r13_c6_rr1;
  assign t1_r13_c6_rr1 = t0_r13_c6_rr2 + t0_r13_c6_rr3;
  assign t1_r13_c6_rr2 = t0_r13_c6_rr4 + t0_r13_c6_rr5;
  assign t1_r13_c6_rr3 = t0_r13_c6_rr6 + t0_r13_c6_rr7;
  assign t1_r13_c6_rr4 = t0_r13_c6_rr8 + t0_r13_c6_rr9;
  assign t1_r13_c6_rr5 = t0_r13_c6_rr10 + t0_r13_c6_rr11;
  assign t1_r13_c6_rr6 = t0_r13_c6_rr12 + t0_r13_c6_rr13;
  assign t1_r13_c6_rr7 = t0_r13_c6_rr14;

  assign t2_r13_c6_rr0 = t1_r13_c6_rr0 + t1_r13_c6_rr1;
  assign t2_r13_c6_rr1 = t1_r13_c6_rr2 + t1_r13_c6_rr3;
  assign t2_r13_c6_rr2 = t1_r13_c6_rr4 + t1_r13_c6_rr5;
  assign t2_r13_c6_rr3 = t1_r13_c6_rr6 + t1_r13_c6_rr7;

  assign t3_r13_c6_rr0 = t2_r13_c6_rr0 + t2_r13_c6_rr1;
  assign t3_r13_c6_rr1 = t2_r13_c6_rr2 + t2_r13_c6_rr3;

  assign t4_r13_c6_rr0 = t3_r13_c6_rr0 + t3_r13_c6_rr1;

  assign c_13_6 = t4_r13_c6_rr0;
  assign t0_r13_c7_rr0 = a_13_0 * b_0_7;
  assign t0_r13_c7_rr1 = a_13_1 * b_1_7;
  assign t0_r13_c7_rr2 = a_13_2 * b_2_7;
  assign t0_r13_c7_rr3 = a_13_3 * b_3_7;
  assign t0_r13_c7_rr4 = a_13_4 * b_4_7;
  assign t0_r13_c7_rr5 = a_13_5 * b_5_7;
  assign t0_r13_c7_rr6 = a_13_6 * b_6_7;
  assign t0_r13_c7_rr7 = a_13_7 * b_7_7;
  assign t0_r13_c7_rr8 = a_13_8 * b_8_7;
  assign t0_r13_c7_rr9 = a_13_9 * b_9_7;
  assign t0_r13_c7_rr10 = a_13_10 * b_10_7;
  assign t0_r13_c7_rr11 = a_13_11 * b_11_7;
  assign t0_r13_c7_rr12 = a_13_12 * b_12_7;
  assign t0_r13_c7_rr13 = a_13_13 * b_13_7;
  assign t0_r13_c7_rr14 = a_13_14 * b_14_7;
  assign t1_r13_c7_rr0 = t0_r13_c7_rr0 + t0_r13_c7_rr1;
  assign t1_r13_c7_rr1 = t0_r13_c7_rr2 + t0_r13_c7_rr3;
  assign t1_r13_c7_rr2 = t0_r13_c7_rr4 + t0_r13_c7_rr5;
  assign t1_r13_c7_rr3 = t0_r13_c7_rr6 + t0_r13_c7_rr7;
  assign t1_r13_c7_rr4 = t0_r13_c7_rr8 + t0_r13_c7_rr9;
  assign t1_r13_c7_rr5 = t0_r13_c7_rr10 + t0_r13_c7_rr11;
  assign t1_r13_c7_rr6 = t0_r13_c7_rr12 + t0_r13_c7_rr13;
  assign t1_r13_c7_rr7 = t0_r13_c7_rr14;

  assign t2_r13_c7_rr0 = t1_r13_c7_rr0 + t1_r13_c7_rr1;
  assign t2_r13_c7_rr1 = t1_r13_c7_rr2 + t1_r13_c7_rr3;
  assign t2_r13_c7_rr2 = t1_r13_c7_rr4 + t1_r13_c7_rr5;
  assign t2_r13_c7_rr3 = t1_r13_c7_rr6 + t1_r13_c7_rr7;

  assign t3_r13_c7_rr0 = t2_r13_c7_rr0 + t2_r13_c7_rr1;
  assign t3_r13_c7_rr1 = t2_r13_c7_rr2 + t2_r13_c7_rr3;

  assign t4_r13_c7_rr0 = t3_r13_c7_rr0 + t3_r13_c7_rr1;

  assign c_13_7 = t4_r13_c7_rr0;
  assign t0_r13_c8_rr0 = a_13_0 * b_0_8;
  assign t0_r13_c8_rr1 = a_13_1 * b_1_8;
  assign t0_r13_c8_rr2 = a_13_2 * b_2_8;
  assign t0_r13_c8_rr3 = a_13_3 * b_3_8;
  assign t0_r13_c8_rr4 = a_13_4 * b_4_8;
  assign t0_r13_c8_rr5 = a_13_5 * b_5_8;
  assign t0_r13_c8_rr6 = a_13_6 * b_6_8;
  assign t0_r13_c8_rr7 = a_13_7 * b_7_8;
  assign t0_r13_c8_rr8 = a_13_8 * b_8_8;
  assign t0_r13_c8_rr9 = a_13_9 * b_9_8;
  assign t0_r13_c8_rr10 = a_13_10 * b_10_8;
  assign t0_r13_c8_rr11 = a_13_11 * b_11_8;
  assign t0_r13_c8_rr12 = a_13_12 * b_12_8;
  assign t0_r13_c8_rr13 = a_13_13 * b_13_8;
  assign t0_r13_c8_rr14 = a_13_14 * b_14_8;
  assign t1_r13_c8_rr0 = t0_r13_c8_rr0 + t0_r13_c8_rr1;
  assign t1_r13_c8_rr1 = t0_r13_c8_rr2 + t0_r13_c8_rr3;
  assign t1_r13_c8_rr2 = t0_r13_c8_rr4 + t0_r13_c8_rr5;
  assign t1_r13_c8_rr3 = t0_r13_c8_rr6 + t0_r13_c8_rr7;
  assign t1_r13_c8_rr4 = t0_r13_c8_rr8 + t0_r13_c8_rr9;
  assign t1_r13_c8_rr5 = t0_r13_c8_rr10 + t0_r13_c8_rr11;
  assign t1_r13_c8_rr6 = t0_r13_c8_rr12 + t0_r13_c8_rr13;
  assign t1_r13_c8_rr7 = t0_r13_c8_rr14;

  assign t2_r13_c8_rr0 = t1_r13_c8_rr0 + t1_r13_c8_rr1;
  assign t2_r13_c8_rr1 = t1_r13_c8_rr2 + t1_r13_c8_rr3;
  assign t2_r13_c8_rr2 = t1_r13_c8_rr4 + t1_r13_c8_rr5;
  assign t2_r13_c8_rr3 = t1_r13_c8_rr6 + t1_r13_c8_rr7;

  assign t3_r13_c8_rr0 = t2_r13_c8_rr0 + t2_r13_c8_rr1;
  assign t3_r13_c8_rr1 = t2_r13_c8_rr2 + t2_r13_c8_rr3;

  assign t4_r13_c8_rr0 = t3_r13_c8_rr0 + t3_r13_c8_rr1;

  assign c_13_8 = t4_r13_c8_rr0;
  assign t0_r13_c9_rr0 = a_13_0 * b_0_9;
  assign t0_r13_c9_rr1 = a_13_1 * b_1_9;
  assign t0_r13_c9_rr2 = a_13_2 * b_2_9;
  assign t0_r13_c9_rr3 = a_13_3 * b_3_9;
  assign t0_r13_c9_rr4 = a_13_4 * b_4_9;
  assign t0_r13_c9_rr5 = a_13_5 * b_5_9;
  assign t0_r13_c9_rr6 = a_13_6 * b_6_9;
  assign t0_r13_c9_rr7 = a_13_7 * b_7_9;
  assign t0_r13_c9_rr8 = a_13_8 * b_8_9;
  assign t0_r13_c9_rr9 = a_13_9 * b_9_9;
  assign t0_r13_c9_rr10 = a_13_10 * b_10_9;
  assign t0_r13_c9_rr11 = a_13_11 * b_11_9;
  assign t0_r13_c9_rr12 = a_13_12 * b_12_9;
  assign t0_r13_c9_rr13 = a_13_13 * b_13_9;
  assign t0_r13_c9_rr14 = a_13_14 * b_14_9;
  assign t1_r13_c9_rr0 = t0_r13_c9_rr0 + t0_r13_c9_rr1;
  assign t1_r13_c9_rr1 = t0_r13_c9_rr2 + t0_r13_c9_rr3;
  assign t1_r13_c9_rr2 = t0_r13_c9_rr4 + t0_r13_c9_rr5;
  assign t1_r13_c9_rr3 = t0_r13_c9_rr6 + t0_r13_c9_rr7;
  assign t1_r13_c9_rr4 = t0_r13_c9_rr8 + t0_r13_c9_rr9;
  assign t1_r13_c9_rr5 = t0_r13_c9_rr10 + t0_r13_c9_rr11;
  assign t1_r13_c9_rr6 = t0_r13_c9_rr12 + t0_r13_c9_rr13;
  assign t1_r13_c9_rr7 = t0_r13_c9_rr14;

  assign t2_r13_c9_rr0 = t1_r13_c9_rr0 + t1_r13_c9_rr1;
  assign t2_r13_c9_rr1 = t1_r13_c9_rr2 + t1_r13_c9_rr3;
  assign t2_r13_c9_rr2 = t1_r13_c9_rr4 + t1_r13_c9_rr5;
  assign t2_r13_c9_rr3 = t1_r13_c9_rr6 + t1_r13_c9_rr7;

  assign t3_r13_c9_rr0 = t2_r13_c9_rr0 + t2_r13_c9_rr1;
  assign t3_r13_c9_rr1 = t2_r13_c9_rr2 + t2_r13_c9_rr3;

  assign t4_r13_c9_rr0 = t3_r13_c9_rr0 + t3_r13_c9_rr1;

  assign c_13_9 = t4_r13_c9_rr0;
  assign t0_r13_c10_rr0 = a_13_0 * b_0_10;
  assign t0_r13_c10_rr1 = a_13_1 * b_1_10;
  assign t0_r13_c10_rr2 = a_13_2 * b_2_10;
  assign t0_r13_c10_rr3 = a_13_3 * b_3_10;
  assign t0_r13_c10_rr4 = a_13_4 * b_4_10;
  assign t0_r13_c10_rr5 = a_13_5 * b_5_10;
  assign t0_r13_c10_rr6 = a_13_6 * b_6_10;
  assign t0_r13_c10_rr7 = a_13_7 * b_7_10;
  assign t0_r13_c10_rr8 = a_13_8 * b_8_10;
  assign t0_r13_c10_rr9 = a_13_9 * b_9_10;
  assign t0_r13_c10_rr10 = a_13_10 * b_10_10;
  assign t0_r13_c10_rr11 = a_13_11 * b_11_10;
  assign t0_r13_c10_rr12 = a_13_12 * b_12_10;
  assign t0_r13_c10_rr13 = a_13_13 * b_13_10;
  assign t0_r13_c10_rr14 = a_13_14 * b_14_10;
  assign t1_r13_c10_rr0 = t0_r13_c10_rr0 + t0_r13_c10_rr1;
  assign t1_r13_c10_rr1 = t0_r13_c10_rr2 + t0_r13_c10_rr3;
  assign t1_r13_c10_rr2 = t0_r13_c10_rr4 + t0_r13_c10_rr5;
  assign t1_r13_c10_rr3 = t0_r13_c10_rr6 + t0_r13_c10_rr7;
  assign t1_r13_c10_rr4 = t0_r13_c10_rr8 + t0_r13_c10_rr9;
  assign t1_r13_c10_rr5 = t0_r13_c10_rr10 + t0_r13_c10_rr11;
  assign t1_r13_c10_rr6 = t0_r13_c10_rr12 + t0_r13_c10_rr13;
  assign t1_r13_c10_rr7 = t0_r13_c10_rr14;

  assign t2_r13_c10_rr0 = t1_r13_c10_rr0 + t1_r13_c10_rr1;
  assign t2_r13_c10_rr1 = t1_r13_c10_rr2 + t1_r13_c10_rr3;
  assign t2_r13_c10_rr2 = t1_r13_c10_rr4 + t1_r13_c10_rr5;
  assign t2_r13_c10_rr3 = t1_r13_c10_rr6 + t1_r13_c10_rr7;

  assign t3_r13_c10_rr0 = t2_r13_c10_rr0 + t2_r13_c10_rr1;
  assign t3_r13_c10_rr1 = t2_r13_c10_rr2 + t2_r13_c10_rr3;

  assign t4_r13_c10_rr0 = t3_r13_c10_rr0 + t3_r13_c10_rr1;

  assign c_13_10 = t4_r13_c10_rr0;
  assign t0_r13_c11_rr0 = a_13_0 * b_0_11;
  assign t0_r13_c11_rr1 = a_13_1 * b_1_11;
  assign t0_r13_c11_rr2 = a_13_2 * b_2_11;
  assign t0_r13_c11_rr3 = a_13_3 * b_3_11;
  assign t0_r13_c11_rr4 = a_13_4 * b_4_11;
  assign t0_r13_c11_rr5 = a_13_5 * b_5_11;
  assign t0_r13_c11_rr6 = a_13_6 * b_6_11;
  assign t0_r13_c11_rr7 = a_13_7 * b_7_11;
  assign t0_r13_c11_rr8 = a_13_8 * b_8_11;
  assign t0_r13_c11_rr9 = a_13_9 * b_9_11;
  assign t0_r13_c11_rr10 = a_13_10 * b_10_11;
  assign t0_r13_c11_rr11 = a_13_11 * b_11_11;
  assign t0_r13_c11_rr12 = a_13_12 * b_12_11;
  assign t0_r13_c11_rr13 = a_13_13 * b_13_11;
  assign t0_r13_c11_rr14 = a_13_14 * b_14_11;
  assign t1_r13_c11_rr0 = t0_r13_c11_rr0 + t0_r13_c11_rr1;
  assign t1_r13_c11_rr1 = t0_r13_c11_rr2 + t0_r13_c11_rr3;
  assign t1_r13_c11_rr2 = t0_r13_c11_rr4 + t0_r13_c11_rr5;
  assign t1_r13_c11_rr3 = t0_r13_c11_rr6 + t0_r13_c11_rr7;
  assign t1_r13_c11_rr4 = t0_r13_c11_rr8 + t0_r13_c11_rr9;
  assign t1_r13_c11_rr5 = t0_r13_c11_rr10 + t0_r13_c11_rr11;
  assign t1_r13_c11_rr6 = t0_r13_c11_rr12 + t0_r13_c11_rr13;
  assign t1_r13_c11_rr7 = t0_r13_c11_rr14;

  assign t2_r13_c11_rr0 = t1_r13_c11_rr0 + t1_r13_c11_rr1;
  assign t2_r13_c11_rr1 = t1_r13_c11_rr2 + t1_r13_c11_rr3;
  assign t2_r13_c11_rr2 = t1_r13_c11_rr4 + t1_r13_c11_rr5;
  assign t2_r13_c11_rr3 = t1_r13_c11_rr6 + t1_r13_c11_rr7;

  assign t3_r13_c11_rr0 = t2_r13_c11_rr0 + t2_r13_c11_rr1;
  assign t3_r13_c11_rr1 = t2_r13_c11_rr2 + t2_r13_c11_rr3;

  assign t4_r13_c11_rr0 = t3_r13_c11_rr0 + t3_r13_c11_rr1;

  assign c_13_11 = t4_r13_c11_rr0;
  assign t0_r13_c12_rr0 = a_13_0 * b_0_12;
  assign t0_r13_c12_rr1 = a_13_1 * b_1_12;
  assign t0_r13_c12_rr2 = a_13_2 * b_2_12;
  assign t0_r13_c12_rr3 = a_13_3 * b_3_12;
  assign t0_r13_c12_rr4 = a_13_4 * b_4_12;
  assign t0_r13_c12_rr5 = a_13_5 * b_5_12;
  assign t0_r13_c12_rr6 = a_13_6 * b_6_12;
  assign t0_r13_c12_rr7 = a_13_7 * b_7_12;
  assign t0_r13_c12_rr8 = a_13_8 * b_8_12;
  assign t0_r13_c12_rr9 = a_13_9 * b_9_12;
  assign t0_r13_c12_rr10 = a_13_10 * b_10_12;
  assign t0_r13_c12_rr11 = a_13_11 * b_11_12;
  assign t0_r13_c12_rr12 = a_13_12 * b_12_12;
  assign t0_r13_c12_rr13 = a_13_13 * b_13_12;
  assign t0_r13_c12_rr14 = a_13_14 * b_14_12;
  assign t1_r13_c12_rr0 = t0_r13_c12_rr0 + t0_r13_c12_rr1;
  assign t1_r13_c12_rr1 = t0_r13_c12_rr2 + t0_r13_c12_rr3;
  assign t1_r13_c12_rr2 = t0_r13_c12_rr4 + t0_r13_c12_rr5;
  assign t1_r13_c12_rr3 = t0_r13_c12_rr6 + t0_r13_c12_rr7;
  assign t1_r13_c12_rr4 = t0_r13_c12_rr8 + t0_r13_c12_rr9;
  assign t1_r13_c12_rr5 = t0_r13_c12_rr10 + t0_r13_c12_rr11;
  assign t1_r13_c12_rr6 = t0_r13_c12_rr12 + t0_r13_c12_rr13;
  assign t1_r13_c12_rr7 = t0_r13_c12_rr14;

  assign t2_r13_c12_rr0 = t1_r13_c12_rr0 + t1_r13_c12_rr1;
  assign t2_r13_c12_rr1 = t1_r13_c12_rr2 + t1_r13_c12_rr3;
  assign t2_r13_c12_rr2 = t1_r13_c12_rr4 + t1_r13_c12_rr5;
  assign t2_r13_c12_rr3 = t1_r13_c12_rr6 + t1_r13_c12_rr7;

  assign t3_r13_c12_rr0 = t2_r13_c12_rr0 + t2_r13_c12_rr1;
  assign t3_r13_c12_rr1 = t2_r13_c12_rr2 + t2_r13_c12_rr3;

  assign t4_r13_c12_rr0 = t3_r13_c12_rr0 + t3_r13_c12_rr1;

  assign c_13_12 = t4_r13_c12_rr0;
  assign t0_r13_c13_rr0 = a_13_0 * b_0_13;
  assign t0_r13_c13_rr1 = a_13_1 * b_1_13;
  assign t0_r13_c13_rr2 = a_13_2 * b_2_13;
  assign t0_r13_c13_rr3 = a_13_3 * b_3_13;
  assign t0_r13_c13_rr4 = a_13_4 * b_4_13;
  assign t0_r13_c13_rr5 = a_13_5 * b_5_13;
  assign t0_r13_c13_rr6 = a_13_6 * b_6_13;
  assign t0_r13_c13_rr7 = a_13_7 * b_7_13;
  assign t0_r13_c13_rr8 = a_13_8 * b_8_13;
  assign t0_r13_c13_rr9 = a_13_9 * b_9_13;
  assign t0_r13_c13_rr10 = a_13_10 * b_10_13;
  assign t0_r13_c13_rr11 = a_13_11 * b_11_13;
  assign t0_r13_c13_rr12 = a_13_12 * b_12_13;
  assign t0_r13_c13_rr13 = a_13_13 * b_13_13;
  assign t0_r13_c13_rr14 = a_13_14 * b_14_13;
  assign t1_r13_c13_rr0 = t0_r13_c13_rr0 + t0_r13_c13_rr1;
  assign t1_r13_c13_rr1 = t0_r13_c13_rr2 + t0_r13_c13_rr3;
  assign t1_r13_c13_rr2 = t0_r13_c13_rr4 + t0_r13_c13_rr5;
  assign t1_r13_c13_rr3 = t0_r13_c13_rr6 + t0_r13_c13_rr7;
  assign t1_r13_c13_rr4 = t0_r13_c13_rr8 + t0_r13_c13_rr9;
  assign t1_r13_c13_rr5 = t0_r13_c13_rr10 + t0_r13_c13_rr11;
  assign t1_r13_c13_rr6 = t0_r13_c13_rr12 + t0_r13_c13_rr13;
  assign t1_r13_c13_rr7 = t0_r13_c13_rr14;

  assign t2_r13_c13_rr0 = t1_r13_c13_rr0 + t1_r13_c13_rr1;
  assign t2_r13_c13_rr1 = t1_r13_c13_rr2 + t1_r13_c13_rr3;
  assign t2_r13_c13_rr2 = t1_r13_c13_rr4 + t1_r13_c13_rr5;
  assign t2_r13_c13_rr3 = t1_r13_c13_rr6 + t1_r13_c13_rr7;

  assign t3_r13_c13_rr0 = t2_r13_c13_rr0 + t2_r13_c13_rr1;
  assign t3_r13_c13_rr1 = t2_r13_c13_rr2 + t2_r13_c13_rr3;

  assign t4_r13_c13_rr0 = t3_r13_c13_rr0 + t3_r13_c13_rr1;

  assign c_13_13 = t4_r13_c13_rr0;
  assign t0_r13_c14_rr0 = a_13_0 * b_0_14;
  assign t0_r13_c14_rr1 = a_13_1 * b_1_14;
  assign t0_r13_c14_rr2 = a_13_2 * b_2_14;
  assign t0_r13_c14_rr3 = a_13_3 * b_3_14;
  assign t0_r13_c14_rr4 = a_13_4 * b_4_14;
  assign t0_r13_c14_rr5 = a_13_5 * b_5_14;
  assign t0_r13_c14_rr6 = a_13_6 * b_6_14;
  assign t0_r13_c14_rr7 = a_13_7 * b_7_14;
  assign t0_r13_c14_rr8 = a_13_8 * b_8_14;
  assign t0_r13_c14_rr9 = a_13_9 * b_9_14;
  assign t0_r13_c14_rr10 = a_13_10 * b_10_14;
  assign t0_r13_c14_rr11 = a_13_11 * b_11_14;
  assign t0_r13_c14_rr12 = a_13_12 * b_12_14;
  assign t0_r13_c14_rr13 = a_13_13 * b_13_14;
  assign t0_r13_c14_rr14 = a_13_14 * b_14_14;
  assign t1_r13_c14_rr0 = t0_r13_c14_rr0 + t0_r13_c14_rr1;
  assign t1_r13_c14_rr1 = t0_r13_c14_rr2 + t0_r13_c14_rr3;
  assign t1_r13_c14_rr2 = t0_r13_c14_rr4 + t0_r13_c14_rr5;
  assign t1_r13_c14_rr3 = t0_r13_c14_rr6 + t0_r13_c14_rr7;
  assign t1_r13_c14_rr4 = t0_r13_c14_rr8 + t0_r13_c14_rr9;
  assign t1_r13_c14_rr5 = t0_r13_c14_rr10 + t0_r13_c14_rr11;
  assign t1_r13_c14_rr6 = t0_r13_c14_rr12 + t0_r13_c14_rr13;
  assign t1_r13_c14_rr7 = t0_r13_c14_rr14;

  assign t2_r13_c14_rr0 = t1_r13_c14_rr0 + t1_r13_c14_rr1;
  assign t2_r13_c14_rr1 = t1_r13_c14_rr2 + t1_r13_c14_rr3;
  assign t2_r13_c14_rr2 = t1_r13_c14_rr4 + t1_r13_c14_rr5;
  assign t2_r13_c14_rr3 = t1_r13_c14_rr6 + t1_r13_c14_rr7;

  assign t3_r13_c14_rr0 = t2_r13_c14_rr0 + t2_r13_c14_rr1;
  assign t3_r13_c14_rr1 = t2_r13_c14_rr2 + t2_r13_c14_rr3;

  assign t4_r13_c14_rr0 = t3_r13_c14_rr0 + t3_r13_c14_rr1;

  assign c_13_14 = t4_r13_c14_rr0;
  assign t0_r14_c0_rr0 = a_14_0 * b_0_0;
  assign t0_r14_c0_rr1 = a_14_1 * b_1_0;
  assign t0_r14_c0_rr2 = a_14_2 * b_2_0;
  assign t0_r14_c0_rr3 = a_14_3 * b_3_0;
  assign t0_r14_c0_rr4 = a_14_4 * b_4_0;
  assign t0_r14_c0_rr5 = a_14_5 * b_5_0;
  assign t0_r14_c0_rr6 = a_14_6 * b_6_0;
  assign t0_r14_c0_rr7 = a_14_7 * b_7_0;
  assign t0_r14_c0_rr8 = a_14_8 * b_8_0;
  assign t0_r14_c0_rr9 = a_14_9 * b_9_0;
  assign t0_r14_c0_rr10 = a_14_10 * b_10_0;
  assign t0_r14_c0_rr11 = a_14_11 * b_11_0;
  assign t0_r14_c0_rr12 = a_14_12 * b_12_0;
  assign t0_r14_c0_rr13 = a_14_13 * b_13_0;
  assign t0_r14_c0_rr14 = a_14_14 * b_14_0;
  assign t1_r14_c0_rr0 = t0_r14_c0_rr0 + t0_r14_c0_rr1;
  assign t1_r14_c0_rr1 = t0_r14_c0_rr2 + t0_r14_c0_rr3;
  assign t1_r14_c0_rr2 = t0_r14_c0_rr4 + t0_r14_c0_rr5;
  assign t1_r14_c0_rr3 = t0_r14_c0_rr6 + t0_r14_c0_rr7;
  assign t1_r14_c0_rr4 = t0_r14_c0_rr8 + t0_r14_c0_rr9;
  assign t1_r14_c0_rr5 = t0_r14_c0_rr10 + t0_r14_c0_rr11;
  assign t1_r14_c0_rr6 = t0_r14_c0_rr12 + t0_r14_c0_rr13;
  assign t1_r14_c0_rr7 = t0_r14_c0_rr14;

  assign t2_r14_c0_rr0 = t1_r14_c0_rr0 + t1_r14_c0_rr1;
  assign t2_r14_c0_rr1 = t1_r14_c0_rr2 + t1_r14_c0_rr3;
  assign t2_r14_c0_rr2 = t1_r14_c0_rr4 + t1_r14_c0_rr5;
  assign t2_r14_c0_rr3 = t1_r14_c0_rr6 + t1_r14_c0_rr7;

  assign t3_r14_c0_rr0 = t2_r14_c0_rr0 + t2_r14_c0_rr1;
  assign t3_r14_c0_rr1 = t2_r14_c0_rr2 + t2_r14_c0_rr3;

  assign t4_r14_c0_rr0 = t3_r14_c0_rr0 + t3_r14_c0_rr1;

  assign c_14_0 = t4_r14_c0_rr0;
  assign t0_r14_c1_rr0 = a_14_0 * b_0_1;
  assign t0_r14_c1_rr1 = a_14_1 * b_1_1;
  assign t0_r14_c1_rr2 = a_14_2 * b_2_1;
  assign t0_r14_c1_rr3 = a_14_3 * b_3_1;
  assign t0_r14_c1_rr4 = a_14_4 * b_4_1;
  assign t0_r14_c1_rr5 = a_14_5 * b_5_1;
  assign t0_r14_c1_rr6 = a_14_6 * b_6_1;
  assign t0_r14_c1_rr7 = a_14_7 * b_7_1;
  assign t0_r14_c1_rr8 = a_14_8 * b_8_1;
  assign t0_r14_c1_rr9 = a_14_9 * b_9_1;
  assign t0_r14_c1_rr10 = a_14_10 * b_10_1;
  assign t0_r14_c1_rr11 = a_14_11 * b_11_1;
  assign t0_r14_c1_rr12 = a_14_12 * b_12_1;
  assign t0_r14_c1_rr13 = a_14_13 * b_13_1;
  assign t0_r14_c1_rr14 = a_14_14 * b_14_1;
  assign t1_r14_c1_rr0 = t0_r14_c1_rr0 + t0_r14_c1_rr1;
  assign t1_r14_c1_rr1 = t0_r14_c1_rr2 + t0_r14_c1_rr3;
  assign t1_r14_c1_rr2 = t0_r14_c1_rr4 + t0_r14_c1_rr5;
  assign t1_r14_c1_rr3 = t0_r14_c1_rr6 + t0_r14_c1_rr7;
  assign t1_r14_c1_rr4 = t0_r14_c1_rr8 + t0_r14_c1_rr9;
  assign t1_r14_c1_rr5 = t0_r14_c1_rr10 + t0_r14_c1_rr11;
  assign t1_r14_c1_rr6 = t0_r14_c1_rr12 + t0_r14_c1_rr13;
  assign t1_r14_c1_rr7 = t0_r14_c1_rr14;

  assign t2_r14_c1_rr0 = t1_r14_c1_rr0 + t1_r14_c1_rr1;
  assign t2_r14_c1_rr1 = t1_r14_c1_rr2 + t1_r14_c1_rr3;
  assign t2_r14_c1_rr2 = t1_r14_c1_rr4 + t1_r14_c1_rr5;
  assign t2_r14_c1_rr3 = t1_r14_c1_rr6 + t1_r14_c1_rr7;

  assign t3_r14_c1_rr0 = t2_r14_c1_rr0 + t2_r14_c1_rr1;
  assign t3_r14_c1_rr1 = t2_r14_c1_rr2 + t2_r14_c1_rr3;

  assign t4_r14_c1_rr0 = t3_r14_c1_rr0 + t3_r14_c1_rr1;

  assign c_14_1 = t4_r14_c1_rr0;
  assign t0_r14_c2_rr0 = a_14_0 * b_0_2;
  assign t0_r14_c2_rr1 = a_14_1 * b_1_2;
  assign t0_r14_c2_rr2 = a_14_2 * b_2_2;
  assign t0_r14_c2_rr3 = a_14_3 * b_3_2;
  assign t0_r14_c2_rr4 = a_14_4 * b_4_2;
  assign t0_r14_c2_rr5 = a_14_5 * b_5_2;
  assign t0_r14_c2_rr6 = a_14_6 * b_6_2;
  assign t0_r14_c2_rr7 = a_14_7 * b_7_2;
  assign t0_r14_c2_rr8 = a_14_8 * b_8_2;
  assign t0_r14_c2_rr9 = a_14_9 * b_9_2;
  assign t0_r14_c2_rr10 = a_14_10 * b_10_2;
  assign t0_r14_c2_rr11 = a_14_11 * b_11_2;
  assign t0_r14_c2_rr12 = a_14_12 * b_12_2;
  assign t0_r14_c2_rr13 = a_14_13 * b_13_2;
  assign t0_r14_c2_rr14 = a_14_14 * b_14_2;
  assign t1_r14_c2_rr0 = t0_r14_c2_rr0 + t0_r14_c2_rr1;
  assign t1_r14_c2_rr1 = t0_r14_c2_rr2 + t0_r14_c2_rr3;
  assign t1_r14_c2_rr2 = t0_r14_c2_rr4 + t0_r14_c2_rr5;
  assign t1_r14_c2_rr3 = t0_r14_c2_rr6 + t0_r14_c2_rr7;
  assign t1_r14_c2_rr4 = t0_r14_c2_rr8 + t0_r14_c2_rr9;
  assign t1_r14_c2_rr5 = t0_r14_c2_rr10 + t0_r14_c2_rr11;
  assign t1_r14_c2_rr6 = t0_r14_c2_rr12 + t0_r14_c2_rr13;
  assign t1_r14_c2_rr7 = t0_r14_c2_rr14;

  assign t2_r14_c2_rr0 = t1_r14_c2_rr0 + t1_r14_c2_rr1;
  assign t2_r14_c2_rr1 = t1_r14_c2_rr2 + t1_r14_c2_rr3;
  assign t2_r14_c2_rr2 = t1_r14_c2_rr4 + t1_r14_c2_rr5;
  assign t2_r14_c2_rr3 = t1_r14_c2_rr6 + t1_r14_c2_rr7;

  assign t3_r14_c2_rr0 = t2_r14_c2_rr0 + t2_r14_c2_rr1;
  assign t3_r14_c2_rr1 = t2_r14_c2_rr2 + t2_r14_c2_rr3;

  assign t4_r14_c2_rr0 = t3_r14_c2_rr0 + t3_r14_c2_rr1;

  assign c_14_2 = t4_r14_c2_rr0;
  assign t0_r14_c3_rr0 = a_14_0 * b_0_3;
  assign t0_r14_c3_rr1 = a_14_1 * b_1_3;
  assign t0_r14_c3_rr2 = a_14_2 * b_2_3;
  assign t0_r14_c3_rr3 = a_14_3 * b_3_3;
  assign t0_r14_c3_rr4 = a_14_4 * b_4_3;
  assign t0_r14_c3_rr5 = a_14_5 * b_5_3;
  assign t0_r14_c3_rr6 = a_14_6 * b_6_3;
  assign t0_r14_c3_rr7 = a_14_7 * b_7_3;
  assign t0_r14_c3_rr8 = a_14_8 * b_8_3;
  assign t0_r14_c3_rr9 = a_14_9 * b_9_3;
  assign t0_r14_c3_rr10 = a_14_10 * b_10_3;
  assign t0_r14_c3_rr11 = a_14_11 * b_11_3;
  assign t0_r14_c3_rr12 = a_14_12 * b_12_3;
  assign t0_r14_c3_rr13 = a_14_13 * b_13_3;
  assign t0_r14_c3_rr14 = a_14_14 * b_14_3;
  assign t1_r14_c3_rr0 = t0_r14_c3_rr0 + t0_r14_c3_rr1;
  assign t1_r14_c3_rr1 = t0_r14_c3_rr2 + t0_r14_c3_rr3;
  assign t1_r14_c3_rr2 = t0_r14_c3_rr4 + t0_r14_c3_rr5;
  assign t1_r14_c3_rr3 = t0_r14_c3_rr6 + t0_r14_c3_rr7;
  assign t1_r14_c3_rr4 = t0_r14_c3_rr8 + t0_r14_c3_rr9;
  assign t1_r14_c3_rr5 = t0_r14_c3_rr10 + t0_r14_c3_rr11;
  assign t1_r14_c3_rr6 = t0_r14_c3_rr12 + t0_r14_c3_rr13;
  assign t1_r14_c3_rr7 = t0_r14_c3_rr14;

  assign t2_r14_c3_rr0 = t1_r14_c3_rr0 + t1_r14_c3_rr1;
  assign t2_r14_c3_rr1 = t1_r14_c3_rr2 + t1_r14_c3_rr3;
  assign t2_r14_c3_rr2 = t1_r14_c3_rr4 + t1_r14_c3_rr5;
  assign t2_r14_c3_rr3 = t1_r14_c3_rr6 + t1_r14_c3_rr7;

  assign t3_r14_c3_rr0 = t2_r14_c3_rr0 + t2_r14_c3_rr1;
  assign t3_r14_c3_rr1 = t2_r14_c3_rr2 + t2_r14_c3_rr3;

  assign t4_r14_c3_rr0 = t3_r14_c3_rr0 + t3_r14_c3_rr1;

  assign c_14_3 = t4_r14_c3_rr0;
  assign t0_r14_c4_rr0 = a_14_0 * b_0_4;
  assign t0_r14_c4_rr1 = a_14_1 * b_1_4;
  assign t0_r14_c4_rr2 = a_14_2 * b_2_4;
  assign t0_r14_c4_rr3 = a_14_3 * b_3_4;
  assign t0_r14_c4_rr4 = a_14_4 * b_4_4;
  assign t0_r14_c4_rr5 = a_14_5 * b_5_4;
  assign t0_r14_c4_rr6 = a_14_6 * b_6_4;
  assign t0_r14_c4_rr7 = a_14_7 * b_7_4;
  assign t0_r14_c4_rr8 = a_14_8 * b_8_4;
  assign t0_r14_c4_rr9 = a_14_9 * b_9_4;
  assign t0_r14_c4_rr10 = a_14_10 * b_10_4;
  assign t0_r14_c4_rr11 = a_14_11 * b_11_4;
  assign t0_r14_c4_rr12 = a_14_12 * b_12_4;
  assign t0_r14_c4_rr13 = a_14_13 * b_13_4;
  assign t0_r14_c4_rr14 = a_14_14 * b_14_4;
  assign t1_r14_c4_rr0 = t0_r14_c4_rr0 + t0_r14_c4_rr1;
  assign t1_r14_c4_rr1 = t0_r14_c4_rr2 + t0_r14_c4_rr3;
  assign t1_r14_c4_rr2 = t0_r14_c4_rr4 + t0_r14_c4_rr5;
  assign t1_r14_c4_rr3 = t0_r14_c4_rr6 + t0_r14_c4_rr7;
  assign t1_r14_c4_rr4 = t0_r14_c4_rr8 + t0_r14_c4_rr9;
  assign t1_r14_c4_rr5 = t0_r14_c4_rr10 + t0_r14_c4_rr11;
  assign t1_r14_c4_rr6 = t0_r14_c4_rr12 + t0_r14_c4_rr13;
  assign t1_r14_c4_rr7 = t0_r14_c4_rr14;

  assign t2_r14_c4_rr0 = t1_r14_c4_rr0 + t1_r14_c4_rr1;
  assign t2_r14_c4_rr1 = t1_r14_c4_rr2 + t1_r14_c4_rr3;
  assign t2_r14_c4_rr2 = t1_r14_c4_rr4 + t1_r14_c4_rr5;
  assign t2_r14_c4_rr3 = t1_r14_c4_rr6 + t1_r14_c4_rr7;

  assign t3_r14_c4_rr0 = t2_r14_c4_rr0 + t2_r14_c4_rr1;
  assign t3_r14_c4_rr1 = t2_r14_c4_rr2 + t2_r14_c4_rr3;

  assign t4_r14_c4_rr0 = t3_r14_c4_rr0 + t3_r14_c4_rr1;

  assign c_14_4 = t4_r14_c4_rr0;
  assign t0_r14_c5_rr0 = a_14_0 * b_0_5;
  assign t0_r14_c5_rr1 = a_14_1 * b_1_5;
  assign t0_r14_c5_rr2 = a_14_2 * b_2_5;
  assign t0_r14_c5_rr3 = a_14_3 * b_3_5;
  assign t0_r14_c5_rr4 = a_14_4 * b_4_5;
  assign t0_r14_c5_rr5 = a_14_5 * b_5_5;
  assign t0_r14_c5_rr6 = a_14_6 * b_6_5;
  assign t0_r14_c5_rr7 = a_14_7 * b_7_5;
  assign t0_r14_c5_rr8 = a_14_8 * b_8_5;
  assign t0_r14_c5_rr9 = a_14_9 * b_9_5;
  assign t0_r14_c5_rr10 = a_14_10 * b_10_5;
  assign t0_r14_c5_rr11 = a_14_11 * b_11_5;
  assign t0_r14_c5_rr12 = a_14_12 * b_12_5;
  assign t0_r14_c5_rr13 = a_14_13 * b_13_5;
  assign t0_r14_c5_rr14 = a_14_14 * b_14_5;
  assign t1_r14_c5_rr0 = t0_r14_c5_rr0 + t0_r14_c5_rr1;
  assign t1_r14_c5_rr1 = t0_r14_c5_rr2 + t0_r14_c5_rr3;
  assign t1_r14_c5_rr2 = t0_r14_c5_rr4 + t0_r14_c5_rr5;
  assign t1_r14_c5_rr3 = t0_r14_c5_rr6 + t0_r14_c5_rr7;
  assign t1_r14_c5_rr4 = t0_r14_c5_rr8 + t0_r14_c5_rr9;
  assign t1_r14_c5_rr5 = t0_r14_c5_rr10 + t0_r14_c5_rr11;
  assign t1_r14_c5_rr6 = t0_r14_c5_rr12 + t0_r14_c5_rr13;
  assign t1_r14_c5_rr7 = t0_r14_c5_rr14;

  assign t2_r14_c5_rr0 = t1_r14_c5_rr0 + t1_r14_c5_rr1;
  assign t2_r14_c5_rr1 = t1_r14_c5_rr2 + t1_r14_c5_rr3;
  assign t2_r14_c5_rr2 = t1_r14_c5_rr4 + t1_r14_c5_rr5;
  assign t2_r14_c5_rr3 = t1_r14_c5_rr6 + t1_r14_c5_rr7;

  assign t3_r14_c5_rr0 = t2_r14_c5_rr0 + t2_r14_c5_rr1;
  assign t3_r14_c5_rr1 = t2_r14_c5_rr2 + t2_r14_c5_rr3;

  assign t4_r14_c5_rr0 = t3_r14_c5_rr0 + t3_r14_c5_rr1;

  assign c_14_5 = t4_r14_c5_rr0;
  assign t0_r14_c6_rr0 = a_14_0 * b_0_6;
  assign t0_r14_c6_rr1 = a_14_1 * b_1_6;
  assign t0_r14_c6_rr2 = a_14_2 * b_2_6;
  assign t0_r14_c6_rr3 = a_14_3 * b_3_6;
  assign t0_r14_c6_rr4 = a_14_4 * b_4_6;
  assign t0_r14_c6_rr5 = a_14_5 * b_5_6;
  assign t0_r14_c6_rr6 = a_14_6 * b_6_6;
  assign t0_r14_c6_rr7 = a_14_7 * b_7_6;
  assign t0_r14_c6_rr8 = a_14_8 * b_8_6;
  assign t0_r14_c6_rr9 = a_14_9 * b_9_6;
  assign t0_r14_c6_rr10 = a_14_10 * b_10_6;
  assign t0_r14_c6_rr11 = a_14_11 * b_11_6;
  assign t0_r14_c6_rr12 = a_14_12 * b_12_6;
  assign t0_r14_c6_rr13 = a_14_13 * b_13_6;
  assign t0_r14_c6_rr14 = a_14_14 * b_14_6;
  assign t1_r14_c6_rr0 = t0_r14_c6_rr0 + t0_r14_c6_rr1;
  assign t1_r14_c6_rr1 = t0_r14_c6_rr2 + t0_r14_c6_rr3;
  assign t1_r14_c6_rr2 = t0_r14_c6_rr4 + t0_r14_c6_rr5;
  assign t1_r14_c6_rr3 = t0_r14_c6_rr6 + t0_r14_c6_rr7;
  assign t1_r14_c6_rr4 = t0_r14_c6_rr8 + t0_r14_c6_rr9;
  assign t1_r14_c6_rr5 = t0_r14_c6_rr10 + t0_r14_c6_rr11;
  assign t1_r14_c6_rr6 = t0_r14_c6_rr12 + t0_r14_c6_rr13;
  assign t1_r14_c6_rr7 = t0_r14_c6_rr14;

  assign t2_r14_c6_rr0 = t1_r14_c6_rr0 + t1_r14_c6_rr1;
  assign t2_r14_c6_rr1 = t1_r14_c6_rr2 + t1_r14_c6_rr3;
  assign t2_r14_c6_rr2 = t1_r14_c6_rr4 + t1_r14_c6_rr5;
  assign t2_r14_c6_rr3 = t1_r14_c6_rr6 + t1_r14_c6_rr7;

  assign t3_r14_c6_rr0 = t2_r14_c6_rr0 + t2_r14_c6_rr1;
  assign t3_r14_c6_rr1 = t2_r14_c6_rr2 + t2_r14_c6_rr3;

  assign t4_r14_c6_rr0 = t3_r14_c6_rr0 + t3_r14_c6_rr1;

  assign c_14_6 = t4_r14_c6_rr0;
  assign t0_r14_c7_rr0 = a_14_0 * b_0_7;
  assign t0_r14_c7_rr1 = a_14_1 * b_1_7;
  assign t0_r14_c7_rr2 = a_14_2 * b_2_7;
  assign t0_r14_c7_rr3 = a_14_3 * b_3_7;
  assign t0_r14_c7_rr4 = a_14_4 * b_4_7;
  assign t0_r14_c7_rr5 = a_14_5 * b_5_7;
  assign t0_r14_c7_rr6 = a_14_6 * b_6_7;
  assign t0_r14_c7_rr7 = a_14_7 * b_7_7;
  assign t0_r14_c7_rr8 = a_14_8 * b_8_7;
  assign t0_r14_c7_rr9 = a_14_9 * b_9_7;
  assign t0_r14_c7_rr10 = a_14_10 * b_10_7;
  assign t0_r14_c7_rr11 = a_14_11 * b_11_7;
  assign t0_r14_c7_rr12 = a_14_12 * b_12_7;
  assign t0_r14_c7_rr13 = a_14_13 * b_13_7;
  assign t0_r14_c7_rr14 = a_14_14 * b_14_7;
  assign t1_r14_c7_rr0 = t0_r14_c7_rr0 + t0_r14_c7_rr1;
  assign t1_r14_c7_rr1 = t0_r14_c7_rr2 + t0_r14_c7_rr3;
  assign t1_r14_c7_rr2 = t0_r14_c7_rr4 + t0_r14_c7_rr5;
  assign t1_r14_c7_rr3 = t0_r14_c7_rr6 + t0_r14_c7_rr7;
  assign t1_r14_c7_rr4 = t0_r14_c7_rr8 + t0_r14_c7_rr9;
  assign t1_r14_c7_rr5 = t0_r14_c7_rr10 + t0_r14_c7_rr11;
  assign t1_r14_c7_rr6 = t0_r14_c7_rr12 + t0_r14_c7_rr13;
  assign t1_r14_c7_rr7 = t0_r14_c7_rr14;

  assign t2_r14_c7_rr0 = t1_r14_c7_rr0 + t1_r14_c7_rr1;
  assign t2_r14_c7_rr1 = t1_r14_c7_rr2 + t1_r14_c7_rr3;
  assign t2_r14_c7_rr2 = t1_r14_c7_rr4 + t1_r14_c7_rr5;
  assign t2_r14_c7_rr3 = t1_r14_c7_rr6 + t1_r14_c7_rr7;

  assign t3_r14_c7_rr0 = t2_r14_c7_rr0 + t2_r14_c7_rr1;
  assign t3_r14_c7_rr1 = t2_r14_c7_rr2 + t2_r14_c7_rr3;

  assign t4_r14_c7_rr0 = t3_r14_c7_rr0 + t3_r14_c7_rr1;

  assign c_14_7 = t4_r14_c7_rr0;
  assign t0_r14_c8_rr0 = a_14_0 * b_0_8;
  assign t0_r14_c8_rr1 = a_14_1 * b_1_8;
  assign t0_r14_c8_rr2 = a_14_2 * b_2_8;
  assign t0_r14_c8_rr3 = a_14_3 * b_3_8;
  assign t0_r14_c8_rr4 = a_14_4 * b_4_8;
  assign t0_r14_c8_rr5 = a_14_5 * b_5_8;
  assign t0_r14_c8_rr6 = a_14_6 * b_6_8;
  assign t0_r14_c8_rr7 = a_14_7 * b_7_8;
  assign t0_r14_c8_rr8 = a_14_8 * b_8_8;
  assign t0_r14_c8_rr9 = a_14_9 * b_9_8;
  assign t0_r14_c8_rr10 = a_14_10 * b_10_8;
  assign t0_r14_c8_rr11 = a_14_11 * b_11_8;
  assign t0_r14_c8_rr12 = a_14_12 * b_12_8;
  assign t0_r14_c8_rr13 = a_14_13 * b_13_8;
  assign t0_r14_c8_rr14 = a_14_14 * b_14_8;
  assign t1_r14_c8_rr0 = t0_r14_c8_rr0 + t0_r14_c8_rr1;
  assign t1_r14_c8_rr1 = t0_r14_c8_rr2 + t0_r14_c8_rr3;
  assign t1_r14_c8_rr2 = t0_r14_c8_rr4 + t0_r14_c8_rr5;
  assign t1_r14_c8_rr3 = t0_r14_c8_rr6 + t0_r14_c8_rr7;
  assign t1_r14_c8_rr4 = t0_r14_c8_rr8 + t0_r14_c8_rr9;
  assign t1_r14_c8_rr5 = t0_r14_c8_rr10 + t0_r14_c8_rr11;
  assign t1_r14_c8_rr6 = t0_r14_c8_rr12 + t0_r14_c8_rr13;
  assign t1_r14_c8_rr7 = t0_r14_c8_rr14;

  assign t2_r14_c8_rr0 = t1_r14_c8_rr0 + t1_r14_c8_rr1;
  assign t2_r14_c8_rr1 = t1_r14_c8_rr2 + t1_r14_c8_rr3;
  assign t2_r14_c8_rr2 = t1_r14_c8_rr4 + t1_r14_c8_rr5;
  assign t2_r14_c8_rr3 = t1_r14_c8_rr6 + t1_r14_c8_rr7;

  assign t3_r14_c8_rr0 = t2_r14_c8_rr0 + t2_r14_c8_rr1;
  assign t3_r14_c8_rr1 = t2_r14_c8_rr2 + t2_r14_c8_rr3;

  assign t4_r14_c8_rr0 = t3_r14_c8_rr0 + t3_r14_c8_rr1;

  assign c_14_8 = t4_r14_c8_rr0;
  assign t0_r14_c9_rr0 = a_14_0 * b_0_9;
  assign t0_r14_c9_rr1 = a_14_1 * b_1_9;
  assign t0_r14_c9_rr2 = a_14_2 * b_2_9;
  assign t0_r14_c9_rr3 = a_14_3 * b_3_9;
  assign t0_r14_c9_rr4 = a_14_4 * b_4_9;
  assign t0_r14_c9_rr5 = a_14_5 * b_5_9;
  assign t0_r14_c9_rr6 = a_14_6 * b_6_9;
  assign t0_r14_c9_rr7 = a_14_7 * b_7_9;
  assign t0_r14_c9_rr8 = a_14_8 * b_8_9;
  assign t0_r14_c9_rr9 = a_14_9 * b_9_9;
  assign t0_r14_c9_rr10 = a_14_10 * b_10_9;
  assign t0_r14_c9_rr11 = a_14_11 * b_11_9;
  assign t0_r14_c9_rr12 = a_14_12 * b_12_9;
  assign t0_r14_c9_rr13 = a_14_13 * b_13_9;
  assign t0_r14_c9_rr14 = a_14_14 * b_14_9;
  assign t1_r14_c9_rr0 = t0_r14_c9_rr0 + t0_r14_c9_rr1;
  assign t1_r14_c9_rr1 = t0_r14_c9_rr2 + t0_r14_c9_rr3;
  assign t1_r14_c9_rr2 = t0_r14_c9_rr4 + t0_r14_c9_rr5;
  assign t1_r14_c9_rr3 = t0_r14_c9_rr6 + t0_r14_c9_rr7;
  assign t1_r14_c9_rr4 = t0_r14_c9_rr8 + t0_r14_c9_rr9;
  assign t1_r14_c9_rr5 = t0_r14_c9_rr10 + t0_r14_c9_rr11;
  assign t1_r14_c9_rr6 = t0_r14_c9_rr12 + t0_r14_c9_rr13;
  assign t1_r14_c9_rr7 = t0_r14_c9_rr14;

  assign t2_r14_c9_rr0 = t1_r14_c9_rr0 + t1_r14_c9_rr1;
  assign t2_r14_c9_rr1 = t1_r14_c9_rr2 + t1_r14_c9_rr3;
  assign t2_r14_c9_rr2 = t1_r14_c9_rr4 + t1_r14_c9_rr5;
  assign t2_r14_c9_rr3 = t1_r14_c9_rr6 + t1_r14_c9_rr7;

  assign t3_r14_c9_rr0 = t2_r14_c9_rr0 + t2_r14_c9_rr1;
  assign t3_r14_c9_rr1 = t2_r14_c9_rr2 + t2_r14_c9_rr3;

  assign t4_r14_c9_rr0 = t3_r14_c9_rr0 + t3_r14_c9_rr1;

  assign c_14_9 = t4_r14_c9_rr0;
  assign t0_r14_c10_rr0 = a_14_0 * b_0_10;
  assign t0_r14_c10_rr1 = a_14_1 * b_1_10;
  assign t0_r14_c10_rr2 = a_14_2 * b_2_10;
  assign t0_r14_c10_rr3 = a_14_3 * b_3_10;
  assign t0_r14_c10_rr4 = a_14_4 * b_4_10;
  assign t0_r14_c10_rr5 = a_14_5 * b_5_10;
  assign t0_r14_c10_rr6 = a_14_6 * b_6_10;
  assign t0_r14_c10_rr7 = a_14_7 * b_7_10;
  assign t0_r14_c10_rr8 = a_14_8 * b_8_10;
  assign t0_r14_c10_rr9 = a_14_9 * b_9_10;
  assign t0_r14_c10_rr10 = a_14_10 * b_10_10;
  assign t0_r14_c10_rr11 = a_14_11 * b_11_10;
  assign t0_r14_c10_rr12 = a_14_12 * b_12_10;
  assign t0_r14_c10_rr13 = a_14_13 * b_13_10;
  assign t0_r14_c10_rr14 = a_14_14 * b_14_10;
  assign t1_r14_c10_rr0 = t0_r14_c10_rr0 + t0_r14_c10_rr1;
  assign t1_r14_c10_rr1 = t0_r14_c10_rr2 + t0_r14_c10_rr3;
  assign t1_r14_c10_rr2 = t0_r14_c10_rr4 + t0_r14_c10_rr5;
  assign t1_r14_c10_rr3 = t0_r14_c10_rr6 + t0_r14_c10_rr7;
  assign t1_r14_c10_rr4 = t0_r14_c10_rr8 + t0_r14_c10_rr9;
  assign t1_r14_c10_rr5 = t0_r14_c10_rr10 + t0_r14_c10_rr11;
  assign t1_r14_c10_rr6 = t0_r14_c10_rr12 + t0_r14_c10_rr13;
  assign t1_r14_c10_rr7 = t0_r14_c10_rr14;

  assign t2_r14_c10_rr0 = t1_r14_c10_rr0 + t1_r14_c10_rr1;
  assign t2_r14_c10_rr1 = t1_r14_c10_rr2 + t1_r14_c10_rr3;
  assign t2_r14_c10_rr2 = t1_r14_c10_rr4 + t1_r14_c10_rr5;
  assign t2_r14_c10_rr3 = t1_r14_c10_rr6 + t1_r14_c10_rr7;

  assign t3_r14_c10_rr0 = t2_r14_c10_rr0 + t2_r14_c10_rr1;
  assign t3_r14_c10_rr1 = t2_r14_c10_rr2 + t2_r14_c10_rr3;

  assign t4_r14_c10_rr0 = t3_r14_c10_rr0 + t3_r14_c10_rr1;

  assign c_14_10 = t4_r14_c10_rr0;
  assign t0_r14_c11_rr0 = a_14_0 * b_0_11;
  assign t0_r14_c11_rr1 = a_14_1 * b_1_11;
  assign t0_r14_c11_rr2 = a_14_2 * b_2_11;
  assign t0_r14_c11_rr3 = a_14_3 * b_3_11;
  assign t0_r14_c11_rr4 = a_14_4 * b_4_11;
  assign t0_r14_c11_rr5 = a_14_5 * b_5_11;
  assign t0_r14_c11_rr6 = a_14_6 * b_6_11;
  assign t0_r14_c11_rr7 = a_14_7 * b_7_11;
  assign t0_r14_c11_rr8 = a_14_8 * b_8_11;
  assign t0_r14_c11_rr9 = a_14_9 * b_9_11;
  assign t0_r14_c11_rr10 = a_14_10 * b_10_11;
  assign t0_r14_c11_rr11 = a_14_11 * b_11_11;
  assign t0_r14_c11_rr12 = a_14_12 * b_12_11;
  assign t0_r14_c11_rr13 = a_14_13 * b_13_11;
  assign t0_r14_c11_rr14 = a_14_14 * b_14_11;
  assign t1_r14_c11_rr0 = t0_r14_c11_rr0 + t0_r14_c11_rr1;
  assign t1_r14_c11_rr1 = t0_r14_c11_rr2 + t0_r14_c11_rr3;
  assign t1_r14_c11_rr2 = t0_r14_c11_rr4 + t0_r14_c11_rr5;
  assign t1_r14_c11_rr3 = t0_r14_c11_rr6 + t0_r14_c11_rr7;
  assign t1_r14_c11_rr4 = t0_r14_c11_rr8 + t0_r14_c11_rr9;
  assign t1_r14_c11_rr5 = t0_r14_c11_rr10 + t0_r14_c11_rr11;
  assign t1_r14_c11_rr6 = t0_r14_c11_rr12 + t0_r14_c11_rr13;
  assign t1_r14_c11_rr7 = t0_r14_c11_rr14;

  assign t2_r14_c11_rr0 = t1_r14_c11_rr0 + t1_r14_c11_rr1;
  assign t2_r14_c11_rr1 = t1_r14_c11_rr2 + t1_r14_c11_rr3;
  assign t2_r14_c11_rr2 = t1_r14_c11_rr4 + t1_r14_c11_rr5;
  assign t2_r14_c11_rr3 = t1_r14_c11_rr6 + t1_r14_c11_rr7;

  assign t3_r14_c11_rr0 = t2_r14_c11_rr0 + t2_r14_c11_rr1;
  assign t3_r14_c11_rr1 = t2_r14_c11_rr2 + t2_r14_c11_rr3;

  assign t4_r14_c11_rr0 = t3_r14_c11_rr0 + t3_r14_c11_rr1;

  assign c_14_11 = t4_r14_c11_rr0;
  assign t0_r14_c12_rr0 = a_14_0 * b_0_12;
  assign t0_r14_c12_rr1 = a_14_1 * b_1_12;
  assign t0_r14_c12_rr2 = a_14_2 * b_2_12;
  assign t0_r14_c12_rr3 = a_14_3 * b_3_12;
  assign t0_r14_c12_rr4 = a_14_4 * b_4_12;
  assign t0_r14_c12_rr5 = a_14_5 * b_5_12;
  assign t0_r14_c12_rr6 = a_14_6 * b_6_12;
  assign t0_r14_c12_rr7 = a_14_7 * b_7_12;
  assign t0_r14_c12_rr8 = a_14_8 * b_8_12;
  assign t0_r14_c12_rr9 = a_14_9 * b_9_12;
  assign t0_r14_c12_rr10 = a_14_10 * b_10_12;
  assign t0_r14_c12_rr11 = a_14_11 * b_11_12;
  assign t0_r14_c12_rr12 = a_14_12 * b_12_12;
  assign t0_r14_c12_rr13 = a_14_13 * b_13_12;
  assign t0_r14_c12_rr14 = a_14_14 * b_14_12;
  assign t1_r14_c12_rr0 = t0_r14_c12_rr0 + t0_r14_c12_rr1;
  assign t1_r14_c12_rr1 = t0_r14_c12_rr2 + t0_r14_c12_rr3;
  assign t1_r14_c12_rr2 = t0_r14_c12_rr4 + t0_r14_c12_rr5;
  assign t1_r14_c12_rr3 = t0_r14_c12_rr6 + t0_r14_c12_rr7;
  assign t1_r14_c12_rr4 = t0_r14_c12_rr8 + t0_r14_c12_rr9;
  assign t1_r14_c12_rr5 = t0_r14_c12_rr10 + t0_r14_c12_rr11;
  assign t1_r14_c12_rr6 = t0_r14_c12_rr12 + t0_r14_c12_rr13;
  assign t1_r14_c12_rr7 = t0_r14_c12_rr14;

  assign t2_r14_c12_rr0 = t1_r14_c12_rr0 + t1_r14_c12_rr1;
  assign t2_r14_c12_rr1 = t1_r14_c12_rr2 + t1_r14_c12_rr3;
  assign t2_r14_c12_rr2 = t1_r14_c12_rr4 + t1_r14_c12_rr5;
  assign t2_r14_c12_rr3 = t1_r14_c12_rr6 + t1_r14_c12_rr7;

  assign t3_r14_c12_rr0 = t2_r14_c12_rr0 + t2_r14_c12_rr1;
  assign t3_r14_c12_rr1 = t2_r14_c12_rr2 + t2_r14_c12_rr3;

  assign t4_r14_c12_rr0 = t3_r14_c12_rr0 + t3_r14_c12_rr1;

  assign c_14_12 = t4_r14_c12_rr0;
  assign t0_r14_c13_rr0 = a_14_0 * b_0_13;
  assign t0_r14_c13_rr1 = a_14_1 * b_1_13;
  assign t0_r14_c13_rr2 = a_14_2 * b_2_13;
  assign t0_r14_c13_rr3 = a_14_3 * b_3_13;
  assign t0_r14_c13_rr4 = a_14_4 * b_4_13;
  assign t0_r14_c13_rr5 = a_14_5 * b_5_13;
  assign t0_r14_c13_rr6 = a_14_6 * b_6_13;
  assign t0_r14_c13_rr7 = a_14_7 * b_7_13;
  assign t0_r14_c13_rr8 = a_14_8 * b_8_13;
  assign t0_r14_c13_rr9 = a_14_9 * b_9_13;
  assign t0_r14_c13_rr10 = a_14_10 * b_10_13;
  assign t0_r14_c13_rr11 = a_14_11 * b_11_13;
  assign t0_r14_c13_rr12 = a_14_12 * b_12_13;
  assign t0_r14_c13_rr13 = a_14_13 * b_13_13;
  assign t0_r14_c13_rr14 = a_14_14 * b_14_13;
  assign t1_r14_c13_rr0 = t0_r14_c13_rr0 + t0_r14_c13_rr1;
  assign t1_r14_c13_rr1 = t0_r14_c13_rr2 + t0_r14_c13_rr3;
  assign t1_r14_c13_rr2 = t0_r14_c13_rr4 + t0_r14_c13_rr5;
  assign t1_r14_c13_rr3 = t0_r14_c13_rr6 + t0_r14_c13_rr7;
  assign t1_r14_c13_rr4 = t0_r14_c13_rr8 + t0_r14_c13_rr9;
  assign t1_r14_c13_rr5 = t0_r14_c13_rr10 + t0_r14_c13_rr11;
  assign t1_r14_c13_rr6 = t0_r14_c13_rr12 + t0_r14_c13_rr13;
  assign t1_r14_c13_rr7 = t0_r14_c13_rr14;

  assign t2_r14_c13_rr0 = t1_r14_c13_rr0 + t1_r14_c13_rr1;
  assign t2_r14_c13_rr1 = t1_r14_c13_rr2 + t1_r14_c13_rr3;
  assign t2_r14_c13_rr2 = t1_r14_c13_rr4 + t1_r14_c13_rr5;
  assign t2_r14_c13_rr3 = t1_r14_c13_rr6 + t1_r14_c13_rr7;

  assign t3_r14_c13_rr0 = t2_r14_c13_rr0 + t2_r14_c13_rr1;
  assign t3_r14_c13_rr1 = t2_r14_c13_rr2 + t2_r14_c13_rr3;

  assign t4_r14_c13_rr0 = t3_r14_c13_rr0 + t3_r14_c13_rr1;

  assign c_14_13 = t4_r14_c13_rr0;
  assign t0_r14_c14_rr0 = a_14_0 * b_0_14;
  assign t0_r14_c14_rr1 = a_14_1 * b_1_14;
  assign t0_r14_c14_rr2 = a_14_2 * b_2_14;
  assign t0_r14_c14_rr3 = a_14_3 * b_3_14;
  assign t0_r14_c14_rr4 = a_14_4 * b_4_14;
  assign t0_r14_c14_rr5 = a_14_5 * b_5_14;
  assign t0_r14_c14_rr6 = a_14_6 * b_6_14;
  assign t0_r14_c14_rr7 = a_14_7 * b_7_14;
  assign t0_r14_c14_rr8 = a_14_8 * b_8_14;
  assign t0_r14_c14_rr9 = a_14_9 * b_9_14;
  assign t0_r14_c14_rr10 = a_14_10 * b_10_14;
  assign t0_r14_c14_rr11 = a_14_11 * b_11_14;
  assign t0_r14_c14_rr12 = a_14_12 * b_12_14;
  assign t0_r14_c14_rr13 = a_14_13 * b_13_14;
  assign t0_r14_c14_rr14 = a_14_14 * b_14_14;
  assign t1_r14_c14_rr0 = t0_r14_c14_rr0 + t0_r14_c14_rr1;
  assign t1_r14_c14_rr1 = t0_r14_c14_rr2 + t0_r14_c14_rr3;
  assign t1_r14_c14_rr2 = t0_r14_c14_rr4 + t0_r14_c14_rr5;
  assign t1_r14_c14_rr3 = t0_r14_c14_rr6 + t0_r14_c14_rr7;
  assign t1_r14_c14_rr4 = t0_r14_c14_rr8 + t0_r14_c14_rr9;
  assign t1_r14_c14_rr5 = t0_r14_c14_rr10 + t0_r14_c14_rr11;
  assign t1_r14_c14_rr6 = t0_r14_c14_rr12 + t0_r14_c14_rr13;
  assign t1_r14_c14_rr7 = t0_r14_c14_rr14;

  assign t2_r14_c14_rr0 = t1_r14_c14_rr0 + t1_r14_c14_rr1;
  assign t2_r14_c14_rr1 = t1_r14_c14_rr2 + t1_r14_c14_rr3;
  assign t2_r14_c14_rr2 = t1_r14_c14_rr4 + t1_r14_c14_rr5;
  assign t2_r14_c14_rr3 = t1_r14_c14_rr6 + t1_r14_c14_rr7;

  assign t3_r14_c14_rr0 = t2_r14_c14_rr0 + t2_r14_c14_rr1;
  assign t3_r14_c14_rr1 = t2_r14_c14_rr2 + t2_r14_c14_rr3;

  assign t4_r14_c14_rr0 = t3_r14_c14_rr0 + t3_r14_c14_rr1;

  assign c_14_14 = t4_r14_c14_rr0;
endmodule
