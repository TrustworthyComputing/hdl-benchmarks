module c7552(N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342, N241_O);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, 0950, 0951, 0952, 0953, 0954, 0955, 0956, 0957, 0958, 0959, 0960, 0961, 0962, 0963, 0964, 0965, 0966, 0967, 0968, 0969, 0970, 0971, 0972, 0973, 0974, 0975, 0976, 0977, 0978, 0979, 0980, 0981, 0982, 0983, 0984, 0985, 0986, 0987, 0988, 0989, 0990, 0991, 0992, 0993, 0994, 0995, 0996, 0997, 0998, 0999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165, 1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187, 1188, 1189, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198, 1199, 1200, 1201, 1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209, 1210, 1211, 1212, 1213, 1214, 1215, 1216, 1217, 1218, 1219, 1220, 1221, 1222, 1223, 1224, 1225, 1226, 1227, 1228, 1229, 1230, 1231, 1232, 1233, 1234, 1235, 1236, 1237, 1238, 1239, 1240, 1241, 1242, 1243, 1244, 1245, 1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264, 1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 1274, 1275, 1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 1286, 1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297, 1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308, 1309, 1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319, 1320, 1321, 1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361, 1362, 1363, 1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371, 1372, 1373, 1374, 1375, 1376, 1377, 1378, 1379, 1380, 1381, 1382, 1383, 1384, 1385, 1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 1394, 1395, 1396, 1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 1418, 1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429, 1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440, 1441, 1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451, 1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495, 1496, 1497, 1498, 1499, 1500, 1501, 1502, 1503, 1504, 1505, 1506, 1507, 1508, 1509, 1510, 1511, 1512, 1513, 1514, 1515, 1516, 1517, 1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550, 1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561, 1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572, 1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1601, 1602, 1603, 1604, 1605, 1606, 1607, 1608, 1609, 1610, 1611, 1612, 1613, 1614, 1615, 1616, 1617, 1618, 1619, 1620, 1621, 1622, 1623, 1624, 1625, 1626, 1627, 1628, 1629, 1630, 1631, 1632, 1633, 1634, 1635, 1636, 1637, 1638, 1639, 1640, 1641, 1642, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1651, 1652, 1653, 1654, 1655, 1656, 1657, 1658, 1659, 1660, 1661, 1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 1670, 1671, 1672, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1681, 1682, 1683, 1684, 1685, 1686, 1687, 1688, 1689, 1690, 1691, 1692, 1693, 1694, 1695, 1696, 1697, 1698, 1699, 1700, 1701, 1702, 1703, 1704, 1705, 1706, 1707, 1708, 1709, 1710, 1711, 1712, 1713, 1714, 1715, 1716, 1717, 1718, 1719, 1720, 1721, 1722, 1723, 1724, 1725, 1726, 1727, 1728, 1729, 1730, 1731, 1732, 1733, 1734, 1735, 1736, 1737, 1738, 1739, 1740, 1741, 1742, 1743, 1744, 1745, 1746, 1747, 1748, 1749, 1750, 1751, 1752, 1753, 1754, 1755, 1756, 1757, 1758, 1759, 1760, 1761, 1762, 1763, 1764, 1765, 1766, 1767, 1768, 1769, 1770, 1771, 1772, 1773, 1774, 1775, 1776, 1777, 1778, 1779, 1780, 1781, 1782, 1783, 1784, 1785, 1786, 1787, 1788, 1789, 1790, 1791, 1792, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1800, 1801, 1802, 1803, 1804, 1805, 1806, 1807, 1808, 1809, 1810, 1811, 1812, 1813, 1814, 1815, 1816, 1817, 1818, 1819, 1820, 1821, 1822, 1823, 1824, 1825, 1826, 1827, 1828, 1829, 1830, 1831, 1832, 1833, 1834, 1835, 1836, 1837, 1838, 1839, 1840, 1841, 1842, 1843, 1844, 1845, 1846, 1847, 1848, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1865, 1866, 1867, 1868, 1869, 1870, 1871, 1872, 1873, 1874, 1875, 1876, 1877, 1878, 1879, 1880, 1881, 1882, 1883, 1884, 1885, 1886, 1887, 1888, 1889, 1890, 1891, 1892, 1893, 1894, 1895, 1896, 1897, 1898, 1899, 1900, 1901, 1902, 1903, 1904, 1905, 1906, 1907, 1908, 1909, 1910, 1911, 1912, 1913, 1914, 1915, 1916, 1917, 1918, 1919, 1920, 1921, 1922, 1923, 1924, 1925, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933, 1934, 1935, 1936, 1937, 1938, 1939, 1940, 1941, 1942, 1943, N10778, N10781, N1116, N1125, N1136, N1147, N1160, N1175, N1182, N1233, N1244, N1249, N1256, N1270, N1277, N1287, N1299, N1308, N1311, N1428, N1431, N1828, N1829, N1830, N1833, N1840, N1841, N1842, N1843, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1913, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1997, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2240, N2267, N2275, N2287, N2293, N2309, N2315, N2331, N2347, N2368, N2384, N2390, N2406, N2412, N590, N614, N625, N636, N657, N676, N682, N689, N750, N871;
  input N1, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N12, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N15, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N18, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N23, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241_I, N242, N245, N248, N251, N254, N257, N26, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N29, N293, N296, N299, N303, N307, N310, N313, N316, N319, N32, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N35, N352, N355, N358, N361, N364, N367, N38, N382, N41, N44, N47, N5, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N9, N94, N97;
  output N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N1110, N1111, N1112, N1113, N1114, N11333, N11334, N11340, N11342, N1489, N1490, N1781, N241_O, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945;
  lut lut_gate1(0xb, N242, N5, N1110);
  lut lut_gate2(0xe, N57, N5, N881);
  lut lut_gate3(0x7, 1744, 1743, N882);
  lut lut_gate4(0x8, N150, N184, 1743);
  lut lut_gate5(0x8, N240, N228, 1744);
  lut lut_gate6(0x7, 1746, 1745, N883);
  lut lut_gate7(0x8, N210, N152, 1745);
  lut lut_gate8(0x8, N230, N218, 1746);
  lut lut_gate9(0x7, 1748, 1747, N884);
  lut lut_gate10(0x8, N183, N182, 1747);
  lut lut_gate11(0x8, N186, N185, 1748);
  lut lut_gate12(0x7, 1750, 1749, N885);
  lut lut_gate13(0x8, N162, N172, 1749);
  lut lut_gate14(0x8, N199, N188, 1750);
  lut lut_gate15(0x7, N134, 1751, N1113);
  lut lut_gate16(0x4, N133, N5, 1751);
  lut lut_gate17(0x6, N367, 1752, N10025);
  lut lut_gate18(0x1, 1755, 1753, 1752);
  lut lut_gate19(0x4, 1754, N310, 1753);
  lut lut_gate20(0x4, N41, N18, 1754);
  lut lut_gate21(0x8, N310, 1756, 1755);
  lut lut_gate22(0x1, N18, N41, 1756);
  lut lut_gate23(0x8, 1760, 1758, 1757);
  lut lut_gate24(0x8, 1759, 1752, 1758);
  lut lut_gate25(0x9, N313, 1484, 1759);
  lut lut_gate26(0x9, N316, 1485, 1760);
  lut lut_gate27(0x9, N319, 1486, 1761);
  lut lut_gate28(0x9, N322, 1487, 1762);
  lut lut_gate29(0x9, 1761, 1763, N10110);
  lut lut_gate30(0x1, 1764, 1483, 1763);
  lut lut_gate31(0x8, N367, 1757, 1764);
  lut lut_gate32(0x6, 1760, 1765, N10111);
  lut lut_gate33(0xb, 1668, 1766, 1765);
  lut lut_gate34(0x8, N367, 1758, 1766);
  lut lut_gate35(0x1, 1769, 1768, 1767);
  lut lut_gate36(0x8, N12, N9, 1768);
  lut lut_gate37(0x4, N18, N215, 1769);
  lut lut_gate38(0x1, 1771, 1768, 1770);
  lut lut_gate39(0x4, N18, N216, 1771);
  lut lut_gate40(0x1, 1773, 1768, 1772);
  lut lut_gate41(0x4, N18, N214, 1773);
  lut lut_gate42(0x1, 1775, 1768, 1774);
  lut lut_gate43(0x4, N18, N213, 1775);
  lut lut_gate44(0x9, N212, 1777, 1776);
  lut lut_gate45(0x6, N209, N211, 1777);
  lut lut_gate46(0x9, 1495, 1494, 1778);
  lut lut_gate47(0x9, 1498, 1497, 1779);
  lut lut_gate48(0x9, 1782, 1781, 1780);
  lut lut_gate49(0x6, 1500, 1499, 1781);
  lut lut_gate50(0x9, 1502, 1501, 1782);
  lut lut_gate51(0x9, 1484, 1485, 1783);
  lut lut_gate52(0x6, 1486, 1487, 1784);
  lut lut_gate53(0x9, 1787, 1786, 1785);
  lut lut_gate54(0x6, 1508, 1507, 1786);
  lut lut_gate55(0x9, 1510, 1509, 1787);
  lut lut_gate56(0x1, 1789, 1768, 1788);
  lut lut_gate57(0x4, N18, N153, 1789);
  lut lut_gate58(0x1, 1791, 1768, 1790);
  lut lut_gate59(0x4, N18, N154, 1791);
  lut lut_gate60(0x1, 1793, 1768, 1792);
  lut lut_gate61(0x4, N18, N156, 1793);
  lut lut_gate62(0x1, 1795, 1768, 1794);
  lut lut_gate63(0x4, N18, N155, 1795);
  lut lut_gate64(0x1, 1797, 1768, 1796);
  lut lut_gate65(0x4, N18, N157, 1797);
  lut lut_gate66(0x9, 1516, 1515, 1798);
  lut lut_gate67(0x9, 1530, 1529, 1799);
  lut lut_gate68(0x9, 1533, 1532, 1800);
  lut lut_gate69(0x6, 1803, 1802, 1801);
  lut lut_gate70(0x9, 1535, 1534, 1802);
  lut lut_gate71(0x6, 1537, 1536, 1803);
  lut lut_gate72(0x9, 1540, 1539, 1804);
  lut lut_gate73(0x9, N267, N263, 1805);
  lut lut_gate74(0x6, N271, N245, 1806);
  lut lut_gate75(0x9, 1542, 1541, 1807);
  lut lut_gate76(0x9, 1812, 1809, 1808);
  lut lut_gate77(0x6, 1811, 1810, 1809);
  lut lut_gate78(0x9, 1544, 1543, 1810);
  lut lut_gate79(0x6, 1546, 1545, 1811);
  lut lut_gate80(0x6, 1548, 1547, 1812);
  lut lut_gate81(0x6, 1550, 1549, 1813);
  lut lut_gate82(0x9, 1556, 1815, 1814);
  lut lut_gate83(0x6, 1555, 1554, 1815);
  lut lut_gate84(0x9, 1559, 1558, 1816);
  lut lut_gate85(0x9, 1562, 1818, 1817);
  lut lut_gate86(0x6, 1561, 1560, 1818);
  lut lut_gate87(0x1, 1820, 1768, 1819);
  lut lut_gate88(0x4, N18, N173, 1820);
  lut lut_gate89(0x1, 1822, 1768, 1821);
  lut lut_gate90(0x4, N18, N174, 1822);
  lut lut_gate91(0x1, 1824, 1768, 1823);
  lut lut_gate92(0x4, N18, N175, 1824);
  lut lut_gate93(0x1, 1826, 1768, 1825);
  lut lut_gate94(0x4, N18, N176, 1826);
  lut lut_gate95(0x1, 1828, 1768, 1827);
  lut lut_gate96(0x4, N18, N177, 1828);
  lut lut_gate97(0x9, 1569, 1568, 1829);
  lut lut_gate98(0x4, N18, N167, 1830);
  lut lut_gate99(0x1, 1832, 1768, 1831);
  lut lut_gate100(0x4, N18, N166, 1832);
  lut lut_gate101(0x9, N165, 1834, 1833);
  lut lut_gate102(0x6, N170, N164, 1834);
  lut lut_gate103(0x1, 1836, 1768, 1835);
  lut lut_gate104(0x4, N18, N168, 1836);
  lut lut_gate105(0x4, N18, N169, 1837);
  lut lut_gate106(0x1, 1837, 1768, 1838);
  lut lut_gate107(0x9, 1841, 1840, 1839);
  lut lut_gate108(0x6, 1574, 1573, 1840);
  lut lut_gate109(0x9, 1576, 1575, 1841);
  lut lut_gate110(0x6, 1844, 1843, 1842);
  lut lut_gate111(0x6, 1579, 1578, 1843);
  lut lut_gate112(0x9, 1581, 1580, 1844);
  lut lut_gate113(0x9, 1849, 1846, 1845);
  lut lut_gate114(0x9, 1848, 1847, 1846);
  lut lut_gate115(0x6, 1585, 1584, 1847);
  lut lut_gate116(0x9, 1587, 1586, 1848);
  lut lut_gate117(0x6, 1851, 1850, 1849);
  lut lut_gate118(0x6, 1589, 1588, 1850);
  lut lut_gate119(0x9, 1591, 1590, 1851);
  lut lut_gate120(0x6, 1879, 1593, N10632);
  lut lut_gate121(0x8, 1875, 1594, 1852);
  lut lut_gate122(0x4, 1507, N328, 1853);
  lut lut_gate123(0x4, 1508, N325, 1854);
  lut lut_gate124(0x4, N328, 1507, 1855);
  lut lut_gate125(0x8, 1860, 1857, 1856);
  lut lut_gate126(0x8, 1859, 1858, 1857);
  lut lut_gate127(0x9, N328, 1507, 1858);
  lut lut_gate128(0x9, N325, 1508, 1859);
  lut lut_gate129(0x6, N331, 1510, 1860);
  lut lut_gate130(0x1, 1865, 1862, 1861);
  lut lut_gate131(0x1, 1864, 1601, 1862);
  lut lut_gate132(0x4, 1496, N340, 1863);
  lut lut_gate133(0x4, 1495, N349, 1864);
  lut lut_gate134(0x4, N349, 1495, 1865);
  lut lut_gate135(0x8, 1872, 1867, 1866);
  lut lut_gate136(0x8, 1871, 1868, 1867);
  lut lut_gate137(0x8, 1870, 1869, 1868);
  lut lut_gate138(0x9, N346, 1497, 1869);
  lut lut_gate139(0x9, N343, 1498, 1870);
  lut lut_gate140(0x9, N340, 1496, 1871);
  lut lut_gate141(0x8, 1874, 1873, 1872);
  lut lut_gate142(0x9, N352, 1494, 1873);
  lut lut_gate143(0x9, N349, 1495, 1874);
  lut lut_gate144(0x8, 1877, 1876, 1875);
  lut lut_gate145(0x9, N358, 1499, 1876);
  lut lut_gate146(0x9, N355, 1500, 1877);
  lut lut_gate147(0x4, 1500, N355, 1878);
  lut lut_gate148(0x6, N277, 1514, 1879);
  lut lut_gate149(0x9, 1902, 1604, N10641);
  lut lut_gate150(0x4, 1895, 1605, 1880);
  lut lut_gate151(0x1, 1883, 1882, 1881);
  lut lut_gate152(0x1, N277, 1514, 1882);
  lut lut_gate153(0x1, N280, 1516, 1883);
  lut lut_gate154(0x8, N280, 1516, 1884);
  lut lut_gate155(0x4, 1511, N286, 1885);
  lut lut_gate156(0x4, N286, 1511, 1886);
  lut lut_gate157(0x8, 1892, 1888, 1887);
  lut lut_gate158(0x8, 1891, 1889, 1888);
  lut lut_gate159(0x8, 1890, 1879, 1889);
  lut lut_gate160(0x6, N280, 1516, 1890);
  lut lut_gate161(0x6, N283, 1515, 1891);
  lut lut_gate162(0x8, 1894, 1893, 1892);
  lut lut_gate163(0x9, N289, 1796, 1893);
  lut lut_gate164(0x9, N286, 1511, 1894);
  lut lut_gate165(0x8, 1899, 1896, 1895);
  lut lut_gate166(0x8, 1898, 1897, 1896);
  lut lut_gate167(0x9, N296, 1794, 1897);
  lut lut_gate168(0x9, N293, 1792, 1898);
  lut lut_gate169(0x9, N299, 1790, 1899);
  lut lut_gate170(0x9, N303, 1788, 1900);
  lut lut_gate171(0x4, 1792, N293, 1901);
  lut lut_gate172(0x9, N251, 1903, 1902);
  lut lut_gate173(0x1, 1904, 1768, 1903);
  lut lut_gate174(0x4, N18, N209, 1904);
  lut lut_gate175(0x4, 1608, 1888, 1905);
  lut lut_gate176(0x1, 1885, 1907, 1906);
  lut lut_gate177(0x1, 1886, 1905, 1907);
  lut lut_gate178(0x4, 1881, 1593, 1908);
  lut lut_gate179(0x8, N277, 1514, 1909);
  lut lut_gate180(0x6, 1923, 1910, N10715);
  lut lut_gate181(0xe, 1614, 1911, 1910);
  lut lut_gate182(0x4, 1912, 1604, 1911);
  lut lut_gate183(0x8, 1917, 1913, 1912);
  lut lut_gate184(0x8, 1902, 1914, 1913);
  lut lut_gate185(0x8, 1916, 1915, 1914);
  lut lut_gate186(0x9, N254, 1770, 1915);
  lut lut_gate187(0x9, N106, 1767, 1916);
  lut lut_gate188(0x9, N257, 1772, 1917);
  lut lut_gate189(0xe, 1922, 1919, 1918);
  lut lut_gate190(0x4, 1920, 1921, 1919);
  lut lut_gate191(0x4, 1903, N251, 1920);
  lut lut_gate192(0x4, N254, 1770, 1921);
  lut lut_gate193(0x4, 1770, N254, 1922);
  lut lut_gate194(0x9, N260, 1774, 1923);
  lut lut_gate195(0x6, 1917, 1924, N10716);
  lut lut_gate196(0xb, 1615, 1925, 1924);
  lut lut_gate197(0x4, 1913, 1604, 1925);
  lut lut_gate198(0x4, 1902, 1604, 1926);
  lut lut_gate199(0x9, 1915, 1927, N10718);
  lut lut_gate200(0x1, 1920, 1926, 1927);
  lut lut_gate201(0x7, 1932, 1928, N10729);
  lut lut_gate202(0x4, 1929, N10574, 1928);
  lut lut_gate203(0x8, 1931, 1930, 1929);
  lut lut_gate204(0x1, N883, N882, 1930);
  lut lut_gate205(0x1, N885, N884, 1931);
  lut lut_gate206(0x1, N10575, N10576, 1932);
  lut lut_gate207(0x6, 1871, 1595, N10827);
  lut lut_gate208(0x9, 1874, 1933, N10869);
  lut lut_gate209(0x1, 1601, 1934, 1933);
  lut lut_gate210(0x8, 1868, 1935, 1934);
  lut lut_gate211(0x8, 1871, 1595, 1935);
  lut lut_gate212(0x6, 1869, 1936, N10870);
  lut lut_gate213(0x1, 1619, 1937, 1936);
  lut lut_gate214(0x1, 1671, 1595, 1937);
  lut lut_gate215(0x4, N340, 1496, 1938);
  lut lut_gate216(0x9, 1870, 1939, N10871);
  lut lut_gate217(0x1, 1863, 1935, 1939);
  lut lut_gate218(0x8, N163, N1, N1781);
  lut lut_gate219(0x8, N382, N263, 1940);
  lut lut_gate220(0x8, N382, N267, 1941);
  lut lut_gate221(0x4, 1560, 1590, 1942);
  lut lut_gate222(0x4, 1592, 1557, 1943);
  lut lut_gate223(0x4, 1590, 1560, 1433);
  lut lut_gate224(0x1, 1436, 1435, 1434);
  lut lut_gate225(0x4, 1587, 1559, 1435);
  lut lut_gate226(0x4, 1586, 1558, 1436);
  lut lut_gate227(0x4, 1559, 1587, 1437);
  lut lut_gate228(0x4, 1440, 1439, 1438);
  lut lut_gate229(0x4, 1558, 1586, 1439);
  lut lut_gate230(0x9, 1585, 1555, 1440);
  lut lut_gate231(0x4, 1585, 1555, 1441);
  lut lut_gate232(0x1, 1444, 1443, 1442);
  lut lut_gate233(0x1, 1838, 1542, 1443);
  lut lut_gate234(0x1, 1835, 1541, 1444);
  lut lut_gate235(0x8, 1835, 1541, 1445);
  lut lut_gate236(0x8, 1825, 1535, 1446);
  lut lut_gate237(0x9, 1821, 1537, 1447);
  lut lut_gate238(0x6, 1448, 1596, N10350);
  lut lut_gate239(0x6, N334, 1509, 1448);
  lut lut_gate240(0x9, 1860, 1449, N10351);
  lut lut_gate241(0x1, 1599, 1450, 1449);
  lut lut_gate242(0x4, 1857, 1685, 1450);
  lut lut_gate243(0x4, N325, 1508, 1451);
  lut lut_gate244(0x9, 1859, 1685, N10353);
  lut lut_gate245(0x9, 1900, 1452, N10760);
  lut lut_gate246(0x4, 1673, 1880, 1452);
  lut lut_gate247(0x9, 1899, 1453, N10761);
  lut lut_gate248(0x4, 1609, 1454, 1453);
  lut lut_gate249(0x4, 1896, 1605, 1454);
  lut lut_gate250(0x4, N293, 1792, 1455);
  lut lut_gate251(0x9, 1898, 1605, N10763);
  lut lut_gate252(0x6, 1941, 1457, 1456);
  lut lut_gate253(0x1, N38, 1940, 1457);
  lut lut_gate254(0x6, 1458, 1621, N10839);
  lut lut_gate255(0x9, N38, 1940, 1458);
  lut lut_gate256(0x6, 1459, 1670, N10905);
  lut lut_gate257(0x9, N364, 1501, 1459);
  lut lut_gate258(0x9, 1461, 1460, N10906);
  lut lut_gate259(0x4, 1602, 1852, 1460);
  lut lut_gate260(0x9, N361, 1502, 1461);
  lut lut_gate261(0x4, 1594, 1463, 1462);
  lut lut_gate262(0x4, N355, 1500, 1463);
  lut lut_gate263(0x6, 1878, 1876, 1464);
  lut lut_gate264(0x6, 1877, 1594, N10908);
  lut lut_gate265(0x6, 1899, 1900, 1465);
  lut lut_gate266(0x6, 1468, 1467, 1466);
  lut lut_gate267(0x6, 1894, 1891, 1467);
  lut lut_gate268(0x6, 1893, 1890, 1468);
  lut lut_gate269(0x1, 1912, 1614, 1469);
  lut lut_gate270(0x4, 1615, 1913, 1470);
  lut lut_gate271(0x4, N251, 1903, 1471);
  lut lut_gate272(0x6, 1474, 1473, 1472);
  lut lut_gate273(0x6, 1916, 1915, 1473);
  lut lut_gate274(0x9, 1917, 1923, 1474);
  lut lut_gate275(0x9, 1477, 1476, 1475);
  lut lut_gate276(0x6, 1870, 1869, 1476);
  lut lut_gate277(0x6, 1874, 1873, 1477);
  lut lut_gate278(0x6, 1448, 1860, 1478);
  lut lut_gate279(0x9, 1481, 1480, 1479);
  lut lut_gate280(0x6, 1761, 1762, 1480);
  lut lut_gate281(0x6, 1759, 1760, 1481);
  lut lut_gate282(0x1, N15, N1111);
  lut lut_gate283(0x2b, 1486, 1483, N319, 1482);
  lut lut_gate284(0x71, 1485, 1668, N316, 1483);
  lut lut_gate285(0xca, N18, N238, N29, 1484);
  lut lut_gate286(0xca, N18, N237, N26, 1485);
  lut lut_gate287(0xca, N18, N236, N23, 1486);
  lut lut_gate288(0xca, N18, N235, N103, 1487);
  lut lut_gate289(0x0b, 1753, N367, 1755, 1488);
  lut lut_gate290(0x9, 1759, 1488, N10112);
  lut lut_gate291(0x6, 1513, 1511, 1489);
  lut lut_gate292(0x1, 1505, 1493, 1490);
  lut lut_gate293(0xca, N18, N227, N115, 1491);
  lut lut_gate294(0x96, 1779, 1496, 1778, 1492);
  lut lut_gate295(0x69, 1780, 1492, 1491, 1493);
  lut lut_gate296(0xca, N18, N223, N47, 1494);
  lut lut_gate297(0xca, N18, N224, N121, 1495);
  lut lut_gate298(0xca, N18, N217, N118, 1496);
  lut lut_gate299(0xca, N18, N225, N94, 1497);
  lut lut_gate300(0xca, N18, N226, N97, 1498);
  lut lut_gate301(0xca, N18, N221, N32, 1499);
  lut lut_gate302(0xca, N18, N222, N35, 1500);
  lut lut_gate303(0xca, N18, N219, N66, 1501);
  lut lut_gate304(0xca, N18, N220, N50, 1502);
  lut lut_gate305(0xca, N18, N239, N44, 1503);
  lut lut_gate306(0x96, 1784, 1783, 1506, 1504);
  lut lut_gate307(0x69, 1785, 1504, 1503, 1505);
  lut lut_gate308(0x53, N18, N41, N229, 1506);
  lut lut_gate309(0xca, N18, N233, N127, 1507);
  lut lut_gate310(0xca, N18, N234, N130, 1508);
  lut lut_gate311(0x35, N18, N231, N100, 1509);
  lut lut_gate312(0x35, N18, N232, N124, 1510);
  lut lut_gate313(0xca, N18, N158, N135, 1511);
  lut lut_gate314(0xca, N18, N161, N141, 1512);
  lut lut_gate315(0x69, 1798, 1514, 1512, 1513);
  lut lut_gate316(0x35, N18, N151, N147, 1514);
  lut lut_gate317(0x35, N18, N159, N144, 1515);
  lut lut_gate318(0x35, N18, N160, N138, 1516);
  lut lut_gate319(0x3a, N18, N310, N69, 1517);
  lut lut_gate320(0x78, 1677, N307, N18, 1518);
  lut lut_gate321(0x4, 1525, 1553, 1519);
  lut lut_gate322(0x6, 1813, 1808, 1520);
  lut lut_gate323(0x9f, 1519, 1520, 1518, N10575);
  lut lut_gate324(0x6, 1805, N248, 1521);
  lut lut_gate325(0x6, 1806, N114, 1522);
  lut lut_gate326(0xca, N18, 1521, 1522, 1523);
  lut lut_gate327(0x96, 1807, 1804, 1538, 1524);
  lut lut_gate328(0x60, 1528, 1524, 1523, 1525);
  lut lut_gate329(0xc5, N18, N274, N82, 1526);
  lut lut_gate330(0x96, 1800, 1531, 1799, 1527);
  lut lut_gate331(0x69, 1801, 1527, 1526, 1528);
  lut lut_gate332(0xc5, N18, N289, N64, 1529);
  lut lut_gate333(0xc5, N18, N286, N85, 1530);
  lut lut_gate334(0xc5, N18, N277, N65, 1531);
  lut lut_gate335(0x3a, N18, N283, N84, 1532);
  lut lut_gate336(0xc5, N18, N280, N83, 1533);
  lut lut_gate337(0x3a, N18, N296, N86, 1534);
  lut lut_gate338(0x3a, N18, N293, N63, 1535);
  lut lut_gate339(0x3a, N18, N303, N110, 1536);
  lut lut_gate340(0xc5, N18, N299, N109, 1537);
  lut lut_gate341(0x3a, N18, N251, N113, 1538);
  lut lut_gate342(0xc5, N18, N260, N88, 1539);
  lut lut_gate343(0xc5, N18, N257, N112, 1540);
  lut lut_gate344(0x3a, N18, N106, N87, 1541);
  lut lut_gate345(0x3a, N18, N254, N111, 1542);
  lut lut_gate346(0xc5, N18, N328, N54, 1543);
  lut lut_gate347(0xc5, N18, N325, N53, 1544);
  lut lut_gate348(0xc5, N18, N331, N55, 1545);
  lut lut_gate349(0x3a, N18, N334, N56, 1546);
  lut lut_gate350(0x3a, N18, N322, N73, 1547);
  lut lut_gate351(0xc5, N18, N319, N75, 1548);
  lut lut_gate352(0x3a, N18, N316, N76, 1549);
  lut lut_gate353(0xc5, N18, N313, N74, 1550);
  lut lut_gate354(0xc5, N18, N337, N58, 1551);
  lut lut_gate355(0x96, 1816, 1557, 1551, 1552);
  lut lut_gate356(0x96, 1817, 1814, 1552, 1553);
  lut lut_gate357(0x3a, N18, N352, N80, 1554);
  lut lut_gate358(0xc5, N18, N349, N81, 1555);
  lut lut_gate359(0xc5, N18, N355, N79, 1556);
  lut lut_gate360(0xc5, N18, N340, N77, 1557);
  lut lut_gate361(0xc5, N18, N346, N59, 1558);
  lut lut_gate362(0xc5, N18, N343, N78, 1559);
  lut lut_gate363(0xc5, N18, N364, N62, 1560);
  lut lut_gate364(0xc5, N18, N361, N61, 1561);
  lut lut_gate365(0x3a, N18, N358, N60, 1562);
  lut lut_gate366(0x94, 1831, 1830, 1768, 1563);
  lut lut_gate367(0xca, N18, N181, N141, 1564);
  lut lut_gate368(0x9, 1566, 1564, 1565);
  lut lut_gate369(0x35, N18, N171, N147, 1566);
  lut lut_gate370(0xca, N18, N178, N135, 1567);
  lut lut_gate371(0x35, N18, N179, N144, 1568);
  lut lut_gate372(0x35, N18, N180, N138, 1569);
  lut lut_gate373(0xca, N18, N208, N44, 1570);
  lut lut_gate374(0x96, 1842, 1577, 1839, 1571);
  lut lut_gate375(0x14, 1571, 1570, 1583, 1572);
  lut lut_gate376(0xca, N18, N206, N26, 1573);
  lut lut_gate377(0xca, N18, N207, N29, 1574);
  lut lut_gate378(0xca, N18, N204, N103, 1575);
  lut lut_gate379(0xca, N18, N205, N23, 1576);
  lut lut_gate380(0x53, N18, N41, N198, 1577);
  lut lut_gate381(0xca, N18, N202, N127, 1578);
  lut lut_gate382(0xca, N18, N203, N130, 1579);
  lut lut_gate383(0x35, N18, N200, N100, 1580);
  lut lut_gate384(0x35, N18, N201, N124, 1581);
  lut lut_gate385(0xca, N18, N197, N115, 1582);
  lut lut_gate386(0x69, 1592, 1845, 1582, 1583);
  lut lut_gate387(0xca, N18, N193, N47, 1584);
  lut lut_gate388(0xca, N18, N194, N121, 1585);
  lut lut_gate389(0xca, N18, N195, N94, 1586);
  lut lut_gate390(0xca, N18, N196, N97, 1587);
  lut lut_gate391(0xca, N18, N191, N32, 1588);
  lut lut_gate392(0xca, N18, N192, N35, 1589);
  lut lut_gate393(0xca, N18, N189, N66, 1590);
  lut lut_gate394(0xca, N18, N190, N50, 1591);
  lut lut_gate395(0xca, N18, N187, N118, 1592);
  lut lut_gate396(0x4, 1501, 1670, N364, 1593);
  lut lut_gate397(0x8f, 1600, 1866, 1595, 1594);
  lut lut_gate398(0x71, 1596, 1509, N334, 1595);
  lut lut_gate399(0xf4, 1598, 1856, 1685, 1596);
  lut lut_gate400(0x71, 1486, 1763, N319, 1597);
  lut lut_gate401(0x71, 1599, 1510, N331, 1598);
  lut lut_gate402(0x4, 1507, 1854, N328, 1599);
  lut lut_gate403(0x2b, 1494, 1861, N352, 1600);
  lut lut_gate404(0x4, 1497, 1671, N346, 1601);
  lut lut_gate405(0x2b, 1499, 1878, N358, 1602);
  lut lut_gate406(0x4, 1673, 1880, 1603);
  lut lut_gate407(0xb2, 1603, 1788, N303, 1604);
  lut lut_gate408(0x07, 1606, 1887, 1593, 1605);
  lut lut_gate409(0x4, 1672, 1796, N289, 1606);
  lut lut_gate410(0x1, 1884, 1881, 1607);
  lut lut_gate411(0xb2, 1515, 1607, N283, 1608);
  lut lut_gate412(0x2b, 1901, 1794, N296, 1609);
  lut lut_gate413(0x70, 1608, 1888, 1593, 1610);
  lut lut_gate414(0x9, 1894, 1610, N10712);
  lut lut_gate415(0x4f, 1907, 1608, 1593, 1611);
  lut lut_gate416(0x4b, 1893, 1611, 1885, N10711);
  lut lut_gate417(0x17, 1516, 1909, N280, 1612);
  lut lut_gate418(0xb4, 1891, 1612, 1908, N10713);
  lut lut_gate419(0x71, 1593, 1514, N277, 1613);
  lut lut_gate420(0x6, 1890, 1613, N10714);
  lut lut_gate421(0x71, 1772, 1615, N257, 1614);
  lut lut_gate422(0x2b, 1918, 1767, N106, 1615);
  lut lut_gate423(0x2b, 1926, 1770, N254, 1616);
  lut lut_gate424(0x4b, 1916, 1616, 1919, N10717);
  lut lut_gate425(0x8f, 1862, 1595, 1867, 1617);
  lut lut_gate426(0xb4, 1873, 1617, 1865, N10868);
  lut lut_gate427(0x0b, 1865, 1862, 1867, 1618);
  lut lut_gate428(0xb2, 1938, 1498, N343, 1619);
  lut lut_gate429(0x1, 1614, 1911, 1620);
  lut lut_gate430(0x71, 1774, 1620, N260, 1621);
  lut lut_gate431(0x2b, 1566, 1531, N10704, 1622);
  lut lut_gate432(0x71, 1546, 1580, 1692, 1623);
  lut lut_gate433(0x4, 1575, 1547, 1695, 1624);
  lut lut_gate434(0x2b, 1573, 1549, 1696, 1625);
  lut lut_gate435(0x17, N89, N70, N41, 1626);
  lut lut_gate436(0x5c, N18, 1626, N89, 1627);
  lut lut_gate437(0xb2, 1629, 1537, 1821, 1628);
  lut lut_gate438(0xe8, 1534, 1446, 1823, 1629);
  lut lut_gate439(0x71, 1508, 1685, N325, 1630);
  lut lut_gate440(0x6, 1858, 1630, N10352);
  lut lut_gate441(0x71, 1792, 1605, N293, 1631);
  lut lut_gate442(0x6, 1897, 1631, N10762);
  lut lut_gate443(0x53, 1621, 1632, 1456, N10837);
  lut lut_gate444(0x78, 1941, 1940, N38, 1632);
  lut lut_gate445(0x3a, 1462, 1876, 1464, N10907);
  lut lut_gate446(0x07, 1606, 1887, 1593, 1633);
  lut lut_gate447(0x69, 1637, 1466, 1702, N11333);
  lut lut_gate448(0xe3, 1673, 1703, 1895, 1634);
  lut lut_gate449(0x6, 1639, 1879, 1635);
  lut lut_gate450(0x3a, 1879, 1641, 1639, 1636);
  lut lut_gate451(0x3a, 1593, 1635, 1636, 1637);
  lut lut_gate452(0xca, 1909, 1883, 1884, 1638);
  lut lut_gate453(0x69, 1906, 1905, 1638, 1639);
  lut lut_gate454(0xca, 1882, 1884, 1883, 1640);
  lut lut_gate455(0x96, 1608, 1640, 1672, 1641);
  lut lut_gate456(0x9e, 1647, 1604, 1902, 1642);
  lut lut_gate457(0x70, 1642, 1650, 1604, 1643);
  lut lut_gate458(0xa3, 1621, 1456, 1632, 1644);
  lut lut_gate459(0x6, 1472, 1644, 1645);
  lut lut_gate460(0x9, 1645, 1643, N11334);
  lut lut_gate461(0xac, 1471, 1921, 1922, 1646);
  lut lut_gate462(0x96, 1470, 1469, 1646, 1647);
  lut lut_gate463(0xca, 1920, 1921, 1922, 1648);
  lut lut_gate464(0x96, 1615, 1614, 1648, 1649);
  lut lut_gate465(0x8, 1649, 1902, 1650);
  lut lut_gate466(0x70, 1600, 1866, 1595, 1651);
  lut lut_gate467(0x69, 1475, 1714, 1708, N11340);
  lut lut_gate468(0xc1, 1601, 1938, 1867, 1652);
  lut lut_gate469(0x96, 1619, 1618, 1652, 1653);
  lut lut_gate470(0x9e, 1657, 1752, N367, 1654);
  lut lut_gate471(0x9, 1661, 1717, N11342);
  lut lut_gate472(0x94, 1483, 1755, 1757, 1655);
  lut lut_gate473(0x43, 1482, 1757, 1761, 1656);
  lut lut_gate474(0x96, 1483, 1482, 1718, 1657);
  lut lut_gate475(0xc1, 1598, 1685, 1856, 1658);
  lut lut_gate476(0xc5, 1685, 1663, 1665, 1659);
  lut lut_gate477(0x6, 1479, 1478, 1660);
  lut lut_gate478(0x69, 1660, 1659, 1658, 1661);
  lut lut_gate479(0x1, 1857, 1853, 1662);
  lut lut_gate480(0xa3, 1451, 1662, 1855, 1663);
  lut lut_gate481(0xf8, 1508, N325, 1855, 1664);
  lut lut_gate482(0x9e, 1664, 1853, N325, 1665);
  lut lut_gate483(0x07, 1483, N367, 1757, 1666);
  lut lut_gate484(0x71, 1486, N319, 1666, 1667);
  lut lut_gate485(0x6, 1762, 1667, N10109);
  lut lut_gate486(0x2b, 1484, 1753, N313, 1668);
  lut lut_gate487(0x4, 1602, 1852, 1669);
  lut lut_gate488(0x71, 1502, 1669, N361, 1670);
  lut lut_gate489(0x4, 1498, 1863, N343, 1671);
  lut lut_gate490(0x71, 1511, 1608, N286, 1672);
  lut lut_gate491(0xb2, 1609, 1790, N299, 1673);
  lut lut_gate492(0x96, 1797, 1795, 1793, 1674);
  lut lut_gate493(0x69, 1674, 1791, 1789, 1675);
  lut lut_gate494(0x4b, 1489, 1675, 1768, 1676);
  lut lut_gate495(0x7f, 1490, 1676, 1721, N10574);
  lut lut_gate496(0xe1, 1517, N70, N18, 1677);
  lut lut_gate497(0x90, N18, 1833, N168, 1678);
  lut lut_gate498(0x41, 1837, 1678, 1768, 1679);
  lut lut_gate499(0xb4, 1820, 1828, 1768, 1680);
  lut lut_gate500(0x96, 1567, 1565, 1829, 1681);
  lut lut_gate501(0x96, 1826, 1824, 1822, 1682);
  lut lut_gate502(0x41, 1680, 1682, 1768, 1683);
  lut lut_gate503(0x90, 1572, 1679, 1563, 1684);
  lut lut_gate504(0x6f, 1684, 1681, 1683, N10576);
  lut lut_gate505(0x2b, 1597, 1487, N322, 1685);
  lut lut_gate506(0x81, 1941, 1940, N38, 1686);
  lut lut_gate507(0xac, 1686, N38, 1621, N10101);
  lut lut_gate508(0x0b, 1628, 1723, 1691, 1687);
  lut lut_gate509(0xb2, 1536, 1687, 1819, 1688);
  lut lut_gate510(0x8, 1724, N382, 1689);
  lut lut_gate511(0x4, 1725, N38, 1689, N10102);
  lut lut_gate512(0x71, 1532, 1568, 1726, 1690);
  lut lut_gate513(0x4, 1529, 1727, 1827, 1691);
  lut lut_gate514(0xe8, 1581, 1545, 1729, 1692);
  lut lut_gate515(0x41, 1592, 1557, 1433, 1693);
  lut lut_gate516(0x71, 1591, 1730, 1561, 1694);
  lut lut_gate517(0xf4, 1433, 1694, 1942, N10704);
  lut lut_gate518(0xb2, 1625, 1576, 1548, 1695);
  lut lut_gate519(0xb2, 1627, 1574, 1550, 1696);
  lut lut_gate520(0x42, 1609, 1790, N299, 1697);
  lut lut_gate521(0x6, 1455, 1697, 1698);
  lut lut_gate522(0x6, 1634, 1898, 1699);
  lut lut_gate523(0xca, 1633, 1698, 1699, 1700);
  lut lut_gate524(0x6, 1465, 1897, 1701);
  lut lut_gate525(0x6, 1701, 1700, 1702);
  lut lut_gate526(0x42, 1455, 1794, N296, 1703);
  lut lut_gate527(0xb0, 1602, 1875, 1651, 1704);
  lut lut_gate528(0xe7, 1502, 1704, N361, 1705);
  lut lut_gate529(0x6, 1459, 1876, 1706);
  lut lut_gate530(0xac, 1651, 1878, 1463, 1707);
  lut lut_gate531(0x96, 1707, 1706, 1705, 1708);
  lut lut_gate532(0x6, 1496, N340, 1709);
  lut lut_gate533(0x6, 1653, 1709, 1710);
  lut lut_gate534(0xb4, 1601, 1498, N343, 1711);
  lut lut_gate535(0x6, 1861, 1711, 1712);
  lut lut_gate536(0x35, 1709, 1653, 1712, 1713);
  lut lut_gate537(0x3a, 1595, 1710, 1713, 1714);
  lut lut_gate538(0xb4, 1656, 1668, 1759, 1715);
  lut lut_gate539(0x60, 1752, 1655, 1715, 1716);
  lut lut_gate540(0x70, 1654, N367, 1716, 1717);
  lut lut_gate541(0x18, 1484, 1753, N313, 1718);
  lut lut_gate542(0x90, N18, 1776, N215, 1719);
  lut lut_gate543(0x96, 1775, 1773, 1771, 1720);
  lut lut_gate544(0xeb, 1720, 1719, 1768, 1721);
  lut lut_gate545(0x60, 1447, 1535, 1825, 1722);
  lut lut_gate546(0x60, 1722, 1534, 1823, 1723);
  lut lut_gate547(0x17, N38, N271, N245, 1724);
  lut lut_gate548(0x2b, 1737, 1539, 1831, 1725);
  lut lut_gate549(0xb2, 1569, 1622, 1533, 1726);
  lut lut_gate550(0x2b, 1690, 1567, 1530, 1727);
  lut lut_gate551(0x2b, 1624, 1579, 1544, 1728);
  lut lut_gate552(0xb2, 1728, 1578, 1543, 1729);
  lut lut_gate553(0x2b, 1588, 1562, 1739, 1730);
  lut lut_gate554(0x4, 1542, 1837, 1731);
  lut lut_gate555(0xfe, 1688, 1538, 1731, 1732);
  lut lut_gate556(0x07, 1445, 1732, 1442, 1733);
  lut lut_gate557(0xe8, 1540, 1733, 1830, 1734);
  lut lut_gate558(0x7f, 1688, 1538, 1442, 1735);
  lut lut_gate559(0x0b, 1540, 1735, 1445, 1736);
  lut lut_gate560(0x3a, 1768, 1736, 1734, 1737);
  lut lut_gate561(0x2b, 1584, 1554, 1742, 1738);
  lut lut_gate562(0xb2, 1738, 1589, 1556, 1739);
  lut lut_gate563(0xf8, 1943, 1693, 1623, 1740);
  lut lut_gate564(0x4f, 1434, 1740, 1437, 1741);
  lut lut_gate565(0x07, 1441, 1741, 1438, 1742);

endmodule
