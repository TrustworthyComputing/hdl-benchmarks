module c6288(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G4, G5, G6, G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266, G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276, G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286, G6287, G6288, G7, G8, G9);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, 0950, 0951, 0952, 0953, 0954, 0955, 0956, 0957, 0958, 0959, 0960, 0961, 0962, 0963, 0964, 0965, 0966, 0967, 0968, 0969, 0970, 0971, 0972, 0973, 0974, 0975, 0976, 0977, 0978, 0979, 0980, 0981, 0982, 0983, 0984, 0985, 0986, 0987, 0988, 0989, 0990, 0991, 0992, 0993, 0994, 0995, 0996, 0997, 0998, 0999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165, 1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187, 1188, 1189, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198, 1199, 1200, 1201, 1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209, 1210, 1211, 1212, 1213, 1214, 1215, 1216, 1217, 1218, 1219, 1220, 1221, 1222, 1223, 1224, 1225, 1226, 1227, 1228, 1229, 1230, 1231, 1232, 1233, 1234, 1235, 1236, 1237, 1238, 1239, 1240, 1241, 1242, 1243, 1244, 1245, 1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264, 1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 1274, 1275, 1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 1286, 1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297, 1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308, 1309, 1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319, 1320, 1321, 1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361, 1362, 1363, 1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371, 1372, 1373, 1374, 1375, 1376, 1377, 1378, 1379, 1380, 1381, 1382, 1383, 1384, 1385, 1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 1394, 1395, 1396, 1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 1418, 1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429, 1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440, 1441, 1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451, 1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495, 1496, 1497, 1498, 1499, 1500, 1501, 1502, 1503, 1504, 1505, 1506, 1507, 1508, 1509, 1510, 1511, 1512, 1513, 1514, 1515, 1516, 1517, 1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550, 1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561, 1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572, 1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1601, 1602, 1603, 1604, 1605, 1606, 1607, 1608, 1609, 1610, 1611, 1612, 1613, 1614, 1615, 1616, 1617, 1618, 1619, 1620, 1621, 1622, 1623, 1624, 1625, 1626, 1627, 1628, 1629, 1630, 1631, 1632, 1633, 1634, 1635, 1636, 1637, 1638, 1639, 1640, 1641, 1642, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1651, 1652, 1653, 1654, 1655, 1656, 1657, 1658, 1659, 1660, 1661, 1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 1670, 1671, 1672, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1681, 1682, 1683, 1684, 1685, 1686, 1687, 1688, 1689, 1690, 1691, 1692, 1693, 1694, 1695, 1696, 1697, 1698, 1699, 1700, 1701, 1702, 1703, 1704, 1705, 1706, 1707, 1708, 1709, 1710, 1711, 1712, 1713, 1714, 1715, 1716, 1717, 1718, 1719, 1720, 1721, 1722, 1723, 1724, 1725, 1726, 1727, 1728, 1729, 1730, 1731, 1732, 1733, 1734, 1735, 1736, 1737, 1738, 1739, 1740, 1741, 1742, 1743, 1744, 1745, 1746, 1747, 1748, 1749, 1750, 1751, 1752, 1753, 1754, 1755, 1756, 1757, 1758, 1759, 1760, 1761, 1762, 1763, 1764, 1765, 1766, 1767, 1768, 1769, 1770, 1771, 1772, 1773, 1774, 1775, 1776, 1777, 1778, 1779, 1780, 1781, 1782, 1783, 1784, 1785, 1786, 1787, 1788, 1789, 1790, 1791, 1792, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1800, 1801, 1802, 1803, 1804, 1805, 1806, 1807, 1808, 1809, 1810, 1811, 1812, 1813, 1814, 1815, 1816, 1817, 1818, 1819, 1820, 1821, 1822, 1823, 1824, 1825, 1826, 1827, 1828, 1829, 1830, 1831, 1832, 1833, 1834, 1835, 1836, 1837, 1838, 1839, 1840, 1841, 1842, 1843, 1844, 1845, 1846, 1847, 1848, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1865, 1866, 1867, 1868, 1869, 1870, 1871, 1872, 1873, 1874, 1875, 1876, 1877, 1878, 1879, 1880, 1881, 1882, 1883, 1884, 1885, 1886, 1887, 1888, 1889, 1890, 1891, 1892, 1893, 1894, 1895, 1896, 1897, 1898, 1899, 1900, 1901, 1902, 1903, 1904, 1905, 1906, 1907, 1908, 1909, 1910, 1911, 1912, 1913, 1914, 1915, 1916, 1917, 1918, 1919, 1920, 1921, 1922, 1923, 1924, 1925, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933, 1934, 1935, 1936, 1937, 1938, 1939, 1940, 1941, 1942, 1943, 1944, 1945, 1946, 1947, 1948, 1949, 1950, 1951, 1952, 1953, 1954, 1955, 1956, 1957, 1958, 1959, 1960, 1961, 1962, 1963, 1964, 1965, 1966, 1967, 1968, 1969, 1970, 1971, 1972, 1973, 1974, 1975, 1976, 1977, 1978, 1979, 1980, 1981, 1982, 1983, 1984, 1985, 1986, 1987, 1988, 1989, 1990, 1991, 1992, 1993, 1994, 1995, 1996, 1997, 1998, 1999, 2000, 2001, 2002, 2003, 2004, 2005, 2006, 2007, 2008, 2009, 2010, 2011, 2012, 2013, 2014, 2015, 2016, 2017, 2018, 2019, 2020, 2021, 2022, 2023, 2024, 2025, 2026, 2027, 2028, 2029, 2030, 2031, 2032, 2033, 2034, 2035, 2036, 2037, 2038, 2039, 2040, 2041, 2042, 2043, 2044, 2045, 2046, 2047, 2048, 2049, 2050, 2051, 2052, 2053, 2054, 2055, 2056, 2057, 2058, 2059, 2060, 2061, 2062, 2063, 2064, 2065, 2066, 2067, 2068, 2069, 2070, 2071, 2072, 2073, 2074, 2075, 2076, 2077, 2078, 2079, 2080, 2081, 2082, 2083, 2084, 2085, 2086, 2087, 2088, 2089, 2090, 2091, 2092, 2093, 2094, 2095, 2096, 2097, 2098, 2099, 2100, 2101, 2102, 2103, 2104, 2105, 2106, 2107, 2108, 2109, 2110, 2111, 2112, 2113, 2114, 2115, 2116, 2117, 2118, 2119, 2120, 2121, 2122, 2123, 2124, 2125, 2126, 2127, 2128, 2129, 2130, 2131, 2132, 2133, 2134, 2135, 2136, 2137, 2138, 2139, 2140, 2141, 2142, 2143, 2144, 2145, 2146, 2147, 2148, 2149, 2150, 2151, 2152, 2153, 2154, 2155, 2156, 2157, 2158, 2159, 2160, 2161, 2162, 2163, 2164, 2165, 2166, 2167, 2168, 2169, 2170, 2171, 2172, 2173, 2174, 2175, 2176, 2177, 2178, 2179, 2180, 2181, 2182, 2183, 2184, 2185, 2186, 2187, 2188, 2189, 2190, 2191, 2192, 2193, 2194, 2195, 2196, 2197, 2198, 2199, 2200, 2201, 2202, 2203, 2204, 2205, 2206, 2207, 2208, 2209, 2210, 2211, 2212, 2213, 2214, 2215, 2216, 2217, 2218, 2219, 2220, 2221, 2222, 2223, 2224, 2225, 2226, 2227, 2228, 2229, 2230, 2231, 2232, 2233, 2234, 2235, 2236, 2237, 2238, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 2246, 2247, 2248, 2249, 2250, 2251, 2252, 2253, 2254, 2255, 2256, 2257, 2258, 2259, 2260, 2261, 2262, 2263, 2264, 2265, 2266, 2267, 2268, 2269, 2270, 2271, 2272, 2273, 2274, 2275, 2276, 2277, 2278, 2279, 2280, 2281, 2282, 2283, 2284, 2285, 2286, 2287, 2288, 2289, 2290, 2291, 2292, 2293, 2294, 2295, 2296, 2297, 2298, 2299, 2300, 2301, 2302, 2303, 2304, 2305, 2306, 2307, 2308, 2309, 2310, 2311, 2312, 2313, 2314, 2315, 2316, 2317, 2318, 2319, 2320, 2321, 2322, 2323, 2324, G1370, G1372, G1374, G1376, G1378, G1380, G1382, G1384, G1386, G1388, G1390, G1392, G1394, G1396, G1398, G6125, G6129;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G4, G5, G6, G7, G8, G9;
  output G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266, G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276, G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286, G6287, G6288;
  lut lut_gate1(0x6, 0081, 0299, G6277);
  lut lut_gate2(0x4, 0302, 0841, 0854);
  lut lut_gate3(0x9, 0797, 0303, 0867);
  lut lut_gate4(0x9, 0756, 0304, 0889);
  lut lut_gate5(0x9, 0718, 0305, 0902);
  lut lut_gate6(0x9, 0683, 0306, 0916);
  lut lut_gate7(0x9, 0651, 0307, 0937);
  lut lut_gate8(0x9, 0622, 0308, 0950);
  lut lut_gate9(0x9, 0596, 0309, 0969);
  lut lut_gate10(0x9, 0573, 0310, 0982);
  lut lut_gate11(0x9, 0553, 0311, 0068);
  lut lut_gate12(0x9, 0536, 0312, 0088);
  lut lut_gate13(0x9, 0317, 0313, 0101);
  lut lut_gate14(0x9, 0244, 0314, 0118);
  lut lut_gate15(0x9, 0195, 0315, 0131);
  lut lut_gate16(0x6, 0167, 0152, 0147);
  lut lut_gate17(0x8, 0162, 0157, 0152);
  lut lut_gate18(0x8, G2, G17, 0157);
  lut lut_gate19(0x8, G18, G1, 0162);
  lut lut_gate20(0x6, 0181, 0177, 0167);
  lut lut_gate21(0x8, G3, G17, 0177);
  lut lut_gate22(0x8, G18, G2, 0181);
  lut lut_gate23(0x8, G19, G1, 0186);
  lut lut_gate24(0x9, 0230, 0204, 0195);
  lut lut_gate25(0x6, 0213, 0208, 0204);
  lut lut_gate26(0x8, 0181, 0177, 0208);
  lut lut_gate27(0x6, 0223, 0218, 0213);
  lut lut_gate28(0x8, G4, G17, 0218);
  lut lut_gate29(0x8, G18, G3, 0223);
  lut lut_gate30(0x8, G19, G2, 0230);
  lut lut_gate31(0x8, G20, G1, 0235);
  lut lut_gate32(0x9, 0297, 0250, 0244);
  lut lut_gate33(0x9, 0267, 0316, 0250);
  lut lut_gate34(0x9, 0296, 0272, 0267);
  lut lut_gate35(0x6, 0283, 0278, 0272);
  lut lut_gate36(0x8, 0223, 0218, 0278);
  lut lut_gate37(0x6, 0293, 0288, 0283);
  lut lut_gate38(0x8, G5, G17, 0288);
  lut lut_gate39(0x8, G4, G18, 0293);
  lut lut_gate40(0x8, G19, G3, 0296);
  lut lut_gate41(0x8, G20, G2, 0297);
  lut lut_gate42(0x8, G21, G1, 0298);
  lut lut_gate43(0x9, 0509, 0328, 0317);
  lut lut_gate44(0x9, 0369, 0318, 0328);
  lut lut_gate45(0x9, 0498, 0380, 0369);
  lut lut_gate46(0x9, 0421, 0319, 0380);
  lut lut_gate47(0x9, 0487, 0432, 0421);
  lut lut_gate48(0x6, 0454, 0443, 0432);
  lut lut_gate49(0x8, 0293, 0288, 0443);
  lut lut_gate50(0x6, 0476, 0465, 0454);
  lut lut_gate51(0x8, G5, G18, 0465);
  lut lut_gate52(0x8, G17, G6, 0476);
  lut lut_gate53(0x8, G4, G19, 0487);
  lut lut_gate54(0x8, G20, G3, 0498);
  lut lut_gate55(0x8, G21, G2, 0509);
  lut lut_gate56(0x8, G22, G1, 0520);
  lut lut_gate57(0x9, 0551, 0537, 0536);
  lut lut_gate58(0x9, 0538, 0320, 0537);
  lut lut_gate59(0x9, 0550, 0539, 0538);
  lut lut_gate60(0x9, 0540, 0321, 0539);
  lut lut_gate61(0x9, 0549, 0541, 0540);
  lut lut_gate62(0x9, 0542, 0322, 0541);
  lut lut_gate63(0x9, 0548, 0543, 0542);
  lut lut_gate64(0x6, 0545, 0544, 0543);
  lut lut_gate65(0x8, 0476, 0465, 0544);
  lut lut_gate66(0x6, 0547, 0546, 0545);
  lut lut_gate67(0x8, G18, G6, 0546);
  lut lut_gate68(0x8, G17, G7, 0547);
  lut lut_gate69(0x8, G5, G19, 0548);
  lut lut_gate70(0x8, G20, G4, 0549);
  lut lut_gate71(0x8, G21, G3, 0550);
  lut lut_gate72(0x8, G22, G2, 0551);
  lut lut_gate73(0x8, G1, G23, 0552);
  lut lut_gate74(0x9, 0571, 0554, 0553);
  lut lut_gate75(0x9, 0555, 0323, 0554);
  lut lut_gate76(0x9, 0570, 0556, 0555);
  lut lut_gate77(0x9, 0557, 0324, 0556);
  lut lut_gate78(0x9, 0569, 0558, 0557);
  lut lut_gate79(0x9, 0559, 0325, 0558);
  lut lut_gate80(0x9, 0568, 0560, 0559);
  lut lut_gate81(0x9, 0561, 0326, 0560);
  lut lut_gate82(0x9, 0567, 0562, 0561);
  lut lut_gate83(0x6, 0564, 0563, 0562);
  lut lut_gate84(0x8, 0547, 0546, 0563);
  lut lut_gate85(0x6, 0566, 0565, 0564);
  lut lut_gate86(0x8, G18, G7, 0565);
  lut lut_gate87(0x8, G17, G8, 0566);
  lut lut_gate88(0x8, G19, G6, 0567);
  lut lut_gate89(0x8, G5, G20, 0568);
  lut lut_gate90(0x8, G21, G4, 0569);
  lut lut_gate91(0x8, G22, G3, 0570);
  lut lut_gate92(0x8, G2, G23, 0571);
  lut lut_gate93(0x8, G1, G24, 0572);
  lut lut_gate94(0x9, 0594, 0574, 0573);
  lut lut_gate95(0x9, 0575, 0327, 0574);
  lut lut_gate96(0x9, 0593, 0576, 0575);
  lut lut_gate97(0x9, 0577, 0329, 0576);
  lut lut_gate98(0x9, 0592, 0578, 0577);
  lut lut_gate99(0x9, 0579, 0330, 0578);
  lut lut_gate100(0x9, 0591, 0580, 0579);
  lut lut_gate101(0x9, 0581, 0331, 0580);
  lut lut_gate102(0x9, 0590, 0582, 0581);
  lut lut_gate103(0x9, 0583, 0332, 0582);
  lut lut_gate104(0x9, 0589, 0584, 0583);
  lut lut_gate105(0x6, 0586, 0585, 0584);
  lut lut_gate106(0x8, 0566, 0565, 0585);
  lut lut_gate107(0x6, 0588, 0587, 0586);
  lut lut_gate108(0x8, G18, G8, 0587);
  lut lut_gate109(0x8, G17, G9, 0588);
  lut lut_gate110(0x8, G19, G7, 0589);
  lut lut_gate111(0x8, G20, G6, 0590);
  lut lut_gate112(0x8, G21, G5, 0591);
  lut lut_gate113(0x8, G22, G4, 0592);
  lut lut_gate114(0x8, G3, G23, 0593);
  lut lut_gate115(0x8, G2, G24, 0594);
  lut lut_gate116(0x8, G1, G25, 0595);
  lut lut_gate117(0x9, 0620, 0597, 0596);
  lut lut_gate118(0x9, 0598, 0333, 0597);
  lut lut_gate119(0x9, 0619, 0599, 0598);
  lut lut_gate120(0x9, 0600, 0334, 0599);
  lut lut_gate121(0x9, 0618, 0601, 0600);
  lut lut_gate122(0x9, 0602, 0335, 0601);
  lut lut_gate123(0x9, 0617, 0603, 0602);
  lut lut_gate124(0x9, 0604, 0336, 0603);
  lut lut_gate125(0x9, 0616, 0605, 0604);
  lut lut_gate126(0x9, 0606, 0337, 0605);
  lut lut_gate127(0x9, 0615, 0607, 0606);
  lut lut_gate128(0x9, 0608, 0338, 0607);
  lut lut_gate129(0x9, 0614, 0609, 0608);
  lut lut_gate130(0x6, 0611, 0610, 0609);
  lut lut_gate131(0x8, 0588, 0587, 0610);
  lut lut_gate132(0x6, 0613, 0612, 0611);
  lut lut_gate133(0x8, G18, G9, 0612);
  lut lut_gate134(0x8, G17, G10, 0613);
  lut lut_gate135(0x8, G19, G8, 0614);
  lut lut_gate136(0x8, G20, G7, 0615);
  lut lut_gate137(0x8, G21, G6, 0616);
  lut lut_gate138(0x8, G22, G5, 0617);
  lut lut_gate139(0x8, G4, G23, 0618);
  lut lut_gate140(0x8, G3, G24, 0619);
  lut lut_gate141(0x8, G2, G25, 0620);
  lut lut_gate142(0x8, G1, G26, 0621);
  lut lut_gate143(0x9, 0649, 0623, 0622);
  lut lut_gate144(0x9, 0624, 0339, 0623);
  lut lut_gate145(0x9, 0648, 0625, 0624);
  lut lut_gate146(0x9, 0626, 0340, 0625);
  lut lut_gate147(0x9, 0647, 0627, 0626);
  lut lut_gate148(0x9, 0628, 0341, 0627);
  lut lut_gate149(0x9, 0646, 0629, 0628);
  lut lut_gate150(0x9, 0630, 0342, 0629);
  lut lut_gate151(0x9, 0645, 0631, 0630);
  lut lut_gate152(0x9, 0632, 0343, 0631);
  lut lut_gate153(0x9, 0644, 0633, 0632);
  lut lut_gate154(0x9, 0634, 0344, 0633);
  lut lut_gate155(0x9, 0643, 0635, 0634);
  lut lut_gate156(0x9, 0636, 0345, 0635);
  lut lut_gate157(0x9, 0642, 0637, 0636);
  lut lut_gate158(0x6, 0639, 0638, 0637);
  lut lut_gate159(0x8, 0613, 0612, 0638);
  lut lut_gate160(0x6, 0641, 0640, 0639);
  lut lut_gate161(0x8, G18, G10, 0640);
  lut lut_gate162(0x8, G17, G11, 0641);
  lut lut_gate163(0x8, G19, G9, 0642);
  lut lut_gate164(0x8, G20, G8, 0643);
  lut lut_gate165(0x8, G21, G7, 0644);
  lut lut_gate166(0x8, G22, G6, 0645);
  lut lut_gate167(0x8, G5, G23, 0646);
  lut lut_gate168(0x8, G4, G24, 0647);
  lut lut_gate169(0x8, G3, G25, 0648);
  lut lut_gate170(0x8, G2, G26, 0649);
  lut lut_gate171(0x8, G1, G27, 0650);
  lut lut_gate172(0x9, 0681, 0652, 0651);
  lut lut_gate173(0x9, 0653, 0346, 0652);
  lut lut_gate174(0x9, 0680, 0654, 0653);
  lut lut_gate175(0x9, 0655, 0347, 0654);
  lut lut_gate176(0x9, 0679, 0656, 0655);
  lut lut_gate177(0x9, 0657, 0348, 0656);
  lut lut_gate178(0x9, 0678, 0658, 0657);
  lut lut_gate179(0x9, 0659, 0349, 0658);
  lut lut_gate180(0x9, 0677, 0660, 0659);
  lut lut_gate181(0x9, 0661, 0350, 0660);
  lut lut_gate182(0x9, 0676, 0662, 0661);
  lut lut_gate183(0x9, 0663, 0351, 0662);
  lut lut_gate184(0x9, 0675, 0664, 0663);
  lut lut_gate185(0x9, 0665, 0352, 0664);
  lut lut_gate186(0x9, 0674, 0666, 0665);
  lut lut_gate187(0x9, 0667, 0353, 0666);
  lut lut_gate188(0x9, 0673, 0668, 0667);
  lut lut_gate189(0x6, 0670, 0669, 0668);
  lut lut_gate190(0x8, 0641, 0640, 0669);
  lut lut_gate191(0x6, 0672, 0671, 0670);
  lut lut_gate192(0x8, G18, G11, 0671);
  lut lut_gate193(0x8, G17, G12, 0672);
  lut lut_gate194(0x8, G19, G10, 0673);
  lut lut_gate195(0x8, G20, G9, 0674);
  lut lut_gate196(0x8, G21, G8, 0675);
  lut lut_gate197(0x8, G22, G7, 0676);
  lut lut_gate198(0x8, G23, G6, 0677);
  lut lut_gate199(0x8, G5, G24, 0678);
  lut lut_gate200(0x8, G4, G25, 0679);
  lut lut_gate201(0x8, G3, G26, 0680);
  lut lut_gate202(0x8, G2, G27, 0681);
  lut lut_gate203(0x8, G1, G28, 0682);
  lut lut_gate204(0x9, 0716, 0684, 0683);
  lut lut_gate205(0x9, 0685, 0354, 0684);
  lut lut_gate206(0x9, 0715, 0686, 0685);
  lut lut_gate207(0x9, 0687, 0355, 0686);
  lut lut_gate208(0x9, 0714, 0688, 0687);
  lut lut_gate209(0x9, 0689, 0356, 0688);
  lut lut_gate210(0x9, 0713, 0690, 0689);
  lut lut_gate211(0x9, 0691, 0357, 0690);
  lut lut_gate212(0x9, 0712, 0692, 0691);
  lut lut_gate213(0x9, 0693, 0358, 0692);
  lut lut_gate214(0x9, 0711, 0694, 0693);
  lut lut_gate215(0x9, 0695, 0359, 0694);
  lut lut_gate216(0x9, 0710, 0696, 0695);
  lut lut_gate217(0x9, 0697, 0360, 0696);
  lut lut_gate218(0x9, 0709, 0698, 0697);
  lut lut_gate219(0x9, 0699, 0361, 0698);
  lut lut_gate220(0x9, 0708, 0700, 0699);
  lut lut_gate221(0x9, 0701, 0362, 0700);
  lut lut_gate222(0x9, 0707, 0702, 0701);
  lut lut_gate223(0x6, 0704, 0703, 0702);
  lut lut_gate224(0x8, 0672, 0671, 0703);
  lut lut_gate225(0x6, 0706, 0705, 0704);
  lut lut_gate226(0x8, G18, G12, 0705);
  lut lut_gate227(0x8, G17, G13, 0706);
  lut lut_gate228(0x8, G19, G11, 0707);
  lut lut_gate229(0x8, G20, G10, 0708);
  lut lut_gate230(0x8, G21, G9, 0709);
  lut lut_gate231(0x8, G22, G8, 0710);
  lut lut_gate232(0x8, G23, G7, 0711);
  lut lut_gate233(0x8, G24, G6, 0712);
  lut lut_gate234(0x8, G5, G25, 0713);
  lut lut_gate235(0x8, G4, G26, 0714);
  lut lut_gate236(0x8, G3, G27, 0715);
  lut lut_gate237(0x8, G2, G28, 0716);
  lut lut_gate238(0x8, G1, G29, 0717);
  lut lut_gate239(0x9, 0754, 0719, 0718);
  lut lut_gate240(0x9, 0720, 0363, 0719);
  lut lut_gate241(0x9, 0753, 0721, 0720);
  lut lut_gate242(0x9, 0722, 0364, 0721);
  lut lut_gate243(0x9, 0752, 0723, 0722);
  lut lut_gate244(0x9, 0724, 0365, 0723);
  lut lut_gate245(0x9, 0751, 0725, 0724);
  lut lut_gate246(0x9, 0726, 0366, 0725);
  lut lut_gate247(0x9, 0750, 0727, 0726);
  lut lut_gate248(0x9, 0728, 0367, 0727);
  lut lut_gate249(0x9, 0749, 0729, 0728);
  lut lut_gate250(0x9, 0730, 0368, 0729);
  lut lut_gate251(0x9, 0748, 0731, 0730);
  lut lut_gate252(0x9, 0732, 0370, 0731);
  lut lut_gate253(0x9, 0747, 0733, 0732);
  lut lut_gate254(0x9, 0734, 0371, 0733);
  lut lut_gate255(0x9, 0746, 0735, 0734);
  lut lut_gate256(0x9, 0736, 0372, 0735);
  lut lut_gate257(0x9, 0745, 0737, 0736);
  lut lut_gate258(0x9, 0738, 0373, 0737);
  lut lut_gate259(0x9, 0744, 0739, 0738);
  lut lut_gate260(0x6, 0741, 0740, 0739);
  lut lut_gate261(0x8, 0706, 0705, 0740);
  lut lut_gate262(0x6, 0743, 0742, 0741);
  lut lut_gate263(0x8, G18, G13, 0742);
  lut lut_gate264(0x8, G17, G14, 0743);
  lut lut_gate265(0x8, G19, G12, 0744);
  lut lut_gate266(0x8, G20, G11, 0745);
  lut lut_gate267(0x8, G21, G10, 0746);
  lut lut_gate268(0x8, G22, G9, 0747);
  lut lut_gate269(0x8, G23, G8, 0748);
  lut lut_gate270(0x8, G24, G7, 0749);
  lut lut_gate271(0x8, G25, G6, 0750);
  lut lut_gate272(0x8, G5, G26, 0751);
  lut lut_gate273(0x8, G4, G27, 0752);
  lut lut_gate274(0x8, G3, G28, 0753);
  lut lut_gate275(0x8, G2, G29, 0754);
  lut lut_gate276(0x8, G1, G30, 0755);
  lut lut_gate277(0x9, 0795, 0757, 0756);
  lut lut_gate278(0x9, 0758, 0374, 0757);
  lut lut_gate279(0x9, 0794, 0759, 0758);
  lut lut_gate280(0x9, 0760, 0375, 0759);
  lut lut_gate281(0x9, 0793, 0761, 0760);
  lut lut_gate282(0x9, 0762, 0376, 0761);
  lut lut_gate283(0x9, 0792, 0763, 0762);
  lut lut_gate284(0x9, 0764, 0377, 0763);
  lut lut_gate285(0x9, 0791, 0765, 0764);
  lut lut_gate286(0x9, 0766, 0378, 0765);
  lut lut_gate287(0x9, 0790, 0767, 0766);
  lut lut_gate288(0x9, 0768, 0379, 0767);
  lut lut_gate289(0x9, 0789, 0769, 0768);
  lut lut_gate290(0x9, 0770, 0381, 0769);
  lut lut_gate291(0x9, 0788, 0771, 0770);
  lut lut_gate292(0x9, 0772, 0382, 0771);
  lut lut_gate293(0x9, 0787, 0773, 0772);
  lut lut_gate294(0x9, 0774, 0383, 0773);
  lut lut_gate295(0x9, 0786, 0775, 0774);
  lut lut_gate296(0x9, 0776, 0384, 0775);
  lut lut_gate297(0x9, 0785, 0777, 0776);
  lut lut_gate298(0x9, 0778, 0385, 0777);
  lut lut_gate299(0x9, 0784, 0779, 0778);
  lut lut_gate300(0x6, 0781, 0780, 0779);
  lut lut_gate301(0x8, 0743, 0742, 0780);
  lut lut_gate302(0x6, 0783, 0782, 0781);
  lut lut_gate303(0x8, G18, G14, 0782);
  lut lut_gate304(0x8, G17, G15, 0783);
  lut lut_gate305(0x8, G19, G13, 0784);
  lut lut_gate306(0x8, G20, G12, 0785);
  lut lut_gate307(0x8, G21, G11, 0786);
  lut lut_gate308(0x8, G22, G10, 0787);
  lut lut_gate309(0x8, G23, G9, 0788);
  lut lut_gate310(0x8, G24, G8, 0789);
  lut lut_gate311(0x8, G25, G7, 0790);
  lut lut_gate312(0x8, G26, G6, 0791);
  lut lut_gate313(0x8, G5, G27, 0792);
  lut lut_gate314(0x8, G4, G28, 0793);
  lut lut_gate315(0x8, G3, G29, 0794);
  lut lut_gate316(0x8, G2, G30, 0795);
  lut lut_gate317(0x8, G1, G31, 0796);
  lut lut_gate318(0x9, 0839, 0798, 0797);
  lut lut_gate319(0x9, 0799, 0386, 0798);
  lut lut_gate320(0x9, 0838, 0800, 0799);
  lut lut_gate321(0x9, 0801, 0387, 0800);
  lut lut_gate322(0x9, 0837, 0802, 0801);
  lut lut_gate323(0x9, 0803, 0388, 0802);
  lut lut_gate324(0x9, 0836, 0804, 0803);
  lut lut_gate325(0x9, 0805, 0389, 0804);
  lut lut_gate326(0x9, 0835, 0806, 0805);
  lut lut_gate327(0x9, 0807, 0390, 0806);
  lut lut_gate328(0x9, 0834, 0808, 0807);
  lut lut_gate329(0x9, 0809, 0391, 0808);
  lut lut_gate330(0x9, 0833, 0810, 0809);
  lut lut_gate331(0x9, 0811, 0392, 0810);
  lut lut_gate332(0x9, 0832, 0812, 0811);
  lut lut_gate333(0x9, 0813, 0393, 0812);
  lut lut_gate334(0x9, 0831, 0814, 0813);
  lut lut_gate335(0x9, 0815, 0394, 0814);
  lut lut_gate336(0x9, 0830, 0816, 0815);
  lut lut_gate337(0x9, 0817, 0395, 0816);
  lut lut_gate338(0x9, 0829, 0818, 0817);
  lut lut_gate339(0x9, 0819, 0396, 0818);
  lut lut_gate340(0x9, 0828, 0820, 0819);
  lut lut_gate341(0x9, 0821, 0397, 0820);
  lut lut_gate342(0x9, 0827, 0822, 0821);
  lut lut_gate343(0x6, 0825, 0823, 0822);
  lut lut_gate344(0x8, 0824, 0743, 0823);
  lut lut_gate345(0x8, G18, G15, 0824);
  lut lut_gate346(0x6, 0826, 0824, 0825);
  lut lut_gate347(0x8, G17, G16, 0826);
  lut lut_gate348(0x8, G19, G14, 0827);
  lut lut_gate349(0x8, G20, G13, 0828);
  lut lut_gate350(0x8, G21, G12, 0829);
  lut lut_gate351(0x8, G22, G11, 0830);
  lut lut_gate352(0x8, G23, G10, 0831);
  lut lut_gate353(0x8, G24, G9, 0832);
  lut lut_gate354(0x8, G25, G8, 0833);
  lut lut_gate355(0x8, G26, G7, 0834);
  lut lut_gate356(0x8, G27, G6, 0835);
  lut lut_gate357(0x8, G5, G28, 0836);
  lut lut_gate358(0x8, G4, G29, 0837);
  lut lut_gate359(0x8, G3, G30, 0838);
  lut lut_gate360(0x8, G2, G31, 0839);
  lut lut_gate361(0x8, G1, G32, 0840);
  lut lut_gate362(0x9, 0885, 0842, 0841);
  lut lut_gate363(0x9, 0843, 0398, 0842);
  lut lut_gate364(0x9, 0884, 0844, 0843);
  lut lut_gate365(0x9, 0845, 0399, 0844);
  lut lut_gate366(0x9, 0883, 0846, 0845);
  lut lut_gate367(0x9, 0847, 0400, 0846);
  lut lut_gate368(0x9, 0882, 0848, 0847);
  lut lut_gate369(0x9, 0849, 0401, 0848);
  lut lut_gate370(0x9, 0881, 0850, 0849);
  lut lut_gate371(0x9, 0851, 0402, 0850);
  lut lut_gate372(0x9, 0880, 0852, 0851);
  lut lut_gate373(0x9, 0853, 0403, 0852);
  lut lut_gate374(0x9, 0879, 0855, 0853);
  lut lut_gate375(0x9, 0856, 0404, 0855);
  lut lut_gate376(0x9, 0878, 0857, 0856);
  lut lut_gate377(0x9, 0858, 0405, 0857);
  lut lut_gate378(0x9, 0877, 0859, 0858);
  lut lut_gate379(0x9, 0860, 0406, 0859);
  lut lut_gate380(0x9, 0876, 0861, 0860);
  lut lut_gate381(0x9, 0862, 0407, 0861);
  lut lut_gate382(0x9, 0875, 0863, 0862);
  lut lut_gate383(0x9, 0864, 0408, 0863);
  lut lut_gate384(0x9, 0874, 0865, 0864);
  lut lut_gate385(0x9, 0866, 0409, 0865);
  lut lut_gate386(0x9, 0873, 0868, 0866);
  lut lut_gate387(0x9, 0869, 0410, 0868);
  lut lut_gate388(0x9, 0872, 0870, 0869);
  lut lut_gate389(0x4, 0871, 0783, 0870);
  lut lut_gate390(0x8, G18, G16, 0871);
  lut lut_gate391(0x8, G19, G15, 0872);
  lut lut_gate392(0x8, G20, G14, 0873);
  lut lut_gate393(0x8, G21, G13, 0874);
  lut lut_gate394(0x8, G22, G12, 0875);
  lut lut_gate395(0x8, G11, G23, 0876);
  lut lut_gate396(0x8, G24, G10, 0877);
  lut lut_gate397(0x8, G25, G9, 0878);
  lut lut_gate398(0x8, G26, G8, 0879);
  lut lut_gate399(0x8, G27, G7, 0880);
  lut lut_gate400(0x8, G6, G28, 0881);
  lut lut_gate401(0x8, G5, G29, 0882);
  lut lut_gate402(0x8, G4, G30, 0883);
  lut lut_gate403(0x8, G3, G31, 0884);
  lut lut_gate404(0x8, G2, G32, 0885);
  lut lut_gate405(0x9, 0887, 0411, 0886);
  lut lut_gate406(0x9, 0929, 0888, 0887);
  lut lut_gate407(0x9, 0890, 0412, 0888);
  lut lut_gate408(0x9, 0928, 0891, 0890);
  lut lut_gate409(0x9, 0892, 0413, 0891);
  lut lut_gate410(0x9, 0927, 0893, 0892);
  lut lut_gate411(0x9, 0894, 0414, 0893);
  lut lut_gate412(0x9, 0926, 0895, 0894);
  lut lut_gate413(0x9, 0896, 0415, 0895);
  lut lut_gate414(0x9, 0925, 0897, 0896);
  lut lut_gate415(0x9, 0898, 0416, 0897);
  lut lut_gate416(0x9, 0924, 0899, 0898);
  lut lut_gate417(0x9, 0900, 0417, 0899);
  lut lut_gate418(0x9, 0923, 0901, 0900);
  lut lut_gate419(0x9, 0903, 0418, 0901);
  lut lut_gate420(0x9, 0922, 0904, 0903);
  lut lut_gate421(0x9, 0905, 0419, 0904);
  lut lut_gate422(0x9, 0921, 0906, 0905);
  lut lut_gate423(0x9, 0907, 0420, 0906);
  lut lut_gate424(0x9, 0920, 0908, 0907);
  lut lut_gate425(0x9, 0909, 0422, 0908);
  lut lut_gate426(0x9, 0919, 0910, 0909);
  lut lut_gate427(0x9, 0911, 0423, 0910);
  lut lut_gate428(0x9, 0918, 0912, 0911);
  lut lut_gate429(0x9, 0913, 0424, 0912);
  lut lut_gate430(0x9, 0917, 0914, 0913);
  lut lut_gate431(0x6, 0915, 0425, 0914);
  lut lut_gate432(0x8, G19, G16, 0915);
  lut lut_gate433(0x8, G20, G15, 0917);
  lut lut_gate434(0x8, G21, G14, 0918);
  lut lut_gate435(0x8, G22, G13, 0919);
  lut lut_gate436(0x8, G12, G23, 0920);
  lut lut_gate437(0x8, G11, G24, 0921);
  lut lut_gate438(0x8, G25, G10, 0922);
  lut lut_gate439(0x8, G26, G9, 0923);
  lut lut_gate440(0x8, G27, G8, 0924);
  lut lut_gate441(0x8, G7, G28, 0925);
  lut lut_gate442(0x8, G6, G29, 0926);
  lut lut_gate443(0x8, G5, G30, 0927);
  lut lut_gate444(0x8, G4, G31, 0928);
  lut lut_gate445(0x8, G3, G32, 0929);
  lut lut_gate446(0x9, 0931, 0426, 0930);
  lut lut_gate447(0x9, 0970, 0932, 0931);
  lut lut_gate448(0x9, 0933, 0427, 0932);
  lut lut_gate449(0x9, 0968, 0934, 0933);
  lut lut_gate450(0x9, 0935, 0428, 0934);
  lut lut_gate451(0x9, 0967, 0936, 0935);
  lut lut_gate452(0x9, 0938, 0429, 0936);
  lut lut_gate453(0x9, 0966, 0939, 0938);
  lut lut_gate454(0x9, 0940, 0430, 0939);
  lut lut_gate455(0x9, 0965, 0941, 0940);
  lut lut_gate456(0x9, 0942, 0431, 0941);
  lut lut_gate457(0x9, 0964, 0943, 0942);
  lut lut_gate458(0x9, 0944, 0433, 0943);
  lut lut_gate459(0x9, 0963, 0945, 0944);
  lut lut_gate460(0x9, 0946, 0434, 0945);
  lut lut_gate461(0x9, 0962, 0947, 0946);
  lut lut_gate462(0x9, 0948, 0435, 0947);
  lut lut_gate463(0x9, 0961, 0949, 0948);
  lut lut_gate464(0x9, 0951, 0436, 0949);
  lut lut_gate465(0x9, 0960, 0952, 0951);
  lut lut_gate466(0x9, 0953, 0437, 0952);
  lut lut_gate467(0x9, 0959, 0954, 0953);
  lut lut_gate468(0x9, 0955, 0438, 0954);
  lut lut_gate469(0x9, 0958, 0956, 0955);
  lut lut_gate470(0x6, 0957, 0439, 0956);
  lut lut_gate471(0x8, G20, G16, 0957);
  lut lut_gate472(0x8, G21, G15, 0958);
  lut lut_gate473(0x8, G22, G14, 0959);
  lut lut_gate474(0x8, G13, G23, 0960);
  lut lut_gate475(0x8, G12, G24, 0961);
  lut lut_gate476(0x8, G11, G25, 0962);
  lut lut_gate477(0x8, G26, G10, 0963);
  lut lut_gate478(0x8, G27, G9, 0964);
  lut lut_gate479(0x8, G8, G28, 0965);
  lut lut_gate480(0x8, G7, G29, 0966);
  lut lut_gate481(0x8, G6, G30, 0967);
  lut lut_gate482(0x8, G5, G31, 0968);
  lut lut_gate483(0x8, G4, G32, 0970);
  lut lut_gate484(0x9, 0972, 0440, 0971);
  lut lut_gate485(0x9, 0080, 0973, 0972);
  lut lut_gate486(0x9, 0974, 0441, 0973);
  lut lut_gate487(0x9, 0079, 0975, 0974);
  lut lut_gate488(0x9, 0976, 0442, 0975);
  lut lut_gate489(0x9, 0078, 0977, 0976);
  lut lut_gate490(0x9, 0978, 0444, 0977);
  lut lut_gate491(0x9, 0077, 0979, 0978);
  lut lut_gate492(0x9, 0980, 0445, 0979);
  lut lut_gate493(0x9, 0076, 0981, 0980);
  lut lut_gate494(0x9, 0983, 0446, 0981);
  lut lut_gate495(0x9, 0075, 0984, 0983);
  lut lut_gate496(0x9, 0985, 0447, 0984);
  lut lut_gate497(0x9, 0074, 0986, 0985);
  lut lut_gate498(0x9, 0987, 0448, 0986);
  lut lut_gate499(0x9, 0073, 0988, 0987);
  lut lut_gate500(0x9, 0989, 0449, 0988);
  lut lut_gate501(0x9, 0072, 0990, 0989);
  lut lut_gate502(0x9, 0064, 0450, 0990);
  lut lut_gate503(0x9, 0071, 0065, 0064);
  lut lut_gate504(0x9, 0066, 0451, 0065);
  lut lut_gate505(0x9, 0070, 0067, 0066);
  lut lut_gate506(0x6, 0069, 0452, 0067);
  lut lut_gate507(0x8, G21, G16, 0069);
  lut lut_gate508(0x8, G22, G15, 0070);
  lut lut_gate509(0x8, G14, G23, 0071);
  lut lut_gate510(0x8, G13, G24, 0072);
  lut lut_gate511(0x8, G12, G25, 0073);
  lut lut_gate512(0x8, G11, G26, 0074);
  lut lut_gate513(0x8, G27, G10, 0075);
  lut lut_gate514(0x8, G9, G28, 0076);
  lut lut_gate515(0x8, G8, G29, 0077);
  lut lut_gate516(0x8, G7, G30, 0078);
  lut lut_gate517(0x8, G6, G31, 0079);
  lut lut_gate518(0x8, G5, G32, 0080);
  lut lut_gate519(0x9, 0082, 0453, 0081);
  lut lut_gate520(0x9, 0114, 0083, 0082);
  lut lut_gate521(0x9, 0084, 0455, 0083);
  lut lut_gate522(0x9, 0113, 0085, 0084);
  lut lut_gate523(0x9, 0086, 0456, 0085);
  lut lut_gate524(0x9, 0112, 0087, 0086);
  lut lut_gate525(0x9, 0089, 0457, 0087);
  lut lut_gate526(0x9, 0111, 0090, 0089);
  lut lut_gate527(0x9, 0091, 0458, 0090);
  lut lut_gate528(0x9, 0110, 0092, 0091);
  lut lut_gate529(0x9, 0093, 0459, 0092);
  lut lut_gate530(0x9, 0109, 0094, 0093);
  lut lut_gate531(0x9, 0095, 0460, 0094);
  lut lut_gate532(0x9, 0108, 0096, 0095);
  lut lut_gate533(0x9, 0097, 0461, 0096);
  lut lut_gate534(0x9, 0107, 0098, 0097);
  lut lut_gate535(0x9, 0099, 0462, 0098);
  lut lut_gate536(0x9, 0106, 0100, 0099);
  lut lut_gate537(0x9, 0102, 0463, 0100);
  lut lut_gate538(0x9, 0105, 0103, 0102);
  lut lut_gate539(0x6, 0104, 0464, 0103);
  lut lut_gate540(0x8, G22, G16, 0104);
  lut lut_gate541(0x8, G15, G23, 0105);
  lut lut_gate542(0x8, G14, G24, 0106);
  lut lut_gate543(0x8, G13, G25, 0107);
  lut lut_gate544(0x8, G12, G26, 0108);
  lut lut_gate545(0x8, G11, G27, 0109);
  lut lut_gate546(0x8, G28, G10, 0110);
  lut lut_gate547(0x8, G29, G9, 0111);
  lut lut_gate548(0x8, G30, G8, 0112);
  lut lut_gate549(0x8, G31, G7, 0113);
  lut lut_gate550(0x8, G32, G6, 0114);
  lut lut_gate551(0x6, 0115, 0466, G6278);
  lut lut_gate552(0x9, 0116, 0467, 0115);
  lut lut_gate553(0x9, 0145, 0117, 0116);
  lut lut_gate554(0x9, 0119, 0468, 0117);
  lut lut_gate555(0x9, 0144, 0120, 0119);
  lut lut_gate556(0x9, 0121, 0469, 0120);
  lut lut_gate557(0x9, 0143, 0122, 0121);
  lut lut_gate558(0x9, 0123, 0470, 0122);
  lut lut_gate559(0x9, 0142, 0124, 0123);
  lut lut_gate560(0x9, 0125, 0471, 0124);
  lut lut_gate561(0x9, 0141, 0126, 0125);
  lut lut_gate562(0x9, 0127, 0472, 0126);
  lut lut_gate563(0x9, 0140, 0128, 0127);
  lut lut_gate564(0x9, 0129, 0473, 0128);
  lut lut_gate565(0x9, 0139, 0130, 0129);
  lut lut_gate566(0x9, 0132, 0474, 0130);
  lut lut_gate567(0x9, 0138, 0133, 0132);
  lut lut_gate568(0x9, 0134, 0475, 0133);
  lut lut_gate569(0x9, 0137, 0135, 0134);
  lut lut_gate570(0x6, 0136, 0477, 0135);
  lut lut_gate571(0x8, G23, G16, 0136);
  lut lut_gate572(0x8, G24, G15, 0137);
  lut lut_gate573(0x8, G25, G14, 0138);
  lut lut_gate574(0x8, G26, G13, 0139);
  lut lut_gate575(0x8, G27, G12, 0140);
  lut lut_gate576(0x8, G11, G28, 0141);
  lut lut_gate577(0x8, G29, G10, 0142);
  lut lut_gate578(0x8, G30, G9, 0143);
  lut lut_gate579(0x8, G31, G8, 0144);
  lut lut_gate580(0x8, G32, G7, 0145);
  lut lut_gate581(0x6, 0146, 0478, G6279);
  lut lut_gate582(0x9, 0148, 0479, 0146);
  lut lut_gate583(0x9, 0176, 0149, 0148);
  lut lut_gate584(0x9, 0150, 0480, 0149);
  lut lut_gate585(0x9, 0175, 0151, 0150);
  lut lut_gate586(0x9, 0153, 0481, 0151);
  lut lut_gate587(0x9, 0174, 0154, 0153);
  lut lut_gate588(0x9, 0155, 0482, 0154);
  lut lut_gate589(0x9, 0173, 0156, 0155);
  lut lut_gate590(0x9, 0158, 0483, 0156);
  lut lut_gate591(0x9, 0172, 0159, 0158);
  lut lut_gate592(0x9, 0160, 0484, 0159);
  lut lut_gate593(0x9, 0171, 0161, 0160);
  lut lut_gate594(0x9, 0163, 0485, 0161);
  lut lut_gate595(0x9, 0170, 0164, 0163);
  lut lut_gate596(0x9, 0165, 0486, 0164);
  lut lut_gate597(0x9, 0169, 0166, 0165);
  lut lut_gate598(0x6, 0168, 0488, 0166);
  lut lut_gate599(0x8, G24, G16, 0168);
  lut lut_gate600(0x8, G25, G15, 0169);
  lut lut_gate601(0x8, G26, G14, 0170);
  lut lut_gate602(0x8, G27, G13, 0171);
  lut lut_gate603(0x8, G12, G28, 0172);
  lut lut_gate604(0x8, G11, G29, 0173);
  lut lut_gate605(0x8, G30, G10, 0174);
  lut lut_gate606(0x8, G31, G9, 0175);
  lut lut_gate607(0x8, G32, G8, 0176);
  lut lut_gate608(0x6, 0178, 0489, G6280);
  lut lut_gate609(0x9, 0179, 0490, 0178);
  lut lut_gate610(0x9, 0203, 0180, 0179);
  lut lut_gate611(0x9, 0182, 0491, 0180);
  lut lut_gate612(0x9, 0202, 0183, 0182);
  lut lut_gate613(0x9, 0184, 0492, 0183);
  lut lut_gate614(0x9, 0201, 0185, 0184);
  lut lut_gate615(0x9, 0187, 0493, 0185);
  lut lut_gate616(0x9, 0200, 0188, 0187);
  lut lut_gate617(0x9, 0189, 0494, 0188);
  lut lut_gate618(0x9, 0199, 0190, 0189);
  lut lut_gate619(0x9, 0191, 0495, 0190);
  lut lut_gate620(0x9, 0198, 0192, 0191);
  lut lut_gate621(0x9, 0193, 0496, 0192);
  lut lut_gate622(0x9, 0197, 0194, 0193);
  lut lut_gate623(0x6, 0196, 0497, 0194);
  lut lut_gate624(0x8, G25, G16, 0196);
  lut lut_gate625(0x8, G26, G15, 0197);
  lut lut_gate626(0x8, G27, G14, 0198);
  lut lut_gate627(0x8, G13, G28, 0199);
  lut lut_gate628(0x8, G12, G29, 0200);
  lut lut_gate629(0x8, G11, G30, 0201);
  lut lut_gate630(0x8, G31, G10, 0202);
  lut lut_gate631(0x8, G32, G9, 0203);
  lut lut_gate632(0x6, 0205, 0499, G6281);
  lut lut_gate633(0x9, 0206, 0500, 0205);
  lut lut_gate634(0x9, 0228, 0207, 0206);
  lut lut_gate635(0x9, 0209, 0501, 0207);
  lut lut_gate636(0x9, 0227, 0210, 0209);
  lut lut_gate637(0x9, 0211, 0502, 0210);
  lut lut_gate638(0x9, 0226, 0212, 0211);
  lut lut_gate639(0x9, 0214, 0503, 0212);
  lut lut_gate640(0x9, 0225, 0215, 0214);
  lut lut_gate641(0x9, 0216, 0504, 0215);
  lut lut_gate642(0x9, 0224, 0217, 0216);
  lut lut_gate643(0x9, 0219, 0505, 0217);
  lut lut_gate644(0x9, 0222, 0220, 0219);
  lut lut_gate645(0x6, 0221, 0506, 0220);
  lut lut_gate646(0x8, G26, G16, 0221);
  lut lut_gate647(0x8, G27, G15, 0222);
  lut lut_gate648(0x8, G14, G28, 0224);
  lut lut_gate649(0x8, G13, G29, 0225);
  lut lut_gate650(0x8, G12, G30, 0226);
  lut lut_gate651(0x8, G11, G31, 0227);
  lut lut_gate652(0x8, G32, G10, 0228);
  lut lut_gate653(0x6, 0229, 0507, G6282);
  lut lut_gate654(0x9, 0231, 0508, 0229);
  lut lut_gate655(0x9, 0248, 0232, 0231);
  lut lut_gate656(0x9, 0233, 0510, 0232);
  lut lut_gate657(0x9, 0247, 0234, 0233);
  lut lut_gate658(0x9, 0236, 0511, 0234);
  lut lut_gate659(0x9, 0246, 0237, 0236);
  lut lut_gate660(0x9, 0238, 0512, 0237);
  lut lut_gate661(0x9, 0245, 0239, 0238);
  lut lut_gate662(0x9, 0240, 0513, 0239);
  lut lut_gate663(0x9, 0243, 0241, 0240);
  lut lut_gate664(0x6, 0242, 0514, 0241);
  lut lut_gate665(0x8, G27, G16, 0242);
  lut lut_gate666(0x8, G15, G28, 0243);
  lut lut_gate667(0x8, G14, G29, 0245);
  lut lut_gate668(0x8, G13, G30, 0246);
  lut lut_gate669(0x8, G12, G31, 0247);
  lut lut_gate670(0x8, G11, G32, 0248);
  lut lut_gate671(0x6, 0249, 0515, G6283);
  lut lut_gate672(0x9, 0251, 0516, 0249);
  lut lut_gate673(0x9, 0263, 0252, 0251);
  lut lut_gate674(0x9, 0253, 0517, 0252);
  lut lut_gate675(0x9, 0262, 0254, 0253);
  lut lut_gate676(0x9, 0255, 0518, 0254);
  lut lut_gate677(0x9, 0261, 0256, 0255);
  lut lut_gate678(0x9, 0257, 0519, 0256);
  lut lut_gate679(0x9, 0260, 0258, 0257);
  lut lut_gate680(0x6, 0259, 0521, 0258);
  lut lut_gate681(0x8, G16, G28, 0259);
  lut lut_gate682(0x8, G15, G29, 0260);
  lut lut_gate683(0x8, G14, G30, 0261);
  lut lut_gate684(0x8, G13, G31, 0262);
  lut lut_gate685(0x8, G12, G32, 0263);
  lut lut_gate686(0x6, 0264, 0522, G6284);
  lut lut_gate687(0x9, 0265, 0523, 0264);
  lut lut_gate688(0x9, 0276, 0266, 0265);
  lut lut_gate689(0x9, 0268, 0524, 0266);
  lut lut_gate690(0x9, 0275, 0269, 0268);
  lut lut_gate691(0x9, 0270, 0525, 0269);
  lut lut_gate692(0x9, 0274, 0271, 0270);
  lut lut_gate693(0x6, 0273, 0526, 0271);
  lut lut_gate694(0x8, G16, G29, 0273);
  lut lut_gate695(0x8, G15, G30, 0274);
  lut lut_gate696(0x8, G14, G31, 0275);
  lut lut_gate697(0x8, G13, G32, 0276);
  lut lut_gate698(0x6, 0277, 0527, G6285);
  lut lut_gate699(0x9, 0279, 0528, 0277);
  lut lut_gate700(0x9, 0286, 0280, 0279);
  lut lut_gate701(0x9, 0281, 0529, 0280);
  lut lut_gate702(0x9, 0285, 0282, 0281);
  lut lut_gate703(0x6, 0284, 0530, 0282);
  lut lut_gate704(0x8, G16, G30, 0284);
  lut lut_gate705(0x8, G15, G31, 0285);
  lut lut_gate706(0x8, G14, G32, 0286);
  lut lut_gate707(0x6, 0287, 0531, G6286);
  lut lut_gate708(0x9, 0289, 0532, 0287);
  lut lut_gate709(0x9, 0292, 0290, 0289);
  lut lut_gate710(0x6, 0291, 0533, 0290);
  lut lut_gate711(0x8, G16, G31, 0291);
  lut lut_gate712(0x8, G15, G32, 0292);
  lut lut_gate713(0x6, 0295, 0535, 0294);
  lut lut_gate714(0x8, G16, G32, 0295);
  lut lut_gate715(0x6, 0294, 0534, G6288);
  lut lut_gate716(0x9, 0841, 0302, G6273);
  lut lut_gate717(0x8, G1, G17, G6257);
  lut lut_gate718(0x6, 0186, 0147, G6259);
  lut lut_gate719(0x6, 0162, 0157, G6258);
  lut lut_gate720(0x6, 0235, 0131, G6260);
  lut lut_gate721(0x6, 0298, 0118, G6261);
  lut lut_gate722(0x6, 0520, 0101, G6262);
  lut lut_gate723(0x6, 0552, 0088, G6263);
  lut lut_gate724(0x6, 0572, 0068, G6264);
  lut lut_gate725(0x6, 0595, 0982, G6265);
  lut lut_gate726(0x6, 0621, 0969, G6266);
  lut lut_gate727(0x6, 0650, 0950, G6267);
  lut lut_gate728(0x6, 0682, 0937, G6268);
  lut lut_gate729(0x6, 0717, 0916, G6269);
  lut lut_gate730(0x6, 0755, 0902, G6270);
  lut lut_gate731(0x6, 0796, 0889, G6271);
  lut lut_gate732(0x6, 0840, 0867, G6272);
  lut lut_gate733(0x6, 0886, 0854, G6274);
  lut lut_gate734(0x6, 0930, 0301, G6275);
  lut lut_gate735(0x6, 0971, 0300, G6276);
  lut lut_gate736(0xb2, 0440, 0972, 0300, 0299);
  lut lut_gate737(0xb2, 0426, 0931, 0301, 0300);
  lut lut_gate738(0xb2, 0411, 0887, 0854, 0301);
  lut lut_gate739(0xb2, 0840, 0797, 0303, 0302);
  lut lut_gate740(0xb2, 0796, 0756, 0304, 0303);
  lut lut_gate741(0xb2, 0755, 0718, 0305, 0304);
  lut lut_gate742(0xb2, 0717, 0683, 0306, 0305);
  lut lut_gate743(0xb2, 0682, 0651, 0307, 0306);
  lut lut_gate744(0xb2, 0650, 0622, 0308, 0307);
  lut lut_gate745(0xb2, 0621, 0596, 0309, 0308);
  lut lut_gate746(0xb2, 0595, 0573, 0310, 0309);
  lut lut_gate747(0xb2, 0572, 0553, 0311, 0310);
  lut lut_gate748(0xb2, 0552, 0536, 0312, 0311);
  lut lut_gate749(0xb2, 0520, 0317, 0313, 0312);
  lut lut_gate750(0xb2, 0298, 0244, 0314, 0313);
  lut lut_gate751(0xb2, 0235, 0195, 0315, 0314);
  lut lut_gate752(0xe8, 0186, 0167, 0152, 0315);
  lut lut_gate753(0xe8, 0230, 0213, 0208, 0316);
  lut lut_gate754(0x4, 0316, 0297, 0267, 0318);
  lut lut_gate755(0xe8, 0296, 0283, 0278, 0319);
  lut lut_gate756(0x4, 0318, 0509, 0369, 0320);
  lut lut_gate757(0x4, 0319, 0498, 0421, 0321);
  lut lut_gate758(0xe8, 0487, 0454, 0443, 0322);
  lut lut_gate759(0x4, 0320, 0551, 0538, 0323);
  lut lut_gate760(0x4, 0321, 0550, 0540, 0324);
  lut lut_gate761(0x4, 0322, 0549, 0542, 0325);
  lut lut_gate762(0xe8, 0548, 0545, 0544, 0326);
  lut lut_gate763(0x4, 0323, 0571, 0555, 0327);
  lut lut_gate764(0x4, 0324, 0570, 0557, 0329);
  lut lut_gate765(0x4, 0325, 0569, 0559, 0330);
  lut lut_gate766(0x4, 0326, 0568, 0561, 0331);
  lut lut_gate767(0xe8, 0567, 0564, 0563, 0332);
  lut lut_gate768(0x4, 0327, 0594, 0575, 0333);
  lut lut_gate769(0x4, 0329, 0593, 0577, 0334);
  lut lut_gate770(0x4, 0330, 0592, 0579, 0335);
  lut lut_gate771(0x4, 0331, 0591, 0581, 0336);
  lut lut_gate772(0x4, 0332, 0590, 0583, 0337);
  lut lut_gate773(0xe8, 0589, 0586, 0585, 0338);
  lut lut_gate774(0x4, 0333, 0620, 0598, 0339);
  lut lut_gate775(0x4, 0334, 0619, 0600, 0340);
  lut lut_gate776(0x4, 0335, 0618, 0602, 0341);
  lut lut_gate777(0x4, 0336, 0617, 0604, 0342);
  lut lut_gate778(0x4, 0337, 0616, 0606, 0343);
  lut lut_gate779(0x4, 0338, 0615, 0608, 0344);
  lut lut_gate780(0xe8, 0614, 0611, 0610, 0345);
  lut lut_gate781(0x4, 0339, 0649, 0624, 0346);
  lut lut_gate782(0x4, 0340, 0648, 0626, 0347);
  lut lut_gate783(0x4, 0341, 0647, 0628, 0348);
  lut lut_gate784(0x4, 0342, 0646, 0630, 0349);
  lut lut_gate785(0x4, 0343, 0645, 0632, 0350);
  lut lut_gate786(0x4, 0344, 0644, 0634, 0351);
  lut lut_gate787(0x4, 0345, 0643, 0636, 0352);
  lut lut_gate788(0xe8, 0642, 0639, 0638, 0353);
  lut lut_gate789(0x4, 0346, 0681, 0653, 0354);
  lut lut_gate790(0x4, 0347, 0680, 0655, 0355);
  lut lut_gate791(0x4, 0348, 0679, 0657, 0356);
  lut lut_gate792(0x4, 0349, 0678, 0659, 0357);
  lut lut_gate793(0x4, 0350, 0677, 0661, 0358);
  lut lut_gate794(0x4, 0351, 0676, 0663, 0359);
  lut lut_gate795(0x4, 0352, 0675, 0665, 0360);
  lut lut_gate796(0x4, 0353, 0674, 0667, 0361);
  lut lut_gate797(0xe8, 0673, 0670, 0669, 0362);
  lut lut_gate798(0x4, 0354, 0716, 0685, 0363);
  lut lut_gate799(0x4, 0355, 0715, 0687, 0364);
  lut lut_gate800(0x4, 0356, 0714, 0689, 0365);
  lut lut_gate801(0x4, 0357, 0713, 0691, 0366);
  lut lut_gate802(0x4, 0358, 0712, 0693, 0367);
  lut lut_gate803(0x4, 0359, 0711, 0695, 0368);
  lut lut_gate804(0x4, 0360, 0710, 0697, 0370);
  lut lut_gate805(0x4, 0361, 0709, 0699, 0371);
  lut lut_gate806(0x4, 0362, 0708, 0701, 0372);
  lut lut_gate807(0xe8, 0707, 0704, 0703, 0373);
  lut lut_gate808(0x4, 0363, 0754, 0720, 0374);
  lut lut_gate809(0x4, 0364, 0753, 0722, 0375);
  lut lut_gate810(0x4, 0365, 0752, 0724, 0376);
  lut lut_gate811(0x4, 0366, 0751, 0726, 0377);
  lut lut_gate812(0x4, 0367, 0750, 0728, 0378);
  lut lut_gate813(0x4, 0368, 0749, 0730, 0379);
  lut lut_gate814(0x4, 0370, 0748, 0732, 0381);
  lut lut_gate815(0x4, 0371, 0747, 0734, 0382);
  lut lut_gate816(0x4, 0372, 0746, 0736, 0383);
  lut lut_gate817(0x4, 0373, 0745, 0738, 0384);
  lut lut_gate818(0xe8, 0744, 0741, 0740, 0385);
  lut lut_gate819(0x4, 0374, 0795, 0758, 0386);
  lut lut_gate820(0x4, 0375, 0794, 0760, 0387);
  lut lut_gate821(0x4, 0376, 0793, 0762, 0388);
  lut lut_gate822(0x4, 0377, 0792, 0764, 0389);
  lut lut_gate823(0x4, 0378, 0791, 0766, 0390);
  lut lut_gate824(0x4, 0379, 0790, 0768, 0391);
  lut lut_gate825(0x4, 0381, 0789, 0770, 0392);
  lut lut_gate826(0x4, 0382, 0788, 0772, 0393);
  lut lut_gate827(0x4, 0383, 0787, 0774, 0394);
  lut lut_gate828(0x4, 0384, 0786, 0776, 0395);
  lut lut_gate829(0x4, 0385, 0785, 0778, 0396);
  lut lut_gate830(0xe8, 0784, 0781, 0780, 0397);
  lut lut_gate831(0x4, 0386, 0839, 0799, 0398);
  lut lut_gate832(0x4, 0387, 0838, 0801, 0399);
  lut lut_gate833(0x4, 0388, 0837, 0803, 0400);
  lut lut_gate834(0x4, 0389, 0836, 0805, 0401);
  lut lut_gate835(0x4, 0390, 0835, 0807, 0402);
  lut lut_gate836(0x4, 0391, 0834, 0809, 0403);
  lut lut_gate837(0x4, 0392, 0833, 0811, 0404);
  lut lut_gate838(0x4, 0393, 0832, 0813, 0405);
  lut lut_gate839(0x4, 0394, 0831, 0815, 0406);
  lut lut_gate840(0x4, 0395, 0830, 0817, 0407);
  lut lut_gate841(0x4, 0396, 0829, 0819, 0408);
  lut lut_gate842(0x4, 0397, 0828, 0821, 0409);
  lut lut_gate843(0xe8, 0827, 0825, 0823, 0410);
  lut lut_gate844(0x4, 0398, 0885, 0843, 0411);
  lut lut_gate845(0x4, 0399, 0884, 0845, 0412);
  lut lut_gate846(0x4, 0400, 0883, 0847, 0413);
  lut lut_gate847(0x4, 0401, 0882, 0849, 0414);
  lut lut_gate848(0x4, 0402, 0881, 0851, 0415);
  lut lut_gate849(0x4, 0403, 0880, 0853, 0416);
  lut lut_gate850(0x4, 0404, 0879, 0856, 0417);
  lut lut_gate851(0x4, 0405, 0878, 0858, 0418);
  lut lut_gate852(0x4, 0406, 0877, 0860, 0419);
  lut lut_gate853(0x4, 0407, 0876, 0862, 0420);
  lut lut_gate854(0x4, 0408, 0875, 0864, 0422);
  lut lut_gate855(0x4, 0409, 0874, 0866, 0423);
  lut lut_gate856(0x4, 0410, 0873, 0869, 0424);
  lut lut_gate857(0xe0, 0871, 0783, 0872, 0425);
  lut lut_gate858(0x4, 0412, 0929, 0890, 0426);
  lut lut_gate859(0x4, 0413, 0928, 0892, 0427);
  lut lut_gate860(0x4, 0414, 0927, 0894, 0428);
  lut lut_gate861(0x4, 0415, 0926, 0896, 0429);
  lut lut_gate862(0x4, 0416, 0925, 0898, 0430);
  lut lut_gate863(0x4, 0417, 0924, 0900, 0431);
  lut lut_gate864(0x4, 0418, 0923, 0903, 0433);
  lut lut_gate865(0x4, 0419, 0922, 0905, 0434);
  lut lut_gate866(0x4, 0420, 0921, 0907, 0435);
  lut lut_gate867(0x4, 0422, 0920, 0909, 0436);
  lut lut_gate868(0x4, 0423, 0919, 0911, 0437);
  lut lut_gate869(0x4, 0424, 0918, 0913, 0438);
  lut lut_gate870(0xe8, 0425, 0917, 0915, 0439);
  lut lut_gate871(0x4, 0427, 0970, 0933, 0440);
  lut lut_gate872(0x4, 0428, 0968, 0935, 0441);
  lut lut_gate873(0x4, 0429, 0967, 0938, 0442);
  lut lut_gate874(0x4, 0430, 0966, 0940, 0444);
  lut lut_gate875(0x4, 0431, 0965, 0942, 0445);
  lut lut_gate876(0x4, 0433, 0964, 0944, 0446);
  lut lut_gate877(0x4, 0434, 0963, 0946, 0447);
  lut lut_gate878(0x4, 0435, 0962, 0948, 0448);
  lut lut_gate879(0x4, 0436, 0961, 0951, 0449);
  lut lut_gate880(0x4, 0437, 0960, 0953, 0450);
  lut lut_gate881(0x4, 0438, 0959, 0955, 0451);
  lut lut_gate882(0xe8, 0439, 0958, 0957, 0452);
  lut lut_gate883(0x4, 0441, 0080, 0974, 0453);
  lut lut_gate884(0x4, 0442, 0079, 0976, 0455);
  lut lut_gate885(0x4, 0444, 0078, 0978, 0456);
  lut lut_gate886(0x4, 0445, 0077, 0980, 0457);
  lut lut_gate887(0x4, 0446, 0076, 0983, 0458);
  lut lut_gate888(0x4, 0447, 0075, 0985, 0459);
  lut lut_gate889(0x4, 0448, 0074, 0987, 0460);
  lut lut_gate890(0x4, 0449, 0073, 0989, 0461);
  lut lut_gate891(0x4, 0450, 0072, 0064, 0462);
  lut lut_gate892(0x4, 0451, 0071, 0066, 0463);
  lut lut_gate893(0xe8, 0452, 0070, 0069, 0464);
  lut lut_gate894(0x4, 0453, 0299, 0082, 0466);
  lut lut_gate895(0x4, 0455, 0114, 0084, 0467);
  lut lut_gate896(0x4, 0456, 0113, 0086, 0468);
  lut lut_gate897(0x4, 0457, 0112, 0089, 0469);
  lut lut_gate898(0x4, 0458, 0111, 0091, 0470);
  lut lut_gate899(0x4, 0459, 0110, 0093, 0471);
  lut lut_gate900(0x4, 0460, 0109, 0095, 0472);
  lut lut_gate901(0x4, 0461, 0108, 0097, 0473);
  lut lut_gate902(0x4, 0462, 0107, 0099, 0474);
  lut lut_gate903(0x4, 0463, 0106, 0102, 0475);
  lut lut_gate904(0xe8, 0464, 0105, 0104, 0477);
  lut lut_gate905(0x4, 0467, 0466, 0116, 0478);
  lut lut_gate906(0x4, 0468, 0145, 0119, 0479);
  lut lut_gate907(0x4, 0469, 0144, 0121, 0480);
  lut lut_gate908(0x4, 0470, 0143, 0123, 0481);
  lut lut_gate909(0x4, 0471, 0142, 0125, 0482);
  lut lut_gate910(0x4, 0472, 0141, 0127, 0483);
  lut lut_gate911(0x4, 0473, 0140, 0129, 0484);
  lut lut_gate912(0x4, 0474, 0139, 0132, 0485);
  lut lut_gate913(0x4, 0475, 0138, 0134, 0486);
  lut lut_gate914(0xe8, 0477, 0137, 0136, 0488);
  lut lut_gate915(0x4, 0479, 0478, 0148, 0489);
  lut lut_gate916(0x4, 0480, 0176, 0150, 0490);
  lut lut_gate917(0x4, 0481, 0175, 0153, 0491);
  lut lut_gate918(0x4, 0482, 0174, 0155, 0492);
  lut lut_gate919(0x4, 0483, 0173, 0158, 0493);
  lut lut_gate920(0x4, 0484, 0172, 0160, 0494);
  lut lut_gate921(0x4, 0485, 0171, 0163, 0495);
  lut lut_gate922(0x4, 0486, 0170, 0165, 0496);
  lut lut_gate923(0xe8, 0488, 0169, 0168, 0497);
  lut lut_gate924(0x4, 0490, 0489, 0179, 0499);
  lut lut_gate925(0x4, 0491, 0203, 0182, 0500);
  lut lut_gate926(0x4, 0492, 0202, 0184, 0501);
  lut lut_gate927(0x4, 0493, 0201, 0187, 0502);
  lut lut_gate928(0x4, 0494, 0200, 0189, 0503);
  lut lut_gate929(0x4, 0495, 0199, 0191, 0504);
  lut lut_gate930(0x4, 0496, 0198, 0193, 0505);
  lut lut_gate931(0xe8, 0497, 0197, 0196, 0506);
  lut lut_gate932(0x4, 0500, 0499, 0206, 0507);
  lut lut_gate933(0x4, 0501, 0228, 0209, 0508);
  lut lut_gate934(0x4, 0502, 0227, 0211, 0510);
  lut lut_gate935(0x4, 0503, 0226, 0214, 0511);
  lut lut_gate936(0x4, 0504, 0225, 0216, 0512);
  lut lut_gate937(0x4, 0505, 0224, 0219, 0513);
  lut lut_gate938(0xe8, 0506, 0222, 0221, 0514);
  lut lut_gate939(0x4, 0508, 0507, 0231, 0515);
  lut lut_gate940(0x4, 0510, 0248, 0233, 0516);
  lut lut_gate941(0x4, 0511, 0247, 0236, 0517);
  lut lut_gate942(0x4, 0512, 0246, 0238, 0518);
  lut lut_gate943(0x4, 0513, 0245, 0240, 0519);
  lut lut_gate944(0xe8, 0514, 0243, 0242, 0521);
  lut lut_gate945(0x4, 0516, 0515, 0251, 0522);
  lut lut_gate946(0x4, 0517, 0263, 0253, 0523);
  lut lut_gate947(0x4, 0518, 0262, 0255, 0524);
  lut lut_gate948(0x4, 0519, 0261, 0257, 0525);
  lut lut_gate949(0xe8, 0521, 0260, 0259, 0526);
  lut lut_gate950(0x4, 0523, 0522, 0265, 0527);
  lut lut_gate951(0x4, 0524, 0276, 0268, 0528);
  lut lut_gate952(0x4, 0525, 0275, 0270, 0529);
  lut lut_gate953(0xe8, 0526, 0274, 0273, 0530);
  lut lut_gate954(0x4, 0528, 0527, 0279, 0531);
  lut lut_gate955(0x4, 0529, 0286, 0281, 0532);
  lut lut_gate956(0xe8, 0530, 0285, 0284, 0533);
  lut lut_gate957(0xe8, 0295, 0535, 0534, G6287);
  lut lut_gate958(0x4, 0532, 0531, 0289, 0534);
  lut lut_gate959(0xe8, 0533, 0292, 0291, 0535);

endmodule
