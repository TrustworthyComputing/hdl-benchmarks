module c880(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G7, G8, G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878, G879, G880, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, G293, G295, G296, G343, G349, G350, G369, G812, G829, G830, G831, G832, G844, G849, G850, G851;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G7, G8, G9;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878, G879, G880;
  lut lut_gate1(0x7f, G6, G16, G8, G855);
  lut lut_gate2(0x7f, G7, G17, G6, G856);
  lut lut_gate3(0x7f, G7, G6, G8, G857);
  lut lut_gate4(0x7, G18, G19, G858);
  lut lut_gate5(0x7fff, G1, G2, G3, G4, G859);
  lut lut_gate6(0x8, 378, G857, G860);
  lut lut_gate7(0x8000, G5, G1, G3, G4, 378);
  lut lut_gate8(0x1f, G23, G21, G20, G864);
  lut lut_gate9(0x4, 378, G857, G865);
  lut lut_gate10(0x7f, G9, G5, G1, G866);
  lut lut_gate11(0x1f, G22, G21, G20, G869);
  lut lut_gate12(0x0700, 308, 296, 297, G52, G872);
  lut lut_gate13(0x60, G51, G58, 297, 296);
  lut lut_gate14(0x9, G48, 298, 297);
  lut lut_gate15(0x4, 301, 299, 298);
  lut lut_gate16(0x40, 300, G10, G60, 299);
  lut lut_gate17(0x4000, G17, G6, G16, G866, 300);
  lut lut_gate18(0xb0bb, G31, 302, G39, 306, 301);
  lut lut_gate19(0xb0bb, 303, G866, 305, 304, 302);
  lut lut_gate20(0x6000, G11, G40, G4, G8, 303);
  lut lut_gate21(0x80, G11, G16, G8, 304);
  lut lut_gate22(0x8000, G9, G1, G2, G4, 305);
  lut lut_gate23(0xef00, G1, G4, G866, 307, 306);
  lut lut_gate24(0x8, G11, G40, 307);
  lut lut_gate25(0x0700, 310, 309, G30, G50, 308);
  lut lut_gate26(0x00f8, 298, G54, G53, G48, 309);
  lut lut_gate27(0x0777, G48, 311, G55, G59, 310);
  lut lut_gate28(0x80, G13, 313, 312, 311);
  lut lut_gate29(0x8000, G10, G1, G2, G3, 312);
  lut lut_gate30(0x8000, G14, G12, G11, G8, 313);
  lut lut_gate31(0x40, 329, 327, 314, G873);
  lut lut_gate32(0x9600, G51, G45, 325, 315, 314);
  lut lut_gate33(0x1, 320, 316, 315);
  lut lut_gate34(0x4, G46, 317, 316);
  lut lut_gate35(0x01, 319, 318, 299, 317);
  lut lut_gate36(0x4, G36, 306, 318);
  lut lut_gate37(0x4, G29, 302, 319);
  lut lut_gate38(0x00, 321, G47, 324, 322, 320);
  lut lut_gate39(0x0001, G46, 319, 318, 299, 321);
  lut lut_gate40(0x000, 323, 299, 306, G37, 322);
  lut lut_gate41(0x4, G30, 302, 323);
  lut lut_gate42(0xe8ee, 301, 299, G58, G48, 324);
  lut lut_gate43(0x0, 326, 306, G35, 325);
  lut lut_gate44(0x0, 299, 302, G28, 326);
  lut lut_gate45(0x70, 328, G50, G27, 327);
  lut lut_gate46(0x0bff, G45, 311, G53, 325, 328);
  lut lut_gate47(0x3f45, 325, G52, G45, G54, 329);
  lut lut_gate48(0x2b, G47, 324, 322, 330);
  lut lut_gate49(0x9, G46, 317, 331);
  lut lut_gate50(0x0, 333, 317, G54, 332);
  lut lut_gate51(0x70, 334, 311, G46, 333);
  lut lut_gate52(0x0777, G28, G50, G56, G55, 334);
  lut lut_gate53(0x0, 371, 335, 322, G54, G875);
  lut lut_gate54(0x60, G51, 324, 336, 335);
  lut lut_gate55(0x9, G47, 322, 336);
  lut lut_gate56(0x0777, G29, G50, G57, G55, 337);
  lut lut_gate57(0xb2, 350, G41, 338, G876);
  lut lut_gate58(0x222b, 347, 339, G42, 348, 338);
  lut lut_gate59(0x7100, 362, G44, 345, 340, 339);
  lut lut_gate60(0x222b, 316, 320, G45, 325, 340);
  lut lut_gate61(0x0, 343, 342, 302, G26, 341);
  lut lut_gate62(0x40, 300, G4, G60, 342);
  lut lut_gate63(0x0777, G37, 344, G34, G4, 343);
  lut lut_gate64(0x10, G10, 307, G866, 344);
  lut lut_gate65(0x0, 346, 342, 302, G27, 345);
  lut lut_gate66(0x0777, G39, 344, G38, G34, 346);
  lut lut_gate67(0x4, G43, 341, 347);
  lut lut_gate68(0x0, 349, 342, 302, G25, 348);
  lut lut_gate69(0x0777, G36, 344, G34, G9, 349);
  lut lut_gate70(0x0, 351, 342, 302, G24, 350);
  lut lut_gate71(0x0777, G35, 344, G34, G2, 351);
  lut lut_gate72(0x0700, 354, 352, 353, G52, G877);
  lut lut_gate73(0x90, G51, 353, 340, 352);
  lut lut_gate74(0x9, G44, 345, 353);
  lut lut_gate75(0x70, 355, 311, G44, 354);
  lut lut_gate76(0x07, 356, G50, G26, 355);
  lut lut_gate77(0x00f8, 345, G54, G44, G53, 356);
  lut lut_gate78(0x7, 373, 358, 338, G51, G878);
  lut lut_gate79(0x7077, G54, 350, G50, G60, 357);
  lut lut_gate80(0x9, G41, 350, 358);
  lut lut_gate81(0x7, 376, 360, 359, G51, G879);
  lut lut_gate82(0x1, 347, 339, 359);
  lut lut_gate83(0x9, G42, 348, 360);
  lut lut_gate84(0xb2, 345, G44, 340, 361);
  lut lut_gate85(0x9, G43, 341, 362);
  lut lut_gate86(0x0, 364, 341, G54, 363);
  lut lut_gate87(0x0777, G43, 311, G50, G25, 364);
  lut lut_gate88(0x80, G11, G17, G16, G861);
  lut lut_gate89(0x80, G11, G7, G17, G862);
  lut lut_gate90(0x80, G11, G7, G8, G863);
  lut lut_gate91(0x7f, G12, G6, 312, G867);
  lut lut_gate92(0x7fff, G15, G12, G11, 312, G868);
  lut lut_gate93(0x9669, G32, G26, G25, 365, G870);
  lut lut_gate94(0x9669, G33, G29, G28, 366, 365);
  lut lut_gate95(0x9669, G24, G27, G31, G30, 366);
  lut lut_gate96(0x6996, G32, G44, G43, 367, G871);
  lut lut_gate97(0x6996, G49, G47, G46, 368, 367);
  lut lut_gate98(0x9669, G42, G41, G45, G48, 368);
  lut lut_gate99(0x15cf, 331, G51, 330, G52, 369);
  lut lut_gate100(0x7000, 332, 369, G53, 316, G874);
  lut lut_gate101(0x35f3, G47, 322, G52, G53, 370);
  lut lut_gate102(0x7000, 337, 370, G47, 311, 371);
  lut lut_gate103(0x35f3, G41, 350, G52, G53, 372);
  lut lut_gate104(0x7000, 357, 372, G41, 311, 373);
  lut lut_gate105(0x0777, G24, G50, 311, G42, 374);
  lut lut_gate106(0x35f3, G42, 348, G52, G53, 375);
  lut lut_gate107(0xb000, 375, 374, G54, 348, 376);
  lut lut_gate108(0x15cf, 362, G51, 361, G52, 377);
  lut lut_gate109(0x7000, 363, 377, G53, 347, G880);

endmodule
