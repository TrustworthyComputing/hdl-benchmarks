module c499(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491, G492, G493, G494, G495, G496, G497, G498, G499, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491, G492, G493, G494, G495, G496, G497, G498, G499;
  lut lut_gate1(0x6, G1, 281, G468);
  lut lut_gate2(0x1000, 293, 282, 301, 300, 281);
  lut lut_gate3(0x4, 288, 283, 282);
  lut lut_gate4(0x9669, 287, 286, 285, 284, 283);
  lut lut_gate5(0x7887, G25, G29, G37, G41, 284);
  lut lut_gate6(0x9, G21, G17, 285);
  lut lut_gate7(0x9669, G7, G8, G6, G5, 286);
  lut lut_gate8(0x9669, G3, G4, G2, G1, 287);
  lut lut_gate9(0x9669, 292, 291, 290, 289, 288);
  lut lut_gate10(0x7887, G26, G30, G38, G41, 289);
  lut lut_gate11(0x9, G22, G18, 290);
  lut lut_gate12(0x9669, G15, G16, G14, G13, 291);
  lut lut_gate13(0x9669, G11, G12, G10, G9, 292);
  lut lut_gate14(0x1, 297, 294, 293);
  lut lut_gate15(0x9669, 296, 295, 291, 286, 294);
  lut lut_gate16(0x8, G40, G41, 295);
  lut lut_gate17(0x9669, G28, G32, G24, G20, 296);
  lut lut_gate18(0x9669, 299, 298, 292, 287, 297);
  lut lut_gate19(0x7887, G27, G31, G39, G41, 298);
  lut lut_gate20(0x9, G23, G19, 299);
  lut lut_gate21(0x6bbf, 240, 232, 301, 237, 300);
  lut lut_gate22(0x9669, 231, 304, 303, 302, 301);
  lut lut_gate23(0x7887, G9, G13, G33, G41, 302);
  lut lut_gate24(0x9, G1, G5, 303);
  lut lut_gate25(0x9669, G23, G24, G21, G22, 304);
  lut lut_gate26(0x9669, G19, G20, G17, G18, 231);
  lut lut_gate27(0x9669, 236, 235, 234, 233, 232);
  lut lut_gate28(0x7887, G14, G10, G34, G41, 233);
  lut lut_gate29(0x9, G6, G2, 234);
  lut lut_gate30(0x9669, G32, G31, G30, G29, 235);
  lut lut_gate31(0x9669, G28, G27, G26, G25, 236);
  lut lut_gate32(0x9669, 239, 238, 235, 304, 237);
  lut lut_gate33(0x8, G36, G41, 238);
  lut lut_gate34(0x9669, G16, G12, G8, G4, 239);
  lut lut_gate35(0x9669, 242, 241, 236, 231, 240);
  lut lut_gate36(0x7887, G15, G11, G35, G41, 241);
  lut lut_gate37(0x9, G7, G3, 242);
  lut lut_gate38(0x6, G2, 243, G469);
  lut lut_gate39(0x1000, 293, 282, 232, 300, 243);
  lut lut_gate40(0x6, G3, 244, G470);
  lut lut_gate41(0x1000, 293, 282, 240, 300, 244);
  lut lut_gate42(0x6, G4, 245, G471);
  lut lut_gate43(0x4000, 237, 282, 293, 300, 245);
  lut lut_gate44(0x6, G5, 246, G472);
  lut lut_gate45(0x1000, 282, 247, 301, 300, 246);
  lut lut_gate46(0x8, 297, 294, 247);
  lut lut_gate47(0x6, G6, 248, G473);
  lut lut_gate48(0x1000, 282, 247, 232, 300, 248);
  lut lut_gate49(0x6, G7, 249, G474);
  lut lut_gate50(0x1000, 282, 247, 240, 300, 249);
  lut lut_gate51(0x6, G8, 250, G475);
  lut lut_gate52(0x4000, 237, 247, 282, 300, 250);
  lut lut_gate53(0x6, G9, 251, G476);
  lut lut_gate54(0x1000, 293, 252, 301, 300, 251);
  lut lut_gate55(0x4, 283, 288, 252);
  lut lut_gate56(0x6, G10, 253, G477);
  lut lut_gate57(0x1000, 293, 252, 232, 300, 253);
  lut lut_gate58(0x6, G11, 254, G478);
  lut lut_gate59(0x1000, 293, 252, 240, 300, 254);
  lut lut_gate60(0x6, G12, 255, G479);
  lut lut_gate61(0x4000, 237, 252, 293, 300, 255);
  lut lut_gate62(0x6, G13, 256, G480);
  lut lut_gate63(0x1000, 247, 252, 301, 300, 256);
  lut lut_gate64(0x6, G14, 257, G481);
  lut lut_gate65(0x1000, 247, 252, 232, 300, 257);
  lut lut_gate66(0x6, G15, 258, G482);
  lut lut_gate67(0x1000, 247, 252, 240, 300, 258);
  lut lut_gate68(0x6, G16, 259, G483);
  lut lut_gate69(0x4000, 237, 252, 247, 300, 259);
  lut lut_gate70(0x6, G17, 260, G484);
  lut lut_gate71(0x1000, 262, 261, 283, 263, 260);
  lut lut_gate72(0x4, 232, 301, 261);
  lut lut_gate73(0x1, 240, 237, 262);
  lut lut_gate74(0x6bbf, 297, 288, 283, 294, 263);
  lut lut_gate75(0x6, G18, 264, G485);
  lut lut_gate76(0x1000, 262, 261, 288, 263, 264);
  lut lut_gate77(0x6, G19, 265, G486);
  lut lut_gate78(0x1000, 262, 261, 297, 263, 265);
  lut lut_gate79(0x6, G20, 266, G487);
  lut lut_gate80(0x4000, 294, 261, 262, 263, 266);
  lut lut_gate81(0x6, G21, 267, G488);
  lut lut_gate82(0x1000, 268, 261, 283, 263, 267);
  lut lut_gate83(0x8, 240, 237, 268);
  lut lut_gate84(0x6, G22, 269, G489);
  lut lut_gate85(0x1000, 268, 261, 288, 263, 269);
  lut lut_gate86(0x6, G23, 270, G490);
  lut lut_gate87(0x1000, 268, 261, 297, 263, 270);
  lut lut_gate88(0x6, G24, 271, G491);
  lut lut_gate89(0x4000, 294, 261, 268, 263, 271);
  lut lut_gate90(0x6, G25, 272, G492);
  lut lut_gate91(0x1000, 262, 273, 283, 263, 272);
  lut lut_gate92(0x4, 301, 232, 273);
  lut lut_gate93(0x6, G26, 274, G493);
  lut lut_gate94(0x1000, 262, 273, 288, 263, 274);
  lut lut_gate95(0x6, G27, 275, G494);
  lut lut_gate96(0x1000, 262, 273, 297, 263, 275);
  lut lut_gate97(0x6, G28, 276, G495);
  lut lut_gate98(0x4000, 294, 273, 262, 263, 276);
  lut lut_gate99(0x6, G29, 277, G496);
  lut lut_gate100(0x1000, 268, 273, 283, 263, 277);
  lut lut_gate101(0x6, G30, 278, G497);
  lut lut_gate102(0x1000, 268, 273, 288, 263, 278);
  lut lut_gate103(0x6, G31, 279, G498);
  lut lut_gate104(0x1000, 268, 273, 297, 263, 279);
  lut lut_gate105(0x6, G32, 280, G499);
  lut lut_gate106(0x4000, 294, 273, 268, 263, 280);

endmodule
