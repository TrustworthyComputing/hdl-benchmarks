module c1908(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893, G1894, G1895, G1896, G1897, G1898, G1899, G19, G1900, G1901, G1902, G1903, G1904, G1905, G1906, G1907, G1908, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G4, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, G313, G314, G315, G316, G317, G318, G319, G320, G321, G322, G323, G324, G325, G326, G327, G328, G335, G338, G341, G344, G347, G350, G356, G359, G362, G368, G374, G377, G395, G398, G401, G404, G407, G410, G413, G416, G419, G425, G428, G431, G437, G440, G443, G446, G449, G452, G455, G458, G467, G470, G473, G476, G479, G482, G485, G488, G491, G494, G497, G500, G506, G509, G512, G515, G518, G521, G524, G527, G530, G715, G716, G718, G719, G720, G721, G723, G728, G772, G774, G776, G778, G780, G782, G784, G786, G787, G789, G790, G792, G795, G805, G807, G808;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G4, G5, G6, G7, G8, G9;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893, G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903, G1904, G1905, G1906, G1907, G1908;
  lut lut_gate1(0x4, 245, 295, 294);
  lut lut_gate2(0x1, 243, 296, 295);
  lut lut_gate3(0x8, 230, 286, 296);
  lut lut_gate4(0x6, 304, 298, 297);
  lut lut_gate5(0x9, 302, 299, 298);
  lut lut_gate6(0x9, G13, 300, 299);
  lut lut_gate7(0x8, G20, 301, 300);
  lut lut_gate8(0x1, G23, G33, 301);
  lut lut_gate9(0x6, G16, 303, 302);
  lut lut_gate10(0x9, G9, G14, 303);
  lut lut_gate11(0x6, G4, 305, 304);
  lut lut_gate12(0x9, G7, G10, 305);
  lut lut_gate13(0x4, G19, 307, 306);
  lut lut_gate14(0x1, G23, G31, 307);
  lut lut_gate15(0x6, 311, 309, 308);
  lut lut_gate16(0x6, G12, 310, 309);
  lut lut_gate17(0x8, G19, 301, 310);
  lut lut_gate18(0x9, 314, 312, 311);
  lut lut_gate19(0x9, G3, 313, 312);
  lut lut_gate20(0x6, G10, G15, 313);
  lut lut_gate21(0x9, G6, G8, 314);
  lut lut_gate22(0x6, 321, 316, 315);
  lut lut_gate23(0x6, 302, 317, 316);
  lut lut_gate24(0x6, 320, 318, 317);
  lut lut_gate25(0x8, G18, 319, 318);
  lut lut_gate26(0x1, G24, G33, 319);
  lut lut_gate27(0x9, G11, G15, 320);
  lut lut_gate28(0x6, G8, 322, 321);
  lut lut_gate29(0x6, G2, G5, 322);
  lut lut_gate30(0x6, 226, 221, 220);
  lut lut_gate31(0x9, 224, 222, 221);
  lut lut_gate32(0x9, G1, 223, 222);
  lut lut_gate33(0x8, G17, 319, 223);
  lut lut_gate34(0x6, G6, 225, 224);
  lut lut_gate35(0x6, G7, G5, 225);
  lut lut_gate36(0x9, 229, 227, 226);
  lut lut_gate37(0x6, G13, 228, 227);
  lut lut_gate38(0x9, G11, G12, 228);
  lut lut_gate39(0x9, G16, 313, 229);
  lut lut_gate40(0x9, 241, 231, 230);
  lut lut_gate41(0x4, 232, G31, 231);
  lut lut_gate42(0x6, 238, 233, 232);
  lut lut_gate43(0x9, 236, 234, 233);
  lut lut_gate44(0x9, 235, 224, 234);
  lut lut_gate45(0x6, G4, G8, 235);
  lut lut_gate46(0x6, G3, 237, 236);
  lut lut_gate47(0x6, G1, G2, 237);
  lut lut_gate48(0x9, 239, 229, 238);
  lut lut_gate49(0x9, G9, 240, 239);
  lut lut_gate50(0x4, G21, G33, 240);
  lut lut_gate51(0x4, G17, 242, 241);
  lut lut_gate52(0x1, G24, G31, 242);
  lut lut_gate53(0x4, 286, 244, 243);
  lut lut_gate54(0x4, G18, 242, 244);
  lut lut_gate55(0x4, 288, 246, 245);
  lut lut_gate56(0x4, 254, 247, 246);
  lut lut_gate57(0x9, G25, 248, 247);
  lut lut_gate58(0x4, 249, G31, 248);
  lut lut_gate59(0x9, 250, 226, 249);
  lut lut_gate60(0x9, 251, 236, 250);
  lut lut_gate61(0x6, 253, 252, 251);
  lut lut_gate62(0x4, G22, G33, 252);
  lut lut_gate63(0x9, G4, G14, 253);
  lut lut_gate64(0x4, G20, 307, 254);
  lut lut_gate65(0x1, G32, G33, 255);
  lut lut_gate66(0x4, G24, G23, 256);
  lut lut_gate67(0x9, G1, 294, G1884);
  lut lut_gate68(0x9, G2, 294, G1885);
  lut lut_gate69(0x9, G3, 294, G1886);
  lut lut_gate70(0x9, G4, 294, G1887);
  lut lut_gate71(0x9, G10, 257, G1888);
  lut lut_gate72(0x4, 258, 295, 257);
  lut lut_gate73(0x4, 290, 246, 258);
  lut lut_gate74(0x9, G15, 257, G1889);
  lut lut_gate75(0x9, G16, 257, G1890);
  lut lut_gate76(0x9, G5, 259, G1891);
  lut lut_gate77(0x8, 288, 260, 259);
  lut lut_gate78(0x4, 261, 295, 260);
  lut lut_gate79(0x8, 254, 247, 261);
  lut lut_gate80(0x9, G6, 259, G1892);
  lut lut_gate81(0x9, G7, 259, G1893);
  lut lut_gate82(0x9, G8, 259, G1894);
  lut lut_gate83(0x9, G9, 262, G1895);
  lut lut_gate84(0x8, 290, 260, 262);
  lut lut_gate85(0x9, G11, 263, G1896);
  lut lut_gate86(0x8, 264, 296, 263);
  lut lut_gate87(0x8, 244, 258, 264);
  lut lut_gate88(0x9, G12, 263, G1897);
  lut lut_gate89(0x9, G13, 263, G1898);
  lut lut_gate90(0x9, G14, 263, G1899);
  lut lut_gate91(0xb, 267, 265, G1900);
  lut lut_gate92(0x4, G32, 266, 265);
  lut lut_gate93(0x1, 257, 294, 266);
  lut lut_gate94(0x1, G33, 268, 267);
  lut lut_gate95(0x8, 269, 243, 268);
  lut lut_gate96(0x8, 270, 230, 269);
  lut lut_gate97(0x4, 247, 254, 270);
  lut lut_gate98(0x4, 272, 266, 271);
  lut lut_gate99(0x4, 241, G31, 272);
  lut lut_gate100(0x4, 273, 255, G1902);
  lut lut_gate101(0x6, 249, 274, 273);
  lut lut_gate102(0x4, G25, 266, 274);
  lut lut_gate103(0x1, 255, 275, G1903);
  lut lut_gate104(0x8, 266, 315, 275);
  lut lut_gate105(0x1, 255, 276, G1904);
  lut lut_gate106(0x4, 266, 308, 276);
  lut lut_gate107(0x1, 255, 277, G1905);
  lut lut_gate108(0x4, 266, 297, 277);
  lut lut_gate109(0x4, 278, 255, G1908);
  lut lut_gate110(0x8, 266, 220, 278);
  lut lut_gate111(0xb4, 233, G21, G33, 279);
  lut lut_gate112(0x3, 279, G33, G29, 280);
  lut lut_gate113(0x6, 294, 280, G1906);
  lut lut_gate114(0x4b, G27, 315, G31, 281);
  lut lut_gate115(0x1e, G28, 308, G31, 282);
  lut lut_gate116(0x1e, 306, 297, G31, 283);
  lut lut_gate117(0x8, 283, 282, 284);
  lut lut_gate118(0x4b, G26, 220, G31, 285);
  lut lut_gate119(0x80, 285, 284, 281, 286);
  lut lut_gate120(0x1f, G32, G31, G29, 287);
  lut lut_gate121(0x10, 287, 256, G33, 288);
  lut lut_gate122(0x1f, G32, G30, G31, 289);
  lut lut_gate123(0x10, 289, 256, G33, 290);
  lut lut_gate124(0x6, 226, 303, 291);
  lut lut_gate125(0xb4, 291, G22, G33, 292);
  lut lut_gate126(0x3, 292, G33, G30, 293);
  lut lut_gate127(0x6, 257, 293, G1907);
  lut lut_gate128(0x14, 271, 232, 255, G1901);

endmodule
