module image_blur (p_0_0, p_0_1, p_0_2, p_0_3, p_0_4, p_0_5, p_0_6, p_0_7, p_0_8, p_0_9, p_0_10, p_0_11, p_0_12, p_0_13, p_0_14, p_0_15, p_0_16, p_0_17, p_0_18, p_0_19, p_0_20, p_0_21, p_0_22, p_0_23, p_0_24, p_0_25, p_0_26, p_0_27, p_0_28, p_0_29, p_0_30, p_0_31, p_0_32, p_0_33, p_0_34, p_0_35, p_0_36, p_0_37, p_0_38, p_0_39, p_0_40, p_0_41, p_0_42, p_0_43, p_0_44, p_0_45, p_0_46, p_0_47, p_0_48, p_0_49, p_0_50, p_0_51, p_0_52, p_0_53, p_0_54, p_0_55, p_0_56, p_0_57, p_0_58, p_0_59, p_0_60, p_0_61, p_0_62, p_0_63, p_0_64, p_0_65, p_1_0, p_1_1, p_1_2, p_1_3, p_1_4, p_1_5, p_1_6, p_1_7, p_1_8, p_1_9, p_1_10, p_1_11, p_1_12, p_1_13, p_1_14, p_1_15, p_1_16, p_1_17, p_1_18, p_1_19, p_1_20, p_1_21, p_1_22, p_1_23, p_1_24, p_1_25, p_1_26, p_1_27, p_1_28, p_1_29, p_1_30, p_1_31, p_1_32, p_1_33, p_1_34, p_1_35, p_1_36, p_1_37, p_1_38, p_1_39, p_1_40, p_1_41, p_1_42, p_1_43, p_1_44, p_1_45, p_1_46, p_1_47, p_1_48, p_1_49, p_1_50, p_1_51, p_1_52, p_1_53, p_1_54, p_1_55, p_1_56, p_1_57, p_1_58, p_1_59, p_1_60, p_1_61, p_1_62, p_1_63, p_1_64, p_1_65, p_2_0, p_2_1, p_2_2, p_2_3, p_2_4, p_2_5, p_2_6, p_2_7, p_2_8, p_2_9, p_2_10, p_2_11, p_2_12, p_2_13, p_2_14, p_2_15, p_2_16, p_2_17, p_2_18, p_2_19, p_2_20, p_2_21, p_2_22, p_2_23, p_2_24, p_2_25, p_2_26, p_2_27, p_2_28, p_2_29, p_2_30, p_2_31, p_2_32, p_2_33, p_2_34, p_2_35, p_2_36, p_2_37, p_2_38, p_2_39, p_2_40, p_2_41, p_2_42, p_2_43, p_2_44, p_2_45, p_2_46, p_2_47, p_2_48, p_2_49, p_2_50, p_2_51, p_2_52, p_2_53, p_2_54, p_2_55, p_2_56, p_2_57, p_2_58, p_2_59, p_2_60, p_2_61, p_2_62, p_2_63, p_2_64, p_2_65, p_3_0, p_3_1, p_3_2, p_3_3, p_3_4, p_3_5, p_3_6, p_3_7, p_3_8, p_3_9, p_3_10, p_3_11, p_3_12, p_3_13, p_3_14, p_3_15, p_3_16, p_3_17, p_3_18, p_3_19, p_3_20, p_3_21, p_3_22, p_3_23, p_3_24, p_3_25, p_3_26, p_3_27, p_3_28, p_3_29, p_3_30, p_3_31, p_3_32, p_3_33, p_3_34, p_3_35, p_3_36, p_3_37, p_3_38, p_3_39, p_3_40, p_3_41, p_3_42, p_3_43, p_3_44, p_3_45, p_3_46, p_3_47, p_3_48, p_3_49, p_3_50, p_3_51, p_3_52, p_3_53, p_3_54, p_3_55, p_3_56, p_3_57, p_3_58, p_3_59, p_3_60, p_3_61, p_3_62, p_3_63, p_3_64, p_3_65, p_4_0, p_4_1, p_4_2, p_4_3, p_4_4, p_4_5, p_4_6, p_4_7, p_4_8, p_4_9, p_4_10, p_4_11, p_4_12, p_4_13, p_4_14, p_4_15, p_4_16, p_4_17, p_4_18, p_4_19, p_4_20, p_4_21, p_4_22, p_4_23, p_4_24, p_4_25, p_4_26, p_4_27, p_4_28, p_4_29, p_4_30, p_4_31, p_4_32, p_4_33, p_4_34, p_4_35, p_4_36, p_4_37, p_4_38, p_4_39, p_4_40, p_4_41, p_4_42, p_4_43, p_4_44, p_4_45, p_4_46, p_4_47, p_4_48, p_4_49, p_4_50, p_4_51, p_4_52, p_4_53, p_4_54, p_4_55, p_4_56, p_4_57, p_4_58, p_4_59, p_4_60, p_4_61, p_4_62, p_4_63, p_4_64, p_4_65, p_5_0, p_5_1, p_5_2, p_5_3, p_5_4, p_5_5, p_5_6, p_5_7, p_5_8, p_5_9, p_5_10, p_5_11, p_5_12, p_5_13, p_5_14, p_5_15, p_5_16, p_5_17, p_5_18, p_5_19, p_5_20, p_5_21, p_5_22, p_5_23, p_5_24, p_5_25, p_5_26, p_5_27, p_5_28, p_5_29, p_5_30, p_5_31, p_5_32, p_5_33, p_5_34, p_5_35, p_5_36, p_5_37, p_5_38, p_5_39, p_5_40, p_5_41, p_5_42, p_5_43, p_5_44, p_5_45, p_5_46, p_5_47, p_5_48, p_5_49, p_5_50, p_5_51, p_5_52, p_5_53, p_5_54, p_5_55, p_5_56, p_5_57, p_5_58, p_5_59, p_5_60, p_5_61, p_5_62, p_5_63, p_5_64, p_5_65, p_6_0, p_6_1, p_6_2, p_6_3, p_6_4, p_6_5, p_6_6, p_6_7, p_6_8, p_6_9, p_6_10, p_6_11, p_6_12, p_6_13, p_6_14, p_6_15, p_6_16, p_6_17, p_6_18, p_6_19, p_6_20, p_6_21, p_6_22, p_6_23, p_6_24, p_6_25, p_6_26, p_6_27, p_6_28, p_6_29, p_6_30, p_6_31, p_6_32, p_6_33, p_6_34, p_6_35, p_6_36, p_6_37, p_6_38, p_6_39, p_6_40, p_6_41, p_6_42, p_6_43, p_6_44, p_6_45, p_6_46, p_6_47, p_6_48, p_6_49, p_6_50, p_6_51, p_6_52, p_6_53, p_6_54, p_6_55, p_6_56, p_6_57, p_6_58, p_6_59, p_6_60, p_6_61, p_6_62, p_6_63, p_6_64, p_6_65, p_7_0, p_7_1, p_7_2, p_7_3, p_7_4, p_7_5, p_7_6, p_7_7, p_7_8, p_7_9, p_7_10, p_7_11, p_7_12, p_7_13, p_7_14, p_7_15, p_7_16, p_7_17, p_7_18, p_7_19, p_7_20, p_7_21, p_7_22, p_7_23, p_7_24, p_7_25, p_7_26, p_7_27, p_7_28, p_7_29, p_7_30, p_7_31, p_7_32, p_7_33, p_7_34, p_7_35, p_7_36, p_7_37, p_7_38, p_7_39, p_7_40, p_7_41, p_7_42, p_7_43, p_7_44, p_7_45, p_7_46, p_7_47, p_7_48, p_7_49, p_7_50, p_7_51, p_7_52, p_7_53, p_7_54, p_7_55, p_7_56, p_7_57, p_7_58, p_7_59, p_7_60, p_7_61, p_7_62, p_7_63, p_7_64, p_7_65, p_8_0, p_8_1, p_8_2, p_8_3, p_8_4, p_8_5, p_8_6, p_8_7, p_8_8, p_8_9, p_8_10, p_8_11, p_8_12, p_8_13, p_8_14, p_8_15, p_8_16, p_8_17, p_8_18, p_8_19, p_8_20, p_8_21, p_8_22, p_8_23, p_8_24, p_8_25, p_8_26, p_8_27, p_8_28, p_8_29, p_8_30, p_8_31, p_8_32, p_8_33, p_8_34, p_8_35, p_8_36, p_8_37, p_8_38, p_8_39, p_8_40, p_8_41, p_8_42, p_8_43, p_8_44, p_8_45, p_8_46, p_8_47, p_8_48, p_8_49, p_8_50, p_8_51, p_8_52, p_8_53, p_8_54, p_8_55, p_8_56, p_8_57, p_8_58, p_8_59, p_8_60, p_8_61, p_8_62, p_8_63, p_8_64, p_8_65, p_9_0, p_9_1, p_9_2, p_9_3, p_9_4, p_9_5, p_9_6, p_9_7, p_9_8, p_9_9, p_9_10, p_9_11, p_9_12, p_9_13, p_9_14, p_9_15, p_9_16, p_9_17, p_9_18, p_9_19, p_9_20, p_9_21, p_9_22, p_9_23, p_9_24, p_9_25, p_9_26, p_9_27, p_9_28, p_9_29, p_9_30, p_9_31, p_9_32, p_9_33, p_9_34, p_9_35, p_9_36, p_9_37, p_9_38, p_9_39, p_9_40, p_9_41, p_9_42, p_9_43, p_9_44, p_9_45, p_9_46, p_9_47, p_9_48, p_9_49, p_9_50, p_9_51, p_9_52, p_9_53, p_9_54, p_9_55, p_9_56, p_9_57, p_9_58, p_9_59, p_9_60, p_9_61, p_9_62, p_9_63, p_9_64, p_9_65, p_10_0, p_10_1, p_10_2, p_10_3, p_10_4, p_10_5, p_10_6, p_10_7, p_10_8, p_10_9, p_10_10, p_10_11, p_10_12, p_10_13, p_10_14, p_10_15, p_10_16, p_10_17, p_10_18, p_10_19, p_10_20, p_10_21, p_10_22, p_10_23, p_10_24, p_10_25, p_10_26, p_10_27, p_10_28, p_10_29, p_10_30, p_10_31, p_10_32, p_10_33, p_10_34, p_10_35, p_10_36, p_10_37, p_10_38, p_10_39, p_10_40, p_10_41, p_10_42, p_10_43, p_10_44, p_10_45, p_10_46, p_10_47, p_10_48, p_10_49, p_10_50, p_10_51, p_10_52, p_10_53, p_10_54, p_10_55, p_10_56, p_10_57, p_10_58, p_10_59, p_10_60, p_10_61, p_10_62, p_10_63, p_10_64, p_10_65, p_11_0, p_11_1, p_11_2, p_11_3, p_11_4, p_11_5, p_11_6, p_11_7, p_11_8, p_11_9, p_11_10, p_11_11, p_11_12, p_11_13, p_11_14, p_11_15, p_11_16, p_11_17, p_11_18, p_11_19, p_11_20, p_11_21, p_11_22, p_11_23, p_11_24, p_11_25, p_11_26, p_11_27, p_11_28, p_11_29, p_11_30, p_11_31, p_11_32, p_11_33, p_11_34, p_11_35, p_11_36, p_11_37, p_11_38, p_11_39, p_11_40, p_11_41, p_11_42, p_11_43, p_11_44, p_11_45, p_11_46, p_11_47, p_11_48, p_11_49, p_11_50, p_11_51, p_11_52, p_11_53, p_11_54, p_11_55, p_11_56, p_11_57, p_11_58, p_11_59, p_11_60, p_11_61, p_11_62, p_11_63, p_11_64, p_11_65, p_12_0, p_12_1, p_12_2, p_12_3, p_12_4, p_12_5, p_12_6, p_12_7, p_12_8, p_12_9, p_12_10, p_12_11, p_12_12, p_12_13, p_12_14, p_12_15, p_12_16, p_12_17, p_12_18, p_12_19, p_12_20, p_12_21, p_12_22, p_12_23, p_12_24, p_12_25, p_12_26, p_12_27, p_12_28, p_12_29, p_12_30, p_12_31, p_12_32, p_12_33, p_12_34, p_12_35, p_12_36, p_12_37, p_12_38, p_12_39, p_12_40, p_12_41, p_12_42, p_12_43, p_12_44, p_12_45, p_12_46, p_12_47, p_12_48, p_12_49, p_12_50, p_12_51, p_12_52, p_12_53, p_12_54, p_12_55, p_12_56, p_12_57, p_12_58, p_12_59, p_12_60, p_12_61, p_12_62, p_12_63, p_12_64, p_12_65, p_13_0, p_13_1, p_13_2, p_13_3, p_13_4, p_13_5, p_13_6, p_13_7, p_13_8, p_13_9, p_13_10, p_13_11, p_13_12, p_13_13, p_13_14, p_13_15, p_13_16, p_13_17, p_13_18, p_13_19, p_13_20, p_13_21, p_13_22, p_13_23, p_13_24, p_13_25, p_13_26, p_13_27, p_13_28, p_13_29, p_13_30, p_13_31, p_13_32, p_13_33, p_13_34, p_13_35, p_13_36, p_13_37, p_13_38, p_13_39, p_13_40, p_13_41, p_13_42, p_13_43, p_13_44, p_13_45, p_13_46, p_13_47, p_13_48, p_13_49, p_13_50, p_13_51, p_13_52, p_13_53, p_13_54, p_13_55, p_13_56, p_13_57, p_13_58, p_13_59, p_13_60, p_13_61, p_13_62, p_13_63, p_13_64, p_13_65, p_14_0, p_14_1, p_14_2, p_14_3, p_14_4, p_14_5, p_14_6, p_14_7, p_14_8, p_14_9, p_14_10, p_14_11, p_14_12, p_14_13, p_14_14, p_14_15, p_14_16, p_14_17, p_14_18, p_14_19, p_14_20, p_14_21, p_14_22, p_14_23, p_14_24, p_14_25, p_14_26, p_14_27, p_14_28, p_14_29, p_14_30, p_14_31, p_14_32, p_14_33, p_14_34, p_14_35, p_14_36, p_14_37, p_14_38, p_14_39, p_14_40, p_14_41, p_14_42, p_14_43, p_14_44, p_14_45, p_14_46, p_14_47, p_14_48, p_14_49, p_14_50, p_14_51, p_14_52, p_14_53, p_14_54, p_14_55, p_14_56, p_14_57, p_14_58, p_14_59, p_14_60, p_14_61, p_14_62, p_14_63, p_14_64, p_14_65, p_15_0, p_15_1, p_15_2, p_15_3, p_15_4, p_15_5, p_15_6, p_15_7, p_15_8, p_15_9, p_15_10, p_15_11, p_15_12, p_15_13, p_15_14, p_15_15, p_15_16, p_15_17, p_15_18, p_15_19, p_15_20, p_15_21, p_15_22, p_15_23, p_15_24, p_15_25, p_15_26, p_15_27, p_15_28, p_15_29, p_15_30, p_15_31, p_15_32, p_15_33, p_15_34, p_15_35, p_15_36, p_15_37, p_15_38, p_15_39, p_15_40, p_15_41, p_15_42, p_15_43, p_15_44, p_15_45, p_15_46, p_15_47, p_15_48, p_15_49, p_15_50, p_15_51, p_15_52, p_15_53, p_15_54, p_15_55, p_15_56, p_15_57, p_15_58, p_15_59, p_15_60, p_15_61, p_15_62, p_15_63, p_15_64, p_15_65, p_16_0, p_16_1, p_16_2, p_16_3, p_16_4, p_16_5, p_16_6, p_16_7, p_16_8, p_16_9, p_16_10, p_16_11, p_16_12, p_16_13, p_16_14, p_16_15, p_16_16, p_16_17, p_16_18, p_16_19, p_16_20, p_16_21, p_16_22, p_16_23, p_16_24, p_16_25, p_16_26, p_16_27, p_16_28, p_16_29, p_16_30, p_16_31, p_16_32, p_16_33, p_16_34, p_16_35, p_16_36, p_16_37, p_16_38, p_16_39, p_16_40, p_16_41, p_16_42, p_16_43, p_16_44, p_16_45, p_16_46, p_16_47, p_16_48, p_16_49, p_16_50, p_16_51, p_16_52, p_16_53, p_16_54, p_16_55, p_16_56, p_16_57, p_16_58, p_16_59, p_16_60, p_16_61, p_16_62, p_16_63, p_16_64, p_16_65, p_17_0, p_17_1, p_17_2, p_17_3, p_17_4, p_17_5, p_17_6, p_17_7, p_17_8, p_17_9, p_17_10, p_17_11, p_17_12, p_17_13, p_17_14, p_17_15, p_17_16, p_17_17, p_17_18, p_17_19, p_17_20, p_17_21, p_17_22, p_17_23, p_17_24, p_17_25, p_17_26, p_17_27, p_17_28, p_17_29, p_17_30, p_17_31, p_17_32, p_17_33, p_17_34, p_17_35, p_17_36, p_17_37, p_17_38, p_17_39, p_17_40, p_17_41, p_17_42, p_17_43, p_17_44, p_17_45, p_17_46, p_17_47, p_17_48, p_17_49, p_17_50, p_17_51, p_17_52, p_17_53, p_17_54, p_17_55, p_17_56, p_17_57, p_17_58, p_17_59, p_17_60, p_17_61, p_17_62, p_17_63, p_17_64, p_17_65, p_18_0, p_18_1, p_18_2, p_18_3, p_18_4, p_18_5, p_18_6, p_18_7, p_18_8, p_18_9, p_18_10, p_18_11, p_18_12, p_18_13, p_18_14, p_18_15, p_18_16, p_18_17, p_18_18, p_18_19, p_18_20, p_18_21, p_18_22, p_18_23, p_18_24, p_18_25, p_18_26, p_18_27, p_18_28, p_18_29, p_18_30, p_18_31, p_18_32, p_18_33, p_18_34, p_18_35, p_18_36, p_18_37, p_18_38, p_18_39, p_18_40, p_18_41, p_18_42, p_18_43, p_18_44, p_18_45, p_18_46, p_18_47, p_18_48, p_18_49, p_18_50, p_18_51, p_18_52, p_18_53, p_18_54, p_18_55, p_18_56, p_18_57, p_18_58, p_18_59, p_18_60, p_18_61, p_18_62, p_18_63, p_18_64, p_18_65, p_19_0, p_19_1, p_19_2, p_19_3, p_19_4, p_19_5, p_19_6, p_19_7, p_19_8, p_19_9, p_19_10, p_19_11, p_19_12, p_19_13, p_19_14, p_19_15, p_19_16, p_19_17, p_19_18, p_19_19, p_19_20, p_19_21, p_19_22, p_19_23, p_19_24, p_19_25, p_19_26, p_19_27, p_19_28, p_19_29, p_19_30, p_19_31, p_19_32, p_19_33, p_19_34, p_19_35, p_19_36, p_19_37, p_19_38, p_19_39, p_19_40, p_19_41, p_19_42, p_19_43, p_19_44, p_19_45, p_19_46, p_19_47, p_19_48, p_19_49, p_19_50, p_19_51, p_19_52, p_19_53, p_19_54, p_19_55, p_19_56, p_19_57, p_19_58, p_19_59, p_19_60, p_19_61, p_19_62, p_19_63, p_19_64, p_19_65, p_20_0, p_20_1, p_20_2, p_20_3, p_20_4, p_20_5, p_20_6, p_20_7, p_20_8, p_20_9, p_20_10, p_20_11, p_20_12, p_20_13, p_20_14, p_20_15, p_20_16, p_20_17, p_20_18, p_20_19, p_20_20, p_20_21, p_20_22, p_20_23, p_20_24, p_20_25, p_20_26, p_20_27, p_20_28, p_20_29, p_20_30, p_20_31, p_20_32, p_20_33, p_20_34, p_20_35, p_20_36, p_20_37, p_20_38, p_20_39, p_20_40, p_20_41, p_20_42, p_20_43, p_20_44, p_20_45, p_20_46, p_20_47, p_20_48, p_20_49, p_20_50, p_20_51, p_20_52, p_20_53, p_20_54, p_20_55, p_20_56, p_20_57, p_20_58, p_20_59, p_20_60, p_20_61, p_20_62, p_20_63, p_20_64, p_20_65, p_21_0, p_21_1, p_21_2, p_21_3, p_21_4, p_21_5, p_21_6, p_21_7, p_21_8, p_21_9, p_21_10, p_21_11, p_21_12, p_21_13, p_21_14, p_21_15, p_21_16, p_21_17, p_21_18, p_21_19, p_21_20, p_21_21, p_21_22, p_21_23, p_21_24, p_21_25, p_21_26, p_21_27, p_21_28, p_21_29, p_21_30, p_21_31, p_21_32, p_21_33, p_21_34, p_21_35, p_21_36, p_21_37, p_21_38, p_21_39, p_21_40, p_21_41, p_21_42, p_21_43, p_21_44, p_21_45, p_21_46, p_21_47, p_21_48, p_21_49, p_21_50, p_21_51, p_21_52, p_21_53, p_21_54, p_21_55, p_21_56, p_21_57, p_21_58, p_21_59, p_21_60, p_21_61, p_21_62, p_21_63, p_21_64, p_21_65, p_22_0, p_22_1, p_22_2, p_22_3, p_22_4, p_22_5, p_22_6, p_22_7, p_22_8, p_22_9, p_22_10, p_22_11, p_22_12, p_22_13, p_22_14, p_22_15, p_22_16, p_22_17, p_22_18, p_22_19, p_22_20, p_22_21, p_22_22, p_22_23, p_22_24, p_22_25, p_22_26, p_22_27, p_22_28, p_22_29, p_22_30, p_22_31, p_22_32, p_22_33, p_22_34, p_22_35, p_22_36, p_22_37, p_22_38, p_22_39, p_22_40, p_22_41, p_22_42, p_22_43, p_22_44, p_22_45, p_22_46, p_22_47, p_22_48, p_22_49, p_22_50, p_22_51, p_22_52, p_22_53, p_22_54, p_22_55, p_22_56, p_22_57, p_22_58, p_22_59, p_22_60, p_22_61, p_22_62, p_22_63, p_22_64, p_22_65, p_23_0, p_23_1, p_23_2, p_23_3, p_23_4, p_23_5, p_23_6, p_23_7, p_23_8, p_23_9, p_23_10, p_23_11, p_23_12, p_23_13, p_23_14, p_23_15, p_23_16, p_23_17, p_23_18, p_23_19, p_23_20, p_23_21, p_23_22, p_23_23, p_23_24, p_23_25, p_23_26, p_23_27, p_23_28, p_23_29, p_23_30, p_23_31, p_23_32, p_23_33, p_23_34, p_23_35, p_23_36, p_23_37, p_23_38, p_23_39, p_23_40, p_23_41, p_23_42, p_23_43, p_23_44, p_23_45, p_23_46, p_23_47, p_23_48, p_23_49, p_23_50, p_23_51, p_23_52, p_23_53, p_23_54, p_23_55, p_23_56, p_23_57, p_23_58, p_23_59, p_23_60, p_23_61, p_23_62, p_23_63, p_23_64, p_23_65, p_24_0, p_24_1, p_24_2, p_24_3, p_24_4, p_24_5, p_24_6, p_24_7, p_24_8, p_24_9, p_24_10, p_24_11, p_24_12, p_24_13, p_24_14, p_24_15, p_24_16, p_24_17, p_24_18, p_24_19, p_24_20, p_24_21, p_24_22, p_24_23, p_24_24, p_24_25, p_24_26, p_24_27, p_24_28, p_24_29, p_24_30, p_24_31, p_24_32, p_24_33, p_24_34, p_24_35, p_24_36, p_24_37, p_24_38, p_24_39, p_24_40, p_24_41, p_24_42, p_24_43, p_24_44, p_24_45, p_24_46, p_24_47, p_24_48, p_24_49, p_24_50, p_24_51, p_24_52, p_24_53, p_24_54, p_24_55, p_24_56, p_24_57, p_24_58, p_24_59, p_24_60, p_24_61, p_24_62, p_24_63, p_24_64, p_24_65, p_25_0, p_25_1, p_25_2, p_25_3, p_25_4, p_25_5, p_25_6, p_25_7, p_25_8, p_25_9, p_25_10, p_25_11, p_25_12, p_25_13, p_25_14, p_25_15, p_25_16, p_25_17, p_25_18, p_25_19, p_25_20, p_25_21, p_25_22, p_25_23, p_25_24, p_25_25, p_25_26, p_25_27, p_25_28, p_25_29, p_25_30, p_25_31, p_25_32, p_25_33, p_25_34, p_25_35, p_25_36, p_25_37, p_25_38, p_25_39, p_25_40, p_25_41, p_25_42, p_25_43, p_25_44, p_25_45, p_25_46, p_25_47, p_25_48, p_25_49, p_25_50, p_25_51, p_25_52, p_25_53, p_25_54, p_25_55, p_25_56, p_25_57, p_25_58, p_25_59, p_25_60, p_25_61, p_25_62, p_25_63, p_25_64, p_25_65, p_26_0, p_26_1, p_26_2, p_26_3, p_26_4, p_26_5, p_26_6, p_26_7, p_26_8, p_26_9, p_26_10, p_26_11, p_26_12, p_26_13, p_26_14, p_26_15, p_26_16, p_26_17, p_26_18, p_26_19, p_26_20, p_26_21, p_26_22, p_26_23, p_26_24, p_26_25, p_26_26, p_26_27, p_26_28, p_26_29, p_26_30, p_26_31, p_26_32, p_26_33, p_26_34, p_26_35, p_26_36, p_26_37, p_26_38, p_26_39, p_26_40, p_26_41, p_26_42, p_26_43, p_26_44, p_26_45, p_26_46, p_26_47, p_26_48, p_26_49, p_26_50, p_26_51, p_26_52, p_26_53, p_26_54, p_26_55, p_26_56, p_26_57, p_26_58, p_26_59, p_26_60, p_26_61, p_26_62, p_26_63, p_26_64, p_26_65, p_27_0, p_27_1, p_27_2, p_27_3, p_27_4, p_27_5, p_27_6, p_27_7, p_27_8, p_27_9, p_27_10, p_27_11, p_27_12, p_27_13, p_27_14, p_27_15, p_27_16, p_27_17, p_27_18, p_27_19, p_27_20, p_27_21, p_27_22, p_27_23, p_27_24, p_27_25, p_27_26, p_27_27, p_27_28, p_27_29, p_27_30, p_27_31, p_27_32, p_27_33, p_27_34, p_27_35, p_27_36, p_27_37, p_27_38, p_27_39, p_27_40, p_27_41, p_27_42, p_27_43, p_27_44, p_27_45, p_27_46, p_27_47, p_27_48, p_27_49, p_27_50, p_27_51, p_27_52, p_27_53, p_27_54, p_27_55, p_27_56, p_27_57, p_27_58, p_27_59, p_27_60, p_27_61, p_27_62, p_27_63, p_27_64, p_27_65, p_28_0, p_28_1, p_28_2, p_28_3, p_28_4, p_28_5, p_28_6, p_28_7, p_28_8, p_28_9, p_28_10, p_28_11, p_28_12, p_28_13, p_28_14, p_28_15, p_28_16, p_28_17, p_28_18, p_28_19, p_28_20, p_28_21, p_28_22, p_28_23, p_28_24, p_28_25, p_28_26, p_28_27, p_28_28, p_28_29, p_28_30, p_28_31, p_28_32, p_28_33, p_28_34, p_28_35, p_28_36, p_28_37, p_28_38, p_28_39, p_28_40, p_28_41, p_28_42, p_28_43, p_28_44, p_28_45, p_28_46, p_28_47, p_28_48, p_28_49, p_28_50, p_28_51, p_28_52, p_28_53, p_28_54, p_28_55, p_28_56, p_28_57, p_28_58, p_28_59, p_28_60, p_28_61, p_28_62, p_28_63, p_28_64, p_28_65, p_29_0, p_29_1, p_29_2, p_29_3, p_29_4, p_29_5, p_29_6, p_29_7, p_29_8, p_29_9, p_29_10, p_29_11, p_29_12, p_29_13, p_29_14, p_29_15, p_29_16, p_29_17, p_29_18, p_29_19, p_29_20, p_29_21, p_29_22, p_29_23, p_29_24, p_29_25, p_29_26, p_29_27, p_29_28, p_29_29, p_29_30, p_29_31, p_29_32, p_29_33, p_29_34, p_29_35, p_29_36, p_29_37, p_29_38, p_29_39, p_29_40, p_29_41, p_29_42, p_29_43, p_29_44, p_29_45, p_29_46, p_29_47, p_29_48, p_29_49, p_29_50, p_29_51, p_29_52, p_29_53, p_29_54, p_29_55, p_29_56, p_29_57, p_29_58, p_29_59, p_29_60, p_29_61, p_29_62, p_29_63, p_29_64, p_29_65, p_30_0, p_30_1, p_30_2, p_30_3, p_30_4, p_30_5, p_30_6, p_30_7, p_30_8, p_30_9, p_30_10, p_30_11, p_30_12, p_30_13, p_30_14, p_30_15, p_30_16, p_30_17, p_30_18, p_30_19, p_30_20, p_30_21, p_30_22, p_30_23, p_30_24, p_30_25, p_30_26, p_30_27, p_30_28, p_30_29, p_30_30, p_30_31, p_30_32, p_30_33, p_30_34, p_30_35, p_30_36, p_30_37, p_30_38, p_30_39, p_30_40, p_30_41, p_30_42, p_30_43, p_30_44, p_30_45, p_30_46, p_30_47, p_30_48, p_30_49, p_30_50, p_30_51, p_30_52, p_30_53, p_30_54, p_30_55, p_30_56, p_30_57, p_30_58, p_30_59, p_30_60, p_30_61, p_30_62, p_30_63, p_30_64, p_30_65, p_31_0, p_31_1, p_31_2, p_31_3, p_31_4, p_31_5, p_31_6, p_31_7, p_31_8, p_31_9, p_31_10, p_31_11, p_31_12, p_31_13, p_31_14, p_31_15, p_31_16, p_31_17, p_31_18, p_31_19, p_31_20, p_31_21, p_31_22, p_31_23, p_31_24, p_31_25, p_31_26, p_31_27, p_31_28, p_31_29, p_31_30, p_31_31, p_31_32, p_31_33, p_31_34, p_31_35, p_31_36, p_31_37, p_31_38, p_31_39, p_31_40, p_31_41, p_31_42, p_31_43, p_31_44, p_31_45, p_31_46, p_31_47, p_31_48, p_31_49, p_31_50, p_31_51, p_31_52, p_31_53, p_31_54, p_31_55, p_31_56, p_31_57, p_31_58, p_31_59, p_31_60, p_31_61, p_31_62, p_31_63, p_31_64, p_31_65, p_32_0, p_32_1, p_32_2, p_32_3, p_32_4, p_32_5, p_32_6, p_32_7, p_32_8, p_32_9, p_32_10, p_32_11, p_32_12, p_32_13, p_32_14, p_32_15, p_32_16, p_32_17, p_32_18, p_32_19, p_32_20, p_32_21, p_32_22, p_32_23, p_32_24, p_32_25, p_32_26, p_32_27, p_32_28, p_32_29, p_32_30, p_32_31, p_32_32, p_32_33, p_32_34, p_32_35, p_32_36, p_32_37, p_32_38, p_32_39, p_32_40, p_32_41, p_32_42, p_32_43, p_32_44, p_32_45, p_32_46, p_32_47, p_32_48, p_32_49, p_32_50, p_32_51, p_32_52, p_32_53, p_32_54, p_32_55, p_32_56, p_32_57, p_32_58, p_32_59, p_32_60, p_32_61, p_32_62, p_32_63, p_32_64, p_32_65, p_33_0, p_33_1, p_33_2, p_33_3, p_33_4, p_33_5, p_33_6, p_33_7, p_33_8, p_33_9, p_33_10, p_33_11, p_33_12, p_33_13, p_33_14, p_33_15, p_33_16, p_33_17, p_33_18, p_33_19, p_33_20, p_33_21, p_33_22, p_33_23, p_33_24, p_33_25, p_33_26, p_33_27, p_33_28, p_33_29, p_33_30, p_33_31, p_33_32, p_33_33, p_33_34, p_33_35, p_33_36, p_33_37, p_33_38, p_33_39, p_33_40, p_33_41, p_33_42, p_33_43, p_33_44, p_33_45, p_33_46, p_33_47, p_33_48, p_33_49, p_33_50, p_33_51, p_33_52, p_33_53, p_33_54, p_33_55, p_33_56, p_33_57, p_33_58, p_33_59, p_33_60, p_33_61, p_33_62, p_33_63, p_33_64, p_33_65, p_34_0, p_34_1, p_34_2, p_34_3, p_34_4, p_34_5, p_34_6, p_34_7, p_34_8, p_34_9, p_34_10, p_34_11, p_34_12, p_34_13, p_34_14, p_34_15, p_34_16, p_34_17, p_34_18, p_34_19, p_34_20, p_34_21, p_34_22, p_34_23, p_34_24, p_34_25, p_34_26, p_34_27, p_34_28, p_34_29, p_34_30, p_34_31, p_34_32, p_34_33, p_34_34, p_34_35, p_34_36, p_34_37, p_34_38, p_34_39, p_34_40, p_34_41, p_34_42, p_34_43, p_34_44, p_34_45, p_34_46, p_34_47, p_34_48, p_34_49, p_34_50, p_34_51, p_34_52, p_34_53, p_34_54, p_34_55, p_34_56, p_34_57, p_34_58, p_34_59, p_34_60, p_34_61, p_34_62, p_34_63, p_34_64, p_34_65, p_35_0, p_35_1, p_35_2, p_35_3, p_35_4, p_35_5, p_35_6, p_35_7, p_35_8, p_35_9, p_35_10, p_35_11, p_35_12, p_35_13, p_35_14, p_35_15, p_35_16, p_35_17, p_35_18, p_35_19, p_35_20, p_35_21, p_35_22, p_35_23, p_35_24, p_35_25, p_35_26, p_35_27, p_35_28, p_35_29, p_35_30, p_35_31, p_35_32, p_35_33, p_35_34, p_35_35, p_35_36, p_35_37, p_35_38, p_35_39, p_35_40, p_35_41, p_35_42, p_35_43, p_35_44, p_35_45, p_35_46, p_35_47, p_35_48, p_35_49, p_35_50, p_35_51, p_35_52, p_35_53, p_35_54, p_35_55, p_35_56, p_35_57, p_35_58, p_35_59, p_35_60, p_35_61, p_35_62, p_35_63, p_35_64, p_35_65, p_36_0, p_36_1, p_36_2, p_36_3, p_36_4, p_36_5, p_36_6, p_36_7, p_36_8, p_36_9, p_36_10, p_36_11, p_36_12, p_36_13, p_36_14, p_36_15, p_36_16, p_36_17, p_36_18, p_36_19, p_36_20, p_36_21, p_36_22, p_36_23, p_36_24, p_36_25, p_36_26, p_36_27, p_36_28, p_36_29, p_36_30, p_36_31, p_36_32, p_36_33, p_36_34, p_36_35, p_36_36, p_36_37, p_36_38, p_36_39, p_36_40, p_36_41, p_36_42, p_36_43, p_36_44, p_36_45, p_36_46, p_36_47, p_36_48, p_36_49, p_36_50, p_36_51, p_36_52, p_36_53, p_36_54, p_36_55, p_36_56, p_36_57, p_36_58, p_36_59, p_36_60, p_36_61, p_36_62, p_36_63, p_36_64, p_36_65, p_37_0, p_37_1, p_37_2, p_37_3, p_37_4, p_37_5, p_37_6, p_37_7, p_37_8, p_37_9, p_37_10, p_37_11, p_37_12, p_37_13, p_37_14, p_37_15, p_37_16, p_37_17, p_37_18, p_37_19, p_37_20, p_37_21, p_37_22, p_37_23, p_37_24, p_37_25, p_37_26, p_37_27, p_37_28, p_37_29, p_37_30, p_37_31, p_37_32, p_37_33, p_37_34, p_37_35, p_37_36, p_37_37, p_37_38, p_37_39, p_37_40, p_37_41, p_37_42, p_37_43, p_37_44, p_37_45, p_37_46, p_37_47, p_37_48, p_37_49, p_37_50, p_37_51, p_37_52, p_37_53, p_37_54, p_37_55, p_37_56, p_37_57, p_37_58, p_37_59, p_37_60, p_37_61, p_37_62, p_37_63, p_37_64, p_37_65, p_38_0, p_38_1, p_38_2, p_38_3, p_38_4, p_38_5, p_38_6, p_38_7, p_38_8, p_38_9, p_38_10, p_38_11, p_38_12, p_38_13, p_38_14, p_38_15, p_38_16, p_38_17, p_38_18, p_38_19, p_38_20, p_38_21, p_38_22, p_38_23, p_38_24, p_38_25, p_38_26, p_38_27, p_38_28, p_38_29, p_38_30, p_38_31, p_38_32, p_38_33, p_38_34, p_38_35, p_38_36, p_38_37, p_38_38, p_38_39, p_38_40, p_38_41, p_38_42, p_38_43, p_38_44, p_38_45, p_38_46, p_38_47, p_38_48, p_38_49, p_38_50, p_38_51, p_38_52, p_38_53, p_38_54, p_38_55, p_38_56, p_38_57, p_38_58, p_38_59, p_38_60, p_38_61, p_38_62, p_38_63, p_38_64, p_38_65, p_39_0, p_39_1, p_39_2, p_39_3, p_39_4, p_39_5, p_39_6, p_39_7, p_39_8, p_39_9, p_39_10, p_39_11, p_39_12, p_39_13, p_39_14, p_39_15, p_39_16, p_39_17, p_39_18, p_39_19, p_39_20, p_39_21, p_39_22, p_39_23, p_39_24, p_39_25, p_39_26, p_39_27, p_39_28, p_39_29, p_39_30, p_39_31, p_39_32, p_39_33, p_39_34, p_39_35, p_39_36, p_39_37, p_39_38, p_39_39, p_39_40, p_39_41, p_39_42, p_39_43, p_39_44, p_39_45, p_39_46, p_39_47, p_39_48, p_39_49, p_39_50, p_39_51, p_39_52, p_39_53, p_39_54, p_39_55, p_39_56, p_39_57, p_39_58, p_39_59, p_39_60, p_39_61, p_39_62, p_39_63, p_39_64, p_39_65, p_40_0, p_40_1, p_40_2, p_40_3, p_40_4, p_40_5, p_40_6, p_40_7, p_40_8, p_40_9, p_40_10, p_40_11, p_40_12, p_40_13, p_40_14, p_40_15, p_40_16, p_40_17, p_40_18, p_40_19, p_40_20, p_40_21, p_40_22, p_40_23, p_40_24, p_40_25, p_40_26, p_40_27, p_40_28, p_40_29, p_40_30, p_40_31, p_40_32, p_40_33, p_40_34, p_40_35, p_40_36, p_40_37, p_40_38, p_40_39, p_40_40, p_40_41, p_40_42, p_40_43, p_40_44, p_40_45, p_40_46, p_40_47, p_40_48, p_40_49, p_40_50, p_40_51, p_40_52, p_40_53, p_40_54, p_40_55, p_40_56, p_40_57, p_40_58, p_40_59, p_40_60, p_40_61, p_40_62, p_40_63, p_40_64, p_40_65, p_41_0, p_41_1, p_41_2, p_41_3, p_41_4, p_41_5, p_41_6, p_41_7, p_41_8, p_41_9, p_41_10, p_41_11, p_41_12, p_41_13, p_41_14, p_41_15, p_41_16, p_41_17, p_41_18, p_41_19, p_41_20, p_41_21, p_41_22, p_41_23, p_41_24, p_41_25, p_41_26, p_41_27, p_41_28, p_41_29, p_41_30, p_41_31, p_41_32, p_41_33, p_41_34, p_41_35, p_41_36, p_41_37, p_41_38, p_41_39, p_41_40, p_41_41, p_41_42, p_41_43, p_41_44, p_41_45, p_41_46, p_41_47, p_41_48, p_41_49, p_41_50, p_41_51, p_41_52, p_41_53, p_41_54, p_41_55, p_41_56, p_41_57, p_41_58, p_41_59, p_41_60, p_41_61, p_41_62, p_41_63, p_41_64, p_41_65, p_42_0, p_42_1, p_42_2, p_42_3, p_42_4, p_42_5, p_42_6, p_42_7, p_42_8, p_42_9, p_42_10, p_42_11, p_42_12, p_42_13, p_42_14, p_42_15, p_42_16, p_42_17, p_42_18, p_42_19, p_42_20, p_42_21, p_42_22, p_42_23, p_42_24, p_42_25, p_42_26, p_42_27, p_42_28, p_42_29, p_42_30, p_42_31, p_42_32, p_42_33, p_42_34, p_42_35, p_42_36, p_42_37, p_42_38, p_42_39, p_42_40, p_42_41, p_42_42, p_42_43, p_42_44, p_42_45, p_42_46, p_42_47, p_42_48, p_42_49, p_42_50, p_42_51, p_42_52, p_42_53, p_42_54, p_42_55, p_42_56, p_42_57, p_42_58, p_42_59, p_42_60, p_42_61, p_42_62, p_42_63, p_42_64, p_42_65, p_43_0, p_43_1, p_43_2, p_43_3, p_43_4, p_43_5, p_43_6, p_43_7, p_43_8, p_43_9, p_43_10, p_43_11, p_43_12, p_43_13, p_43_14, p_43_15, p_43_16, p_43_17, p_43_18, p_43_19, p_43_20, p_43_21, p_43_22, p_43_23, p_43_24, p_43_25, p_43_26, p_43_27, p_43_28, p_43_29, p_43_30, p_43_31, p_43_32, p_43_33, p_43_34, p_43_35, p_43_36, p_43_37, p_43_38, p_43_39, p_43_40, p_43_41, p_43_42, p_43_43, p_43_44, p_43_45, p_43_46, p_43_47, p_43_48, p_43_49, p_43_50, p_43_51, p_43_52, p_43_53, p_43_54, p_43_55, p_43_56, p_43_57, p_43_58, p_43_59, p_43_60, p_43_61, p_43_62, p_43_63, p_43_64, p_43_65, p_44_0, p_44_1, p_44_2, p_44_3, p_44_4, p_44_5, p_44_6, p_44_7, p_44_8, p_44_9, p_44_10, p_44_11, p_44_12, p_44_13, p_44_14, p_44_15, p_44_16, p_44_17, p_44_18, p_44_19, p_44_20, p_44_21, p_44_22, p_44_23, p_44_24, p_44_25, p_44_26, p_44_27, p_44_28, p_44_29, p_44_30, p_44_31, p_44_32, p_44_33, p_44_34, p_44_35, p_44_36, p_44_37, p_44_38, p_44_39, p_44_40, p_44_41, p_44_42, p_44_43, p_44_44, p_44_45, p_44_46, p_44_47, p_44_48, p_44_49, p_44_50, p_44_51, p_44_52, p_44_53, p_44_54, p_44_55, p_44_56, p_44_57, p_44_58, p_44_59, p_44_60, p_44_61, p_44_62, p_44_63, p_44_64, p_44_65, out_1_1, out_1_2, out_1_3, out_1_4, out_1_5, out_1_6, out_1_7, out_1_8, out_1_9, out_1_10, out_1_11, out_1_12, out_1_13, out_1_14, out_1_15, out_1_16, out_1_17, out_1_18, out_1_19, out_1_20, out_1_21, out_1_22, out_1_23, out_1_24, out_1_25, out_1_26, out_1_27, out_1_28, out_1_29, out_1_30, out_1_31, out_1_32, out_1_33, out_1_34, out_1_35, out_1_36, out_1_37, out_1_38, out_1_39, out_1_40, out_1_41, out_1_42, out_1_43, out_1_44, out_1_45, out_1_46, out_1_47, out_1_48, out_1_49, out_1_50, out_1_51, out_1_52, out_1_53, out_1_54, out_1_55, out_1_56, out_1_57, out_1_58, out_1_59, out_1_60, out_1_61, out_1_62, out_1_63, out_1_64, out_2_1, out_2_2, out_2_3, out_2_4, out_2_5, out_2_6, out_2_7, out_2_8, out_2_9, out_2_10, out_2_11, out_2_12, out_2_13, out_2_14, out_2_15, out_2_16, out_2_17, out_2_18, out_2_19, out_2_20, out_2_21, out_2_22, out_2_23, out_2_24, out_2_25, out_2_26, out_2_27, out_2_28, out_2_29, out_2_30, out_2_31, out_2_32, out_2_33, out_2_34, out_2_35, out_2_36, out_2_37, out_2_38, out_2_39, out_2_40, out_2_41, out_2_42, out_2_43, out_2_44, out_2_45, out_2_46, out_2_47, out_2_48, out_2_49, out_2_50, out_2_51, out_2_52, out_2_53, out_2_54, out_2_55, out_2_56, out_2_57, out_2_58, out_2_59, out_2_60, out_2_61, out_2_62, out_2_63, out_2_64, out_3_1, out_3_2, out_3_3, out_3_4, out_3_5, out_3_6, out_3_7, out_3_8, out_3_9, out_3_10, out_3_11, out_3_12, out_3_13, out_3_14, out_3_15, out_3_16, out_3_17, out_3_18, out_3_19, out_3_20, out_3_21, out_3_22, out_3_23, out_3_24, out_3_25, out_3_26, out_3_27, out_3_28, out_3_29, out_3_30, out_3_31, out_3_32, out_3_33, out_3_34, out_3_35, out_3_36, out_3_37, out_3_38, out_3_39, out_3_40, out_3_41, out_3_42, out_3_43, out_3_44, out_3_45, out_3_46, out_3_47, out_3_48, out_3_49, out_3_50, out_3_51, out_3_52, out_3_53, out_3_54, out_3_55, out_3_56, out_3_57, out_3_58, out_3_59, out_3_60, out_3_61, out_3_62, out_3_63, out_3_64, out_4_1, out_4_2, out_4_3, out_4_4, out_4_5, out_4_6, out_4_7, out_4_8, out_4_9, out_4_10, out_4_11, out_4_12, out_4_13, out_4_14, out_4_15, out_4_16, out_4_17, out_4_18, out_4_19, out_4_20, out_4_21, out_4_22, out_4_23, out_4_24, out_4_25, out_4_26, out_4_27, out_4_28, out_4_29, out_4_30, out_4_31, out_4_32, out_4_33, out_4_34, out_4_35, out_4_36, out_4_37, out_4_38, out_4_39, out_4_40, out_4_41, out_4_42, out_4_43, out_4_44, out_4_45, out_4_46, out_4_47, out_4_48, out_4_49, out_4_50, out_4_51, out_4_52, out_4_53, out_4_54, out_4_55, out_4_56, out_4_57, out_4_58, out_4_59, out_4_60, out_4_61, out_4_62, out_4_63, out_4_64, out_5_1, out_5_2, out_5_3, out_5_4, out_5_5, out_5_6, out_5_7, out_5_8, out_5_9, out_5_10, out_5_11, out_5_12, out_5_13, out_5_14, out_5_15, out_5_16, out_5_17, out_5_18, out_5_19, out_5_20, out_5_21, out_5_22, out_5_23, out_5_24, out_5_25, out_5_26, out_5_27, out_5_28, out_5_29, out_5_30, out_5_31, out_5_32, out_5_33, out_5_34, out_5_35, out_5_36, out_5_37, out_5_38, out_5_39, out_5_40, out_5_41, out_5_42, out_5_43, out_5_44, out_5_45, out_5_46, out_5_47, out_5_48, out_5_49, out_5_50, out_5_51, out_5_52, out_5_53, out_5_54, out_5_55, out_5_56, out_5_57, out_5_58, out_5_59, out_5_60, out_5_61, out_5_62, out_5_63, out_5_64, out_6_1, out_6_2, out_6_3, out_6_4, out_6_5, out_6_6, out_6_7, out_6_8, out_6_9, out_6_10, out_6_11, out_6_12, out_6_13, out_6_14, out_6_15, out_6_16, out_6_17, out_6_18, out_6_19, out_6_20, out_6_21, out_6_22, out_6_23, out_6_24, out_6_25, out_6_26, out_6_27, out_6_28, out_6_29, out_6_30, out_6_31, out_6_32, out_6_33, out_6_34, out_6_35, out_6_36, out_6_37, out_6_38, out_6_39, out_6_40, out_6_41, out_6_42, out_6_43, out_6_44, out_6_45, out_6_46, out_6_47, out_6_48, out_6_49, out_6_50, out_6_51, out_6_52, out_6_53, out_6_54, out_6_55, out_6_56, out_6_57, out_6_58, out_6_59, out_6_60, out_6_61, out_6_62, out_6_63, out_6_64, out_7_1, out_7_2, out_7_3, out_7_4, out_7_5, out_7_6, out_7_7, out_7_8, out_7_9, out_7_10, out_7_11, out_7_12, out_7_13, out_7_14, out_7_15, out_7_16, out_7_17, out_7_18, out_7_19, out_7_20, out_7_21, out_7_22, out_7_23, out_7_24, out_7_25, out_7_26, out_7_27, out_7_28, out_7_29, out_7_30, out_7_31, out_7_32, out_7_33, out_7_34, out_7_35, out_7_36, out_7_37, out_7_38, out_7_39, out_7_40, out_7_41, out_7_42, out_7_43, out_7_44, out_7_45, out_7_46, out_7_47, out_7_48, out_7_49, out_7_50, out_7_51, out_7_52, out_7_53, out_7_54, out_7_55, out_7_56, out_7_57, out_7_58, out_7_59, out_7_60, out_7_61, out_7_62, out_7_63, out_7_64, out_8_1, out_8_2, out_8_3, out_8_4, out_8_5, out_8_6, out_8_7, out_8_8, out_8_9, out_8_10, out_8_11, out_8_12, out_8_13, out_8_14, out_8_15, out_8_16, out_8_17, out_8_18, out_8_19, out_8_20, out_8_21, out_8_22, out_8_23, out_8_24, out_8_25, out_8_26, out_8_27, out_8_28, out_8_29, out_8_30, out_8_31, out_8_32, out_8_33, out_8_34, out_8_35, out_8_36, out_8_37, out_8_38, out_8_39, out_8_40, out_8_41, out_8_42, out_8_43, out_8_44, out_8_45, out_8_46, out_8_47, out_8_48, out_8_49, out_8_50, out_8_51, out_8_52, out_8_53, out_8_54, out_8_55, out_8_56, out_8_57, out_8_58, out_8_59, out_8_60, out_8_61, out_8_62, out_8_63, out_8_64, out_9_1, out_9_2, out_9_3, out_9_4, out_9_5, out_9_6, out_9_7, out_9_8, out_9_9, out_9_10, out_9_11, out_9_12, out_9_13, out_9_14, out_9_15, out_9_16, out_9_17, out_9_18, out_9_19, out_9_20, out_9_21, out_9_22, out_9_23, out_9_24, out_9_25, out_9_26, out_9_27, out_9_28, out_9_29, out_9_30, out_9_31, out_9_32, out_9_33, out_9_34, out_9_35, out_9_36, out_9_37, out_9_38, out_9_39, out_9_40, out_9_41, out_9_42, out_9_43, out_9_44, out_9_45, out_9_46, out_9_47, out_9_48, out_9_49, out_9_50, out_9_51, out_9_52, out_9_53, out_9_54, out_9_55, out_9_56, out_9_57, out_9_58, out_9_59, out_9_60, out_9_61, out_9_62, out_9_63, out_9_64, out_10_1, out_10_2, out_10_3, out_10_4, out_10_5, out_10_6, out_10_7, out_10_8, out_10_9, out_10_10, out_10_11, out_10_12, out_10_13, out_10_14, out_10_15, out_10_16, out_10_17, out_10_18, out_10_19, out_10_20, out_10_21, out_10_22, out_10_23, out_10_24, out_10_25, out_10_26, out_10_27, out_10_28, out_10_29, out_10_30, out_10_31, out_10_32, out_10_33, out_10_34, out_10_35, out_10_36, out_10_37, out_10_38, out_10_39, out_10_40, out_10_41, out_10_42, out_10_43, out_10_44, out_10_45, out_10_46, out_10_47, out_10_48, out_10_49, out_10_50, out_10_51, out_10_52, out_10_53, out_10_54, out_10_55, out_10_56, out_10_57, out_10_58, out_10_59, out_10_60, out_10_61, out_10_62, out_10_63, out_10_64, out_11_1, out_11_2, out_11_3, out_11_4, out_11_5, out_11_6, out_11_7, out_11_8, out_11_9, out_11_10, out_11_11, out_11_12, out_11_13, out_11_14, out_11_15, out_11_16, out_11_17, out_11_18, out_11_19, out_11_20, out_11_21, out_11_22, out_11_23, out_11_24, out_11_25, out_11_26, out_11_27, out_11_28, out_11_29, out_11_30, out_11_31, out_11_32, out_11_33, out_11_34, out_11_35, out_11_36, out_11_37, out_11_38, out_11_39, out_11_40, out_11_41, out_11_42, out_11_43, out_11_44, out_11_45, out_11_46, out_11_47, out_11_48, out_11_49, out_11_50, out_11_51, out_11_52, out_11_53, out_11_54, out_11_55, out_11_56, out_11_57, out_11_58, out_11_59, out_11_60, out_11_61, out_11_62, out_11_63, out_11_64, out_12_1, out_12_2, out_12_3, out_12_4, out_12_5, out_12_6, out_12_7, out_12_8, out_12_9, out_12_10, out_12_11, out_12_12, out_12_13, out_12_14, out_12_15, out_12_16, out_12_17, out_12_18, out_12_19, out_12_20, out_12_21, out_12_22, out_12_23, out_12_24, out_12_25, out_12_26, out_12_27, out_12_28, out_12_29, out_12_30, out_12_31, out_12_32, out_12_33, out_12_34, out_12_35, out_12_36, out_12_37, out_12_38, out_12_39, out_12_40, out_12_41, out_12_42, out_12_43, out_12_44, out_12_45, out_12_46, out_12_47, out_12_48, out_12_49, out_12_50, out_12_51, out_12_52, out_12_53, out_12_54, out_12_55, out_12_56, out_12_57, out_12_58, out_12_59, out_12_60, out_12_61, out_12_62, out_12_63, out_12_64, out_13_1, out_13_2, out_13_3, out_13_4, out_13_5, out_13_6, out_13_7, out_13_8, out_13_9, out_13_10, out_13_11, out_13_12, out_13_13, out_13_14, out_13_15, out_13_16, out_13_17, out_13_18, out_13_19, out_13_20, out_13_21, out_13_22, out_13_23, out_13_24, out_13_25, out_13_26, out_13_27, out_13_28, out_13_29, out_13_30, out_13_31, out_13_32, out_13_33, out_13_34, out_13_35, out_13_36, out_13_37, out_13_38, out_13_39, out_13_40, out_13_41, out_13_42, out_13_43, out_13_44, out_13_45, out_13_46, out_13_47, out_13_48, out_13_49, out_13_50, out_13_51, out_13_52, out_13_53, out_13_54, out_13_55, out_13_56, out_13_57, out_13_58, out_13_59, out_13_60, out_13_61, out_13_62, out_13_63, out_13_64, out_14_1, out_14_2, out_14_3, out_14_4, out_14_5, out_14_6, out_14_7, out_14_8, out_14_9, out_14_10, out_14_11, out_14_12, out_14_13, out_14_14, out_14_15, out_14_16, out_14_17, out_14_18, out_14_19, out_14_20, out_14_21, out_14_22, out_14_23, out_14_24, out_14_25, out_14_26, out_14_27, out_14_28, out_14_29, out_14_30, out_14_31, out_14_32, out_14_33, out_14_34, out_14_35, out_14_36, out_14_37, out_14_38, out_14_39, out_14_40, out_14_41, out_14_42, out_14_43, out_14_44, out_14_45, out_14_46, out_14_47, out_14_48, out_14_49, out_14_50, out_14_51, out_14_52, out_14_53, out_14_54, out_14_55, out_14_56, out_14_57, out_14_58, out_14_59, out_14_60, out_14_61, out_14_62, out_14_63, out_14_64, out_15_1, out_15_2, out_15_3, out_15_4, out_15_5, out_15_6, out_15_7, out_15_8, out_15_9, out_15_10, out_15_11, out_15_12, out_15_13, out_15_14, out_15_15, out_15_16, out_15_17, out_15_18, out_15_19, out_15_20, out_15_21, out_15_22, out_15_23, out_15_24, out_15_25, out_15_26, out_15_27, out_15_28, out_15_29, out_15_30, out_15_31, out_15_32, out_15_33, out_15_34, out_15_35, out_15_36, out_15_37, out_15_38, out_15_39, out_15_40, out_15_41, out_15_42, out_15_43, out_15_44, out_15_45, out_15_46, out_15_47, out_15_48, out_15_49, out_15_50, out_15_51, out_15_52, out_15_53, out_15_54, out_15_55, out_15_56, out_15_57, out_15_58, out_15_59, out_15_60, out_15_61, out_15_62, out_15_63, out_15_64, out_16_1, out_16_2, out_16_3, out_16_4, out_16_5, out_16_6, out_16_7, out_16_8, out_16_9, out_16_10, out_16_11, out_16_12, out_16_13, out_16_14, out_16_15, out_16_16, out_16_17, out_16_18, out_16_19, out_16_20, out_16_21, out_16_22, out_16_23, out_16_24, out_16_25, out_16_26, out_16_27, out_16_28, out_16_29, out_16_30, out_16_31, out_16_32, out_16_33, out_16_34, out_16_35, out_16_36, out_16_37, out_16_38, out_16_39, out_16_40, out_16_41, out_16_42, out_16_43, out_16_44, out_16_45, out_16_46, out_16_47, out_16_48, out_16_49, out_16_50, out_16_51, out_16_52, out_16_53, out_16_54, out_16_55, out_16_56, out_16_57, out_16_58, out_16_59, out_16_60, out_16_61, out_16_62, out_16_63, out_16_64, out_17_1, out_17_2, out_17_3, out_17_4, out_17_5, out_17_6, out_17_7, out_17_8, out_17_9, out_17_10, out_17_11, out_17_12, out_17_13, out_17_14, out_17_15, out_17_16, out_17_17, out_17_18, out_17_19, out_17_20, out_17_21, out_17_22, out_17_23, out_17_24, out_17_25, out_17_26, out_17_27, out_17_28, out_17_29, out_17_30, out_17_31, out_17_32, out_17_33, out_17_34, out_17_35, out_17_36, out_17_37, out_17_38, out_17_39, out_17_40, out_17_41, out_17_42, out_17_43, out_17_44, out_17_45, out_17_46, out_17_47, out_17_48, out_17_49, out_17_50, out_17_51, out_17_52, out_17_53, out_17_54, out_17_55, out_17_56, out_17_57, out_17_58, out_17_59, out_17_60, out_17_61, out_17_62, out_17_63, out_17_64, out_18_1, out_18_2, out_18_3, out_18_4, out_18_5, out_18_6, out_18_7, out_18_8, out_18_9, out_18_10, out_18_11, out_18_12, out_18_13, out_18_14, out_18_15, out_18_16, out_18_17, out_18_18, out_18_19, out_18_20, out_18_21, out_18_22, out_18_23, out_18_24, out_18_25, out_18_26, out_18_27, out_18_28, out_18_29, out_18_30, out_18_31, out_18_32, out_18_33, out_18_34, out_18_35, out_18_36, out_18_37, out_18_38, out_18_39, out_18_40, out_18_41, out_18_42, out_18_43, out_18_44, out_18_45, out_18_46, out_18_47, out_18_48, out_18_49, out_18_50, out_18_51, out_18_52, out_18_53, out_18_54, out_18_55, out_18_56, out_18_57, out_18_58, out_18_59, out_18_60, out_18_61, out_18_62, out_18_63, out_18_64, out_19_1, out_19_2, out_19_3, out_19_4, out_19_5, out_19_6, out_19_7, out_19_8, out_19_9, out_19_10, out_19_11, out_19_12, out_19_13, out_19_14, out_19_15, out_19_16, out_19_17, out_19_18, out_19_19, out_19_20, out_19_21, out_19_22, out_19_23, out_19_24, out_19_25, out_19_26, out_19_27, out_19_28, out_19_29, out_19_30, out_19_31, out_19_32, out_19_33, out_19_34, out_19_35, out_19_36, out_19_37, out_19_38, out_19_39, out_19_40, out_19_41, out_19_42, out_19_43, out_19_44, out_19_45, out_19_46, out_19_47, out_19_48, out_19_49, out_19_50, out_19_51, out_19_52, out_19_53, out_19_54, out_19_55, out_19_56, out_19_57, out_19_58, out_19_59, out_19_60, out_19_61, out_19_62, out_19_63, out_19_64, out_20_1, out_20_2, out_20_3, out_20_4, out_20_5, out_20_6, out_20_7, out_20_8, out_20_9, out_20_10, out_20_11, out_20_12, out_20_13, out_20_14, out_20_15, out_20_16, out_20_17, out_20_18, out_20_19, out_20_20, out_20_21, out_20_22, out_20_23, out_20_24, out_20_25, out_20_26, out_20_27, out_20_28, out_20_29, out_20_30, out_20_31, out_20_32, out_20_33, out_20_34, out_20_35, out_20_36, out_20_37, out_20_38, out_20_39, out_20_40, out_20_41, out_20_42, out_20_43, out_20_44, out_20_45, out_20_46, out_20_47, out_20_48, out_20_49, out_20_50, out_20_51, out_20_52, out_20_53, out_20_54, out_20_55, out_20_56, out_20_57, out_20_58, out_20_59, out_20_60, out_20_61, out_20_62, out_20_63, out_20_64, out_21_1, out_21_2, out_21_3, out_21_4, out_21_5, out_21_6, out_21_7, out_21_8, out_21_9, out_21_10, out_21_11, out_21_12, out_21_13, out_21_14, out_21_15, out_21_16, out_21_17, out_21_18, out_21_19, out_21_20, out_21_21, out_21_22, out_21_23, out_21_24, out_21_25, out_21_26, out_21_27, out_21_28, out_21_29, out_21_30, out_21_31, out_21_32, out_21_33, out_21_34, out_21_35, out_21_36, out_21_37, out_21_38, out_21_39, out_21_40, out_21_41, out_21_42, out_21_43, out_21_44, out_21_45, out_21_46, out_21_47, out_21_48, out_21_49, out_21_50, out_21_51, out_21_52, out_21_53, out_21_54, out_21_55, out_21_56, out_21_57, out_21_58, out_21_59, out_21_60, out_21_61, out_21_62, out_21_63, out_21_64, out_22_1, out_22_2, out_22_3, out_22_4, out_22_5, out_22_6, out_22_7, out_22_8, out_22_9, out_22_10, out_22_11, out_22_12, out_22_13, out_22_14, out_22_15, out_22_16, out_22_17, out_22_18, out_22_19, out_22_20, out_22_21, out_22_22, out_22_23, out_22_24, out_22_25, out_22_26, out_22_27, out_22_28, out_22_29, out_22_30, out_22_31, out_22_32, out_22_33, out_22_34, out_22_35, out_22_36, out_22_37, out_22_38, out_22_39, out_22_40, out_22_41, out_22_42, out_22_43, out_22_44, out_22_45, out_22_46, out_22_47, out_22_48, out_22_49, out_22_50, out_22_51, out_22_52, out_22_53, out_22_54, out_22_55, out_22_56, out_22_57, out_22_58, out_22_59, out_22_60, out_22_61, out_22_62, out_22_63, out_22_64, out_23_1, out_23_2, out_23_3, out_23_4, out_23_5, out_23_6, out_23_7, out_23_8, out_23_9, out_23_10, out_23_11, out_23_12, out_23_13, out_23_14, out_23_15, out_23_16, out_23_17, out_23_18, out_23_19, out_23_20, out_23_21, out_23_22, out_23_23, out_23_24, out_23_25, out_23_26, out_23_27, out_23_28, out_23_29, out_23_30, out_23_31, out_23_32, out_23_33, out_23_34, out_23_35, out_23_36, out_23_37, out_23_38, out_23_39, out_23_40, out_23_41, out_23_42, out_23_43, out_23_44, out_23_45, out_23_46, out_23_47, out_23_48, out_23_49, out_23_50, out_23_51, out_23_52, out_23_53, out_23_54, out_23_55, out_23_56, out_23_57, out_23_58, out_23_59, out_23_60, out_23_61, out_23_62, out_23_63, out_23_64, out_24_1, out_24_2, out_24_3, out_24_4, out_24_5, out_24_6, out_24_7, out_24_8, out_24_9, out_24_10, out_24_11, out_24_12, out_24_13, out_24_14, out_24_15, out_24_16, out_24_17, out_24_18, out_24_19, out_24_20, out_24_21, out_24_22, out_24_23, out_24_24, out_24_25, out_24_26, out_24_27, out_24_28, out_24_29, out_24_30, out_24_31, out_24_32, out_24_33, out_24_34, out_24_35, out_24_36, out_24_37, out_24_38, out_24_39, out_24_40, out_24_41, out_24_42, out_24_43, out_24_44, out_24_45, out_24_46, out_24_47, out_24_48, out_24_49, out_24_50, out_24_51, out_24_52, out_24_53, out_24_54, out_24_55, out_24_56, out_24_57, out_24_58, out_24_59, out_24_60, out_24_61, out_24_62, out_24_63, out_24_64, out_25_1, out_25_2, out_25_3, out_25_4, out_25_5, out_25_6, out_25_7, out_25_8, out_25_9, out_25_10, out_25_11, out_25_12, out_25_13, out_25_14, out_25_15, out_25_16, out_25_17, out_25_18, out_25_19, out_25_20, out_25_21, out_25_22, out_25_23, out_25_24, out_25_25, out_25_26, out_25_27, out_25_28, out_25_29, out_25_30, out_25_31, out_25_32, out_25_33, out_25_34, out_25_35, out_25_36, out_25_37, out_25_38, out_25_39, out_25_40, out_25_41, out_25_42, out_25_43, out_25_44, out_25_45, out_25_46, out_25_47, out_25_48, out_25_49, out_25_50, out_25_51, out_25_52, out_25_53, out_25_54, out_25_55, out_25_56, out_25_57, out_25_58, out_25_59, out_25_60, out_25_61, out_25_62, out_25_63, out_25_64, out_26_1, out_26_2, out_26_3, out_26_4, out_26_5, out_26_6, out_26_7, out_26_8, out_26_9, out_26_10, out_26_11, out_26_12, out_26_13, out_26_14, out_26_15, out_26_16, out_26_17, out_26_18, out_26_19, out_26_20, out_26_21, out_26_22, out_26_23, out_26_24, out_26_25, out_26_26, out_26_27, out_26_28, out_26_29, out_26_30, out_26_31, out_26_32, out_26_33, out_26_34, out_26_35, out_26_36, out_26_37, out_26_38, out_26_39, out_26_40, out_26_41, out_26_42, out_26_43, out_26_44, out_26_45, out_26_46, out_26_47, out_26_48, out_26_49, out_26_50, out_26_51, out_26_52, out_26_53, out_26_54, out_26_55, out_26_56, out_26_57, out_26_58, out_26_59, out_26_60, out_26_61, out_26_62, out_26_63, out_26_64, out_27_1, out_27_2, out_27_3, out_27_4, out_27_5, out_27_6, out_27_7, out_27_8, out_27_9, out_27_10, out_27_11, out_27_12, out_27_13, out_27_14, out_27_15, out_27_16, out_27_17, out_27_18, out_27_19, out_27_20, out_27_21, out_27_22, out_27_23, out_27_24, out_27_25, out_27_26, out_27_27, out_27_28, out_27_29, out_27_30, out_27_31, out_27_32, out_27_33, out_27_34, out_27_35, out_27_36, out_27_37, out_27_38, out_27_39, out_27_40, out_27_41, out_27_42, out_27_43, out_27_44, out_27_45, out_27_46, out_27_47, out_27_48, out_27_49, out_27_50, out_27_51, out_27_52, out_27_53, out_27_54, out_27_55, out_27_56, out_27_57, out_27_58, out_27_59, out_27_60, out_27_61, out_27_62, out_27_63, out_27_64, out_28_1, out_28_2, out_28_3, out_28_4, out_28_5, out_28_6, out_28_7, out_28_8, out_28_9, out_28_10, out_28_11, out_28_12, out_28_13, out_28_14, out_28_15, out_28_16, out_28_17, out_28_18, out_28_19, out_28_20, out_28_21, out_28_22, out_28_23, out_28_24, out_28_25, out_28_26, out_28_27, out_28_28, out_28_29, out_28_30, out_28_31, out_28_32, out_28_33, out_28_34, out_28_35, out_28_36, out_28_37, out_28_38, out_28_39, out_28_40, out_28_41, out_28_42, out_28_43, out_28_44, out_28_45, out_28_46, out_28_47, out_28_48, out_28_49, out_28_50, out_28_51, out_28_52, out_28_53, out_28_54, out_28_55, out_28_56, out_28_57, out_28_58, out_28_59, out_28_60, out_28_61, out_28_62, out_28_63, out_28_64, out_29_1, out_29_2, out_29_3, out_29_4, out_29_5, out_29_6, out_29_7, out_29_8, out_29_9, out_29_10, out_29_11, out_29_12, out_29_13, out_29_14, out_29_15, out_29_16, out_29_17, out_29_18, out_29_19, out_29_20, out_29_21, out_29_22, out_29_23, out_29_24, out_29_25, out_29_26, out_29_27, out_29_28, out_29_29, out_29_30, out_29_31, out_29_32, out_29_33, out_29_34, out_29_35, out_29_36, out_29_37, out_29_38, out_29_39, out_29_40, out_29_41, out_29_42, out_29_43, out_29_44, out_29_45, out_29_46, out_29_47, out_29_48, out_29_49, out_29_50, out_29_51, out_29_52, out_29_53, out_29_54, out_29_55, out_29_56, out_29_57, out_29_58, out_29_59, out_29_60, out_29_61, out_29_62, out_29_63, out_29_64, out_30_1, out_30_2, out_30_3, out_30_4, out_30_5, out_30_6, out_30_7, out_30_8, out_30_9, out_30_10, out_30_11, out_30_12, out_30_13, out_30_14, out_30_15, out_30_16, out_30_17, out_30_18, out_30_19, out_30_20, out_30_21, out_30_22, out_30_23, out_30_24, out_30_25, out_30_26, out_30_27, out_30_28, out_30_29, out_30_30, out_30_31, out_30_32, out_30_33, out_30_34, out_30_35, out_30_36, out_30_37, out_30_38, out_30_39, out_30_40, out_30_41, out_30_42, out_30_43, out_30_44, out_30_45, out_30_46, out_30_47, out_30_48, out_30_49, out_30_50, out_30_51, out_30_52, out_30_53, out_30_54, out_30_55, out_30_56, out_30_57, out_30_58, out_30_59, out_30_60, out_30_61, out_30_62, out_30_63, out_30_64, out_31_1, out_31_2, out_31_3, out_31_4, out_31_5, out_31_6, out_31_7, out_31_8, out_31_9, out_31_10, out_31_11, out_31_12, out_31_13, out_31_14, out_31_15, out_31_16, out_31_17, out_31_18, out_31_19, out_31_20, out_31_21, out_31_22, out_31_23, out_31_24, out_31_25, out_31_26, out_31_27, out_31_28, out_31_29, out_31_30, out_31_31, out_31_32, out_31_33, out_31_34, out_31_35, out_31_36, out_31_37, out_31_38, out_31_39, out_31_40, out_31_41, out_31_42, out_31_43, out_31_44, out_31_45, out_31_46, out_31_47, out_31_48, out_31_49, out_31_50, out_31_51, out_31_52, out_31_53, out_31_54, out_31_55, out_31_56, out_31_57, out_31_58, out_31_59, out_31_60, out_31_61, out_31_62, out_31_63, out_31_64, out_32_1, out_32_2, out_32_3, out_32_4, out_32_5, out_32_6, out_32_7, out_32_8, out_32_9, out_32_10, out_32_11, out_32_12, out_32_13, out_32_14, out_32_15, out_32_16, out_32_17, out_32_18, out_32_19, out_32_20, out_32_21, out_32_22, out_32_23, out_32_24, out_32_25, out_32_26, out_32_27, out_32_28, out_32_29, out_32_30, out_32_31, out_32_32, out_32_33, out_32_34, out_32_35, out_32_36, out_32_37, out_32_38, out_32_39, out_32_40, out_32_41, out_32_42, out_32_43, out_32_44, out_32_45, out_32_46, out_32_47, out_32_48, out_32_49, out_32_50, out_32_51, out_32_52, out_32_53, out_32_54, out_32_55, out_32_56, out_32_57, out_32_58, out_32_59, out_32_60, out_32_61, out_32_62, out_32_63, out_32_64, out_33_1, out_33_2, out_33_3, out_33_4, out_33_5, out_33_6, out_33_7, out_33_8, out_33_9, out_33_10, out_33_11, out_33_12, out_33_13, out_33_14, out_33_15, out_33_16, out_33_17, out_33_18, out_33_19, out_33_20, out_33_21, out_33_22, out_33_23, out_33_24, out_33_25, out_33_26, out_33_27, out_33_28, out_33_29, out_33_30, out_33_31, out_33_32, out_33_33, out_33_34, out_33_35, out_33_36, out_33_37, out_33_38, out_33_39, out_33_40, out_33_41, out_33_42, out_33_43, out_33_44, out_33_45, out_33_46, out_33_47, out_33_48, out_33_49, out_33_50, out_33_51, out_33_52, out_33_53, out_33_54, out_33_55, out_33_56, out_33_57, out_33_58, out_33_59, out_33_60, out_33_61, out_33_62, out_33_63, out_33_64, out_34_1, out_34_2, out_34_3, out_34_4, out_34_5, out_34_6, out_34_7, out_34_8, out_34_9, out_34_10, out_34_11, out_34_12, out_34_13, out_34_14, out_34_15, out_34_16, out_34_17, out_34_18, out_34_19, out_34_20, out_34_21, out_34_22, out_34_23, out_34_24, out_34_25, out_34_26, out_34_27, out_34_28, out_34_29, out_34_30, out_34_31, out_34_32, out_34_33, out_34_34, out_34_35, out_34_36, out_34_37, out_34_38, out_34_39, out_34_40, out_34_41, out_34_42, out_34_43, out_34_44, out_34_45, out_34_46, out_34_47, out_34_48, out_34_49, out_34_50, out_34_51, out_34_52, out_34_53, out_34_54, out_34_55, out_34_56, out_34_57, out_34_58, out_34_59, out_34_60, out_34_61, out_34_62, out_34_63, out_34_64, out_35_1, out_35_2, out_35_3, out_35_4, out_35_5, out_35_6, out_35_7, out_35_8, out_35_9, out_35_10, out_35_11, out_35_12, out_35_13, out_35_14, out_35_15, out_35_16, out_35_17, out_35_18, out_35_19, out_35_20, out_35_21, out_35_22, out_35_23, out_35_24, out_35_25, out_35_26, out_35_27, out_35_28, out_35_29, out_35_30, out_35_31, out_35_32, out_35_33, out_35_34, out_35_35, out_35_36, out_35_37, out_35_38, out_35_39, out_35_40, out_35_41, out_35_42, out_35_43, out_35_44, out_35_45, out_35_46, out_35_47, out_35_48, out_35_49, out_35_50, out_35_51, out_35_52, out_35_53, out_35_54, out_35_55, out_35_56, out_35_57, out_35_58, out_35_59, out_35_60, out_35_61, out_35_62, out_35_63, out_35_64, out_36_1, out_36_2, out_36_3, out_36_4, out_36_5, out_36_6, out_36_7, out_36_8, out_36_9, out_36_10, out_36_11, out_36_12, out_36_13, out_36_14, out_36_15, out_36_16, out_36_17, out_36_18, out_36_19, out_36_20, out_36_21, out_36_22, out_36_23, out_36_24, out_36_25, out_36_26, out_36_27, out_36_28, out_36_29, out_36_30, out_36_31, out_36_32, out_36_33, out_36_34, out_36_35, out_36_36, out_36_37, out_36_38, out_36_39, out_36_40, out_36_41, out_36_42, out_36_43, out_36_44, out_36_45, out_36_46, out_36_47, out_36_48, out_36_49, out_36_50, out_36_51, out_36_52, out_36_53, out_36_54, out_36_55, out_36_56, out_36_57, out_36_58, out_36_59, out_36_60, out_36_61, out_36_62, out_36_63, out_36_64, out_37_1, out_37_2, out_37_3, out_37_4, out_37_5, out_37_6, out_37_7, out_37_8, out_37_9, out_37_10, out_37_11, out_37_12, out_37_13, out_37_14, out_37_15, out_37_16, out_37_17, out_37_18, out_37_19, out_37_20, out_37_21, out_37_22, out_37_23, out_37_24, out_37_25, out_37_26, out_37_27, out_37_28, out_37_29, out_37_30, out_37_31, out_37_32, out_37_33, out_37_34, out_37_35, out_37_36, out_37_37, out_37_38, out_37_39, out_37_40, out_37_41, out_37_42, out_37_43, out_37_44, out_37_45, out_37_46, out_37_47, out_37_48, out_37_49, out_37_50, out_37_51, out_37_52, out_37_53, out_37_54, out_37_55, out_37_56, out_37_57, out_37_58, out_37_59, out_37_60, out_37_61, out_37_62, out_37_63, out_37_64, out_38_1, out_38_2, out_38_3, out_38_4, out_38_5, out_38_6, out_38_7, out_38_8, out_38_9, out_38_10, out_38_11, out_38_12, out_38_13, out_38_14, out_38_15, out_38_16, out_38_17, out_38_18, out_38_19, out_38_20, out_38_21, out_38_22, out_38_23, out_38_24, out_38_25, out_38_26, out_38_27, out_38_28, out_38_29, out_38_30, out_38_31, out_38_32, out_38_33, out_38_34, out_38_35, out_38_36, out_38_37, out_38_38, out_38_39, out_38_40, out_38_41, out_38_42, out_38_43, out_38_44, out_38_45, out_38_46, out_38_47, out_38_48, out_38_49, out_38_50, out_38_51, out_38_52, out_38_53, out_38_54, out_38_55, out_38_56, out_38_57, out_38_58, out_38_59, out_38_60, out_38_61, out_38_62, out_38_63, out_38_64, out_39_1, out_39_2, out_39_3, out_39_4, out_39_5, out_39_6, out_39_7, out_39_8, out_39_9, out_39_10, out_39_11, out_39_12, out_39_13, out_39_14, out_39_15, out_39_16, out_39_17, out_39_18, out_39_19, out_39_20, out_39_21, out_39_22, out_39_23, out_39_24, out_39_25, out_39_26, out_39_27, out_39_28, out_39_29, out_39_30, out_39_31, out_39_32, out_39_33, out_39_34, out_39_35, out_39_36, out_39_37, out_39_38, out_39_39, out_39_40, out_39_41, out_39_42, out_39_43, out_39_44, out_39_45, out_39_46, out_39_47, out_39_48, out_39_49, out_39_50, out_39_51, out_39_52, out_39_53, out_39_54, out_39_55, out_39_56, out_39_57, out_39_58, out_39_59, out_39_60, out_39_61, out_39_62, out_39_63, out_39_64, out_40_1, out_40_2, out_40_3, out_40_4, out_40_5, out_40_6, out_40_7, out_40_8, out_40_9, out_40_10, out_40_11, out_40_12, out_40_13, out_40_14, out_40_15, out_40_16, out_40_17, out_40_18, out_40_19, out_40_20, out_40_21, out_40_22, out_40_23, out_40_24, out_40_25, out_40_26, out_40_27, out_40_28, out_40_29, out_40_30, out_40_31, out_40_32, out_40_33, out_40_34, out_40_35, out_40_36, out_40_37, out_40_38, out_40_39, out_40_40, out_40_41, out_40_42, out_40_43, out_40_44, out_40_45, out_40_46, out_40_47, out_40_48, out_40_49, out_40_50, out_40_51, out_40_52, out_40_53, out_40_54, out_40_55, out_40_56, out_40_57, out_40_58, out_40_59, out_40_60, out_40_61, out_40_62, out_40_63, out_40_64, out_41_1, out_41_2, out_41_3, out_41_4, out_41_5, out_41_6, out_41_7, out_41_8, out_41_9, out_41_10, out_41_11, out_41_12, out_41_13, out_41_14, out_41_15, out_41_16, out_41_17, out_41_18, out_41_19, out_41_20, out_41_21, out_41_22, out_41_23, out_41_24, out_41_25, out_41_26, out_41_27, out_41_28, out_41_29, out_41_30, out_41_31, out_41_32, out_41_33, out_41_34, out_41_35, out_41_36, out_41_37, out_41_38, out_41_39, out_41_40, out_41_41, out_41_42, out_41_43, out_41_44, out_41_45, out_41_46, out_41_47, out_41_48, out_41_49, out_41_50, out_41_51, out_41_52, out_41_53, out_41_54, out_41_55, out_41_56, out_41_57, out_41_58, out_41_59, out_41_60, out_41_61, out_41_62, out_41_63, out_41_64, out_42_1, out_42_2, out_42_3, out_42_4, out_42_5, out_42_6, out_42_7, out_42_8, out_42_9, out_42_10, out_42_11, out_42_12, out_42_13, out_42_14, out_42_15, out_42_16, out_42_17, out_42_18, out_42_19, out_42_20, out_42_21, out_42_22, out_42_23, out_42_24, out_42_25, out_42_26, out_42_27, out_42_28, out_42_29, out_42_30, out_42_31, out_42_32, out_42_33, out_42_34, out_42_35, out_42_36, out_42_37, out_42_38, out_42_39, out_42_40, out_42_41, out_42_42, out_42_43, out_42_44, out_42_45, out_42_46, out_42_47, out_42_48, out_42_49, out_42_50, out_42_51, out_42_52, out_42_53, out_42_54, out_42_55, out_42_56, out_42_57, out_42_58, out_42_59, out_42_60, out_42_61, out_42_62, out_42_63, out_42_64, out_43_1, out_43_2, out_43_3, out_43_4, out_43_5, out_43_6, out_43_7, out_43_8, out_43_9, out_43_10, out_43_11, out_43_12, out_43_13, out_43_14, out_43_15, out_43_16, out_43_17, out_43_18, out_43_19, out_43_20, out_43_21, out_43_22, out_43_23, out_43_24, out_43_25, out_43_26, out_43_27, out_43_28, out_43_29, out_43_30, out_43_31, out_43_32, out_43_33, out_43_34, out_43_35, out_43_36, out_43_37, out_43_38, out_43_39, out_43_40, out_43_41, out_43_42, out_43_43, out_43_44, out_43_45, out_43_46, out_43_47, out_43_48, out_43_49, out_43_50, out_43_51, out_43_52, out_43_53, out_43_54, out_43_55, out_43_56, out_43_57, out_43_58, out_43_59, out_43_60, out_43_61, out_43_62, out_43_63, out_43_64);

  input [7:0] p_0_0;
  input [7:0] p_0_1;
  input [7:0] p_0_2;
  input [7:0] p_0_3;
  input [7:0] p_0_4;
  input [7:0] p_0_5;
  input [7:0] p_0_6;
  input [7:0] p_0_7;
  input [7:0] p_0_8;
  input [7:0] p_0_9;
  input [7:0] p_0_10;
  input [7:0] p_0_11;
  input [7:0] p_0_12;
  input [7:0] p_0_13;
  input [7:0] p_0_14;
  input [7:0] p_0_15;
  input [7:0] p_0_16;
  input [7:0] p_0_17;
  input [7:0] p_0_18;
  input [7:0] p_0_19;
  input [7:0] p_0_20;
  input [7:0] p_0_21;
  input [7:0] p_0_22;
  input [7:0] p_0_23;
  input [7:0] p_0_24;
  input [7:0] p_0_25;
  input [7:0] p_0_26;
  input [7:0] p_0_27;
  input [7:0] p_0_28;
  input [7:0] p_0_29;
  input [7:0] p_0_30;
  input [7:0] p_0_31;
  input [7:0] p_0_32;
  input [7:0] p_0_33;
  input [7:0] p_0_34;
  input [7:0] p_0_35;
  input [7:0] p_0_36;
  input [7:0] p_0_37;
  input [7:0] p_0_38;
  input [7:0] p_0_39;
  input [7:0] p_0_40;
  input [7:0] p_0_41;
  input [7:0] p_0_42;
  input [7:0] p_0_43;
  input [7:0] p_0_44;
  input [7:0] p_0_45;
  input [7:0] p_0_46;
  input [7:0] p_0_47;
  input [7:0] p_0_48;
  input [7:0] p_0_49;
  input [7:0] p_0_50;
  input [7:0] p_0_51;
  input [7:0] p_0_52;
  input [7:0] p_0_53;
  input [7:0] p_0_54;
  input [7:0] p_0_55;
  input [7:0] p_0_56;
  input [7:0] p_0_57;
  input [7:0] p_0_58;
  input [7:0] p_0_59;
  input [7:0] p_0_60;
  input [7:0] p_0_61;
  input [7:0] p_0_62;
  input [7:0] p_0_63;
  input [7:0] p_0_64;
  input [7:0] p_0_65;
  input [7:0] p_1_0;
  input [7:0] p_1_1;
  input [7:0] p_1_2;
  input [7:0] p_1_3;
  input [7:0] p_1_4;
  input [7:0] p_1_5;
  input [7:0] p_1_6;
  input [7:0] p_1_7;
  input [7:0] p_1_8;
  input [7:0] p_1_9;
  input [7:0] p_1_10;
  input [7:0] p_1_11;
  input [7:0] p_1_12;
  input [7:0] p_1_13;
  input [7:0] p_1_14;
  input [7:0] p_1_15;
  input [7:0] p_1_16;
  input [7:0] p_1_17;
  input [7:0] p_1_18;
  input [7:0] p_1_19;
  input [7:0] p_1_20;
  input [7:0] p_1_21;
  input [7:0] p_1_22;
  input [7:0] p_1_23;
  input [7:0] p_1_24;
  input [7:0] p_1_25;
  input [7:0] p_1_26;
  input [7:0] p_1_27;
  input [7:0] p_1_28;
  input [7:0] p_1_29;
  input [7:0] p_1_30;
  input [7:0] p_1_31;
  input [7:0] p_1_32;
  input [7:0] p_1_33;
  input [7:0] p_1_34;
  input [7:0] p_1_35;
  input [7:0] p_1_36;
  input [7:0] p_1_37;
  input [7:0] p_1_38;
  input [7:0] p_1_39;
  input [7:0] p_1_40;
  input [7:0] p_1_41;
  input [7:0] p_1_42;
  input [7:0] p_1_43;
  input [7:0] p_1_44;
  input [7:0] p_1_45;
  input [7:0] p_1_46;
  input [7:0] p_1_47;
  input [7:0] p_1_48;
  input [7:0] p_1_49;
  input [7:0] p_1_50;
  input [7:0] p_1_51;
  input [7:0] p_1_52;
  input [7:0] p_1_53;
  input [7:0] p_1_54;
  input [7:0] p_1_55;
  input [7:0] p_1_56;
  input [7:0] p_1_57;
  input [7:0] p_1_58;
  input [7:0] p_1_59;
  input [7:0] p_1_60;
  input [7:0] p_1_61;
  input [7:0] p_1_62;
  input [7:0] p_1_63;
  input [7:0] p_1_64;
  input [7:0] p_1_65;
  input [7:0] p_2_0;
  input [7:0] p_2_1;
  input [7:0] p_2_2;
  input [7:0] p_2_3;
  input [7:0] p_2_4;
  input [7:0] p_2_5;
  input [7:0] p_2_6;
  input [7:0] p_2_7;
  input [7:0] p_2_8;
  input [7:0] p_2_9;
  input [7:0] p_2_10;
  input [7:0] p_2_11;
  input [7:0] p_2_12;
  input [7:0] p_2_13;
  input [7:0] p_2_14;
  input [7:0] p_2_15;
  input [7:0] p_2_16;
  input [7:0] p_2_17;
  input [7:0] p_2_18;
  input [7:0] p_2_19;
  input [7:0] p_2_20;
  input [7:0] p_2_21;
  input [7:0] p_2_22;
  input [7:0] p_2_23;
  input [7:0] p_2_24;
  input [7:0] p_2_25;
  input [7:0] p_2_26;
  input [7:0] p_2_27;
  input [7:0] p_2_28;
  input [7:0] p_2_29;
  input [7:0] p_2_30;
  input [7:0] p_2_31;
  input [7:0] p_2_32;
  input [7:0] p_2_33;
  input [7:0] p_2_34;
  input [7:0] p_2_35;
  input [7:0] p_2_36;
  input [7:0] p_2_37;
  input [7:0] p_2_38;
  input [7:0] p_2_39;
  input [7:0] p_2_40;
  input [7:0] p_2_41;
  input [7:0] p_2_42;
  input [7:0] p_2_43;
  input [7:0] p_2_44;
  input [7:0] p_2_45;
  input [7:0] p_2_46;
  input [7:0] p_2_47;
  input [7:0] p_2_48;
  input [7:0] p_2_49;
  input [7:0] p_2_50;
  input [7:0] p_2_51;
  input [7:0] p_2_52;
  input [7:0] p_2_53;
  input [7:0] p_2_54;
  input [7:0] p_2_55;
  input [7:0] p_2_56;
  input [7:0] p_2_57;
  input [7:0] p_2_58;
  input [7:0] p_2_59;
  input [7:0] p_2_60;
  input [7:0] p_2_61;
  input [7:0] p_2_62;
  input [7:0] p_2_63;
  input [7:0] p_2_64;
  input [7:0] p_2_65;
  input [7:0] p_3_0;
  input [7:0] p_3_1;
  input [7:0] p_3_2;
  input [7:0] p_3_3;
  input [7:0] p_3_4;
  input [7:0] p_3_5;
  input [7:0] p_3_6;
  input [7:0] p_3_7;
  input [7:0] p_3_8;
  input [7:0] p_3_9;
  input [7:0] p_3_10;
  input [7:0] p_3_11;
  input [7:0] p_3_12;
  input [7:0] p_3_13;
  input [7:0] p_3_14;
  input [7:0] p_3_15;
  input [7:0] p_3_16;
  input [7:0] p_3_17;
  input [7:0] p_3_18;
  input [7:0] p_3_19;
  input [7:0] p_3_20;
  input [7:0] p_3_21;
  input [7:0] p_3_22;
  input [7:0] p_3_23;
  input [7:0] p_3_24;
  input [7:0] p_3_25;
  input [7:0] p_3_26;
  input [7:0] p_3_27;
  input [7:0] p_3_28;
  input [7:0] p_3_29;
  input [7:0] p_3_30;
  input [7:0] p_3_31;
  input [7:0] p_3_32;
  input [7:0] p_3_33;
  input [7:0] p_3_34;
  input [7:0] p_3_35;
  input [7:0] p_3_36;
  input [7:0] p_3_37;
  input [7:0] p_3_38;
  input [7:0] p_3_39;
  input [7:0] p_3_40;
  input [7:0] p_3_41;
  input [7:0] p_3_42;
  input [7:0] p_3_43;
  input [7:0] p_3_44;
  input [7:0] p_3_45;
  input [7:0] p_3_46;
  input [7:0] p_3_47;
  input [7:0] p_3_48;
  input [7:0] p_3_49;
  input [7:0] p_3_50;
  input [7:0] p_3_51;
  input [7:0] p_3_52;
  input [7:0] p_3_53;
  input [7:0] p_3_54;
  input [7:0] p_3_55;
  input [7:0] p_3_56;
  input [7:0] p_3_57;
  input [7:0] p_3_58;
  input [7:0] p_3_59;
  input [7:0] p_3_60;
  input [7:0] p_3_61;
  input [7:0] p_3_62;
  input [7:0] p_3_63;
  input [7:0] p_3_64;
  input [7:0] p_3_65;
  input [7:0] p_4_0;
  input [7:0] p_4_1;
  input [7:0] p_4_2;
  input [7:0] p_4_3;
  input [7:0] p_4_4;
  input [7:0] p_4_5;
  input [7:0] p_4_6;
  input [7:0] p_4_7;
  input [7:0] p_4_8;
  input [7:0] p_4_9;
  input [7:0] p_4_10;
  input [7:0] p_4_11;
  input [7:0] p_4_12;
  input [7:0] p_4_13;
  input [7:0] p_4_14;
  input [7:0] p_4_15;
  input [7:0] p_4_16;
  input [7:0] p_4_17;
  input [7:0] p_4_18;
  input [7:0] p_4_19;
  input [7:0] p_4_20;
  input [7:0] p_4_21;
  input [7:0] p_4_22;
  input [7:0] p_4_23;
  input [7:0] p_4_24;
  input [7:0] p_4_25;
  input [7:0] p_4_26;
  input [7:0] p_4_27;
  input [7:0] p_4_28;
  input [7:0] p_4_29;
  input [7:0] p_4_30;
  input [7:0] p_4_31;
  input [7:0] p_4_32;
  input [7:0] p_4_33;
  input [7:0] p_4_34;
  input [7:0] p_4_35;
  input [7:0] p_4_36;
  input [7:0] p_4_37;
  input [7:0] p_4_38;
  input [7:0] p_4_39;
  input [7:0] p_4_40;
  input [7:0] p_4_41;
  input [7:0] p_4_42;
  input [7:0] p_4_43;
  input [7:0] p_4_44;
  input [7:0] p_4_45;
  input [7:0] p_4_46;
  input [7:0] p_4_47;
  input [7:0] p_4_48;
  input [7:0] p_4_49;
  input [7:0] p_4_50;
  input [7:0] p_4_51;
  input [7:0] p_4_52;
  input [7:0] p_4_53;
  input [7:0] p_4_54;
  input [7:0] p_4_55;
  input [7:0] p_4_56;
  input [7:0] p_4_57;
  input [7:0] p_4_58;
  input [7:0] p_4_59;
  input [7:0] p_4_60;
  input [7:0] p_4_61;
  input [7:0] p_4_62;
  input [7:0] p_4_63;
  input [7:0] p_4_64;
  input [7:0] p_4_65;
  input [7:0] p_5_0;
  input [7:0] p_5_1;
  input [7:0] p_5_2;
  input [7:0] p_5_3;
  input [7:0] p_5_4;
  input [7:0] p_5_5;
  input [7:0] p_5_6;
  input [7:0] p_5_7;
  input [7:0] p_5_8;
  input [7:0] p_5_9;
  input [7:0] p_5_10;
  input [7:0] p_5_11;
  input [7:0] p_5_12;
  input [7:0] p_5_13;
  input [7:0] p_5_14;
  input [7:0] p_5_15;
  input [7:0] p_5_16;
  input [7:0] p_5_17;
  input [7:0] p_5_18;
  input [7:0] p_5_19;
  input [7:0] p_5_20;
  input [7:0] p_5_21;
  input [7:0] p_5_22;
  input [7:0] p_5_23;
  input [7:0] p_5_24;
  input [7:0] p_5_25;
  input [7:0] p_5_26;
  input [7:0] p_5_27;
  input [7:0] p_5_28;
  input [7:0] p_5_29;
  input [7:0] p_5_30;
  input [7:0] p_5_31;
  input [7:0] p_5_32;
  input [7:0] p_5_33;
  input [7:0] p_5_34;
  input [7:0] p_5_35;
  input [7:0] p_5_36;
  input [7:0] p_5_37;
  input [7:0] p_5_38;
  input [7:0] p_5_39;
  input [7:0] p_5_40;
  input [7:0] p_5_41;
  input [7:0] p_5_42;
  input [7:0] p_5_43;
  input [7:0] p_5_44;
  input [7:0] p_5_45;
  input [7:0] p_5_46;
  input [7:0] p_5_47;
  input [7:0] p_5_48;
  input [7:0] p_5_49;
  input [7:0] p_5_50;
  input [7:0] p_5_51;
  input [7:0] p_5_52;
  input [7:0] p_5_53;
  input [7:0] p_5_54;
  input [7:0] p_5_55;
  input [7:0] p_5_56;
  input [7:0] p_5_57;
  input [7:0] p_5_58;
  input [7:0] p_5_59;
  input [7:0] p_5_60;
  input [7:0] p_5_61;
  input [7:0] p_5_62;
  input [7:0] p_5_63;
  input [7:0] p_5_64;
  input [7:0] p_5_65;
  input [7:0] p_6_0;
  input [7:0] p_6_1;
  input [7:0] p_6_2;
  input [7:0] p_6_3;
  input [7:0] p_6_4;
  input [7:0] p_6_5;
  input [7:0] p_6_6;
  input [7:0] p_6_7;
  input [7:0] p_6_8;
  input [7:0] p_6_9;
  input [7:0] p_6_10;
  input [7:0] p_6_11;
  input [7:0] p_6_12;
  input [7:0] p_6_13;
  input [7:0] p_6_14;
  input [7:0] p_6_15;
  input [7:0] p_6_16;
  input [7:0] p_6_17;
  input [7:0] p_6_18;
  input [7:0] p_6_19;
  input [7:0] p_6_20;
  input [7:0] p_6_21;
  input [7:0] p_6_22;
  input [7:0] p_6_23;
  input [7:0] p_6_24;
  input [7:0] p_6_25;
  input [7:0] p_6_26;
  input [7:0] p_6_27;
  input [7:0] p_6_28;
  input [7:0] p_6_29;
  input [7:0] p_6_30;
  input [7:0] p_6_31;
  input [7:0] p_6_32;
  input [7:0] p_6_33;
  input [7:0] p_6_34;
  input [7:0] p_6_35;
  input [7:0] p_6_36;
  input [7:0] p_6_37;
  input [7:0] p_6_38;
  input [7:0] p_6_39;
  input [7:0] p_6_40;
  input [7:0] p_6_41;
  input [7:0] p_6_42;
  input [7:0] p_6_43;
  input [7:0] p_6_44;
  input [7:0] p_6_45;
  input [7:0] p_6_46;
  input [7:0] p_6_47;
  input [7:0] p_6_48;
  input [7:0] p_6_49;
  input [7:0] p_6_50;
  input [7:0] p_6_51;
  input [7:0] p_6_52;
  input [7:0] p_6_53;
  input [7:0] p_6_54;
  input [7:0] p_6_55;
  input [7:0] p_6_56;
  input [7:0] p_6_57;
  input [7:0] p_6_58;
  input [7:0] p_6_59;
  input [7:0] p_6_60;
  input [7:0] p_6_61;
  input [7:0] p_6_62;
  input [7:0] p_6_63;
  input [7:0] p_6_64;
  input [7:0] p_6_65;
  input [7:0] p_7_0;
  input [7:0] p_7_1;
  input [7:0] p_7_2;
  input [7:0] p_7_3;
  input [7:0] p_7_4;
  input [7:0] p_7_5;
  input [7:0] p_7_6;
  input [7:0] p_7_7;
  input [7:0] p_7_8;
  input [7:0] p_7_9;
  input [7:0] p_7_10;
  input [7:0] p_7_11;
  input [7:0] p_7_12;
  input [7:0] p_7_13;
  input [7:0] p_7_14;
  input [7:0] p_7_15;
  input [7:0] p_7_16;
  input [7:0] p_7_17;
  input [7:0] p_7_18;
  input [7:0] p_7_19;
  input [7:0] p_7_20;
  input [7:0] p_7_21;
  input [7:0] p_7_22;
  input [7:0] p_7_23;
  input [7:0] p_7_24;
  input [7:0] p_7_25;
  input [7:0] p_7_26;
  input [7:0] p_7_27;
  input [7:0] p_7_28;
  input [7:0] p_7_29;
  input [7:0] p_7_30;
  input [7:0] p_7_31;
  input [7:0] p_7_32;
  input [7:0] p_7_33;
  input [7:0] p_7_34;
  input [7:0] p_7_35;
  input [7:0] p_7_36;
  input [7:0] p_7_37;
  input [7:0] p_7_38;
  input [7:0] p_7_39;
  input [7:0] p_7_40;
  input [7:0] p_7_41;
  input [7:0] p_7_42;
  input [7:0] p_7_43;
  input [7:0] p_7_44;
  input [7:0] p_7_45;
  input [7:0] p_7_46;
  input [7:0] p_7_47;
  input [7:0] p_7_48;
  input [7:0] p_7_49;
  input [7:0] p_7_50;
  input [7:0] p_7_51;
  input [7:0] p_7_52;
  input [7:0] p_7_53;
  input [7:0] p_7_54;
  input [7:0] p_7_55;
  input [7:0] p_7_56;
  input [7:0] p_7_57;
  input [7:0] p_7_58;
  input [7:0] p_7_59;
  input [7:0] p_7_60;
  input [7:0] p_7_61;
  input [7:0] p_7_62;
  input [7:0] p_7_63;
  input [7:0] p_7_64;
  input [7:0] p_7_65;
  input [7:0] p_8_0;
  input [7:0] p_8_1;
  input [7:0] p_8_2;
  input [7:0] p_8_3;
  input [7:0] p_8_4;
  input [7:0] p_8_5;
  input [7:0] p_8_6;
  input [7:0] p_8_7;
  input [7:0] p_8_8;
  input [7:0] p_8_9;
  input [7:0] p_8_10;
  input [7:0] p_8_11;
  input [7:0] p_8_12;
  input [7:0] p_8_13;
  input [7:0] p_8_14;
  input [7:0] p_8_15;
  input [7:0] p_8_16;
  input [7:0] p_8_17;
  input [7:0] p_8_18;
  input [7:0] p_8_19;
  input [7:0] p_8_20;
  input [7:0] p_8_21;
  input [7:0] p_8_22;
  input [7:0] p_8_23;
  input [7:0] p_8_24;
  input [7:0] p_8_25;
  input [7:0] p_8_26;
  input [7:0] p_8_27;
  input [7:0] p_8_28;
  input [7:0] p_8_29;
  input [7:0] p_8_30;
  input [7:0] p_8_31;
  input [7:0] p_8_32;
  input [7:0] p_8_33;
  input [7:0] p_8_34;
  input [7:0] p_8_35;
  input [7:0] p_8_36;
  input [7:0] p_8_37;
  input [7:0] p_8_38;
  input [7:0] p_8_39;
  input [7:0] p_8_40;
  input [7:0] p_8_41;
  input [7:0] p_8_42;
  input [7:0] p_8_43;
  input [7:0] p_8_44;
  input [7:0] p_8_45;
  input [7:0] p_8_46;
  input [7:0] p_8_47;
  input [7:0] p_8_48;
  input [7:0] p_8_49;
  input [7:0] p_8_50;
  input [7:0] p_8_51;
  input [7:0] p_8_52;
  input [7:0] p_8_53;
  input [7:0] p_8_54;
  input [7:0] p_8_55;
  input [7:0] p_8_56;
  input [7:0] p_8_57;
  input [7:0] p_8_58;
  input [7:0] p_8_59;
  input [7:0] p_8_60;
  input [7:0] p_8_61;
  input [7:0] p_8_62;
  input [7:0] p_8_63;
  input [7:0] p_8_64;
  input [7:0] p_8_65;
  input [7:0] p_9_0;
  input [7:0] p_9_1;
  input [7:0] p_9_2;
  input [7:0] p_9_3;
  input [7:0] p_9_4;
  input [7:0] p_9_5;
  input [7:0] p_9_6;
  input [7:0] p_9_7;
  input [7:0] p_9_8;
  input [7:0] p_9_9;
  input [7:0] p_9_10;
  input [7:0] p_9_11;
  input [7:0] p_9_12;
  input [7:0] p_9_13;
  input [7:0] p_9_14;
  input [7:0] p_9_15;
  input [7:0] p_9_16;
  input [7:0] p_9_17;
  input [7:0] p_9_18;
  input [7:0] p_9_19;
  input [7:0] p_9_20;
  input [7:0] p_9_21;
  input [7:0] p_9_22;
  input [7:0] p_9_23;
  input [7:0] p_9_24;
  input [7:0] p_9_25;
  input [7:0] p_9_26;
  input [7:0] p_9_27;
  input [7:0] p_9_28;
  input [7:0] p_9_29;
  input [7:0] p_9_30;
  input [7:0] p_9_31;
  input [7:0] p_9_32;
  input [7:0] p_9_33;
  input [7:0] p_9_34;
  input [7:0] p_9_35;
  input [7:0] p_9_36;
  input [7:0] p_9_37;
  input [7:0] p_9_38;
  input [7:0] p_9_39;
  input [7:0] p_9_40;
  input [7:0] p_9_41;
  input [7:0] p_9_42;
  input [7:0] p_9_43;
  input [7:0] p_9_44;
  input [7:0] p_9_45;
  input [7:0] p_9_46;
  input [7:0] p_9_47;
  input [7:0] p_9_48;
  input [7:0] p_9_49;
  input [7:0] p_9_50;
  input [7:0] p_9_51;
  input [7:0] p_9_52;
  input [7:0] p_9_53;
  input [7:0] p_9_54;
  input [7:0] p_9_55;
  input [7:0] p_9_56;
  input [7:0] p_9_57;
  input [7:0] p_9_58;
  input [7:0] p_9_59;
  input [7:0] p_9_60;
  input [7:0] p_9_61;
  input [7:0] p_9_62;
  input [7:0] p_9_63;
  input [7:0] p_9_64;
  input [7:0] p_9_65;
  input [7:0] p_10_0;
  input [7:0] p_10_1;
  input [7:0] p_10_2;
  input [7:0] p_10_3;
  input [7:0] p_10_4;
  input [7:0] p_10_5;
  input [7:0] p_10_6;
  input [7:0] p_10_7;
  input [7:0] p_10_8;
  input [7:0] p_10_9;
  input [7:0] p_10_10;
  input [7:0] p_10_11;
  input [7:0] p_10_12;
  input [7:0] p_10_13;
  input [7:0] p_10_14;
  input [7:0] p_10_15;
  input [7:0] p_10_16;
  input [7:0] p_10_17;
  input [7:0] p_10_18;
  input [7:0] p_10_19;
  input [7:0] p_10_20;
  input [7:0] p_10_21;
  input [7:0] p_10_22;
  input [7:0] p_10_23;
  input [7:0] p_10_24;
  input [7:0] p_10_25;
  input [7:0] p_10_26;
  input [7:0] p_10_27;
  input [7:0] p_10_28;
  input [7:0] p_10_29;
  input [7:0] p_10_30;
  input [7:0] p_10_31;
  input [7:0] p_10_32;
  input [7:0] p_10_33;
  input [7:0] p_10_34;
  input [7:0] p_10_35;
  input [7:0] p_10_36;
  input [7:0] p_10_37;
  input [7:0] p_10_38;
  input [7:0] p_10_39;
  input [7:0] p_10_40;
  input [7:0] p_10_41;
  input [7:0] p_10_42;
  input [7:0] p_10_43;
  input [7:0] p_10_44;
  input [7:0] p_10_45;
  input [7:0] p_10_46;
  input [7:0] p_10_47;
  input [7:0] p_10_48;
  input [7:0] p_10_49;
  input [7:0] p_10_50;
  input [7:0] p_10_51;
  input [7:0] p_10_52;
  input [7:0] p_10_53;
  input [7:0] p_10_54;
  input [7:0] p_10_55;
  input [7:0] p_10_56;
  input [7:0] p_10_57;
  input [7:0] p_10_58;
  input [7:0] p_10_59;
  input [7:0] p_10_60;
  input [7:0] p_10_61;
  input [7:0] p_10_62;
  input [7:0] p_10_63;
  input [7:0] p_10_64;
  input [7:0] p_10_65;
  input [7:0] p_11_0;
  input [7:0] p_11_1;
  input [7:0] p_11_2;
  input [7:0] p_11_3;
  input [7:0] p_11_4;
  input [7:0] p_11_5;
  input [7:0] p_11_6;
  input [7:0] p_11_7;
  input [7:0] p_11_8;
  input [7:0] p_11_9;
  input [7:0] p_11_10;
  input [7:0] p_11_11;
  input [7:0] p_11_12;
  input [7:0] p_11_13;
  input [7:0] p_11_14;
  input [7:0] p_11_15;
  input [7:0] p_11_16;
  input [7:0] p_11_17;
  input [7:0] p_11_18;
  input [7:0] p_11_19;
  input [7:0] p_11_20;
  input [7:0] p_11_21;
  input [7:0] p_11_22;
  input [7:0] p_11_23;
  input [7:0] p_11_24;
  input [7:0] p_11_25;
  input [7:0] p_11_26;
  input [7:0] p_11_27;
  input [7:0] p_11_28;
  input [7:0] p_11_29;
  input [7:0] p_11_30;
  input [7:0] p_11_31;
  input [7:0] p_11_32;
  input [7:0] p_11_33;
  input [7:0] p_11_34;
  input [7:0] p_11_35;
  input [7:0] p_11_36;
  input [7:0] p_11_37;
  input [7:0] p_11_38;
  input [7:0] p_11_39;
  input [7:0] p_11_40;
  input [7:0] p_11_41;
  input [7:0] p_11_42;
  input [7:0] p_11_43;
  input [7:0] p_11_44;
  input [7:0] p_11_45;
  input [7:0] p_11_46;
  input [7:0] p_11_47;
  input [7:0] p_11_48;
  input [7:0] p_11_49;
  input [7:0] p_11_50;
  input [7:0] p_11_51;
  input [7:0] p_11_52;
  input [7:0] p_11_53;
  input [7:0] p_11_54;
  input [7:0] p_11_55;
  input [7:0] p_11_56;
  input [7:0] p_11_57;
  input [7:0] p_11_58;
  input [7:0] p_11_59;
  input [7:0] p_11_60;
  input [7:0] p_11_61;
  input [7:0] p_11_62;
  input [7:0] p_11_63;
  input [7:0] p_11_64;
  input [7:0] p_11_65;
  input [7:0] p_12_0;
  input [7:0] p_12_1;
  input [7:0] p_12_2;
  input [7:0] p_12_3;
  input [7:0] p_12_4;
  input [7:0] p_12_5;
  input [7:0] p_12_6;
  input [7:0] p_12_7;
  input [7:0] p_12_8;
  input [7:0] p_12_9;
  input [7:0] p_12_10;
  input [7:0] p_12_11;
  input [7:0] p_12_12;
  input [7:0] p_12_13;
  input [7:0] p_12_14;
  input [7:0] p_12_15;
  input [7:0] p_12_16;
  input [7:0] p_12_17;
  input [7:0] p_12_18;
  input [7:0] p_12_19;
  input [7:0] p_12_20;
  input [7:0] p_12_21;
  input [7:0] p_12_22;
  input [7:0] p_12_23;
  input [7:0] p_12_24;
  input [7:0] p_12_25;
  input [7:0] p_12_26;
  input [7:0] p_12_27;
  input [7:0] p_12_28;
  input [7:0] p_12_29;
  input [7:0] p_12_30;
  input [7:0] p_12_31;
  input [7:0] p_12_32;
  input [7:0] p_12_33;
  input [7:0] p_12_34;
  input [7:0] p_12_35;
  input [7:0] p_12_36;
  input [7:0] p_12_37;
  input [7:0] p_12_38;
  input [7:0] p_12_39;
  input [7:0] p_12_40;
  input [7:0] p_12_41;
  input [7:0] p_12_42;
  input [7:0] p_12_43;
  input [7:0] p_12_44;
  input [7:0] p_12_45;
  input [7:0] p_12_46;
  input [7:0] p_12_47;
  input [7:0] p_12_48;
  input [7:0] p_12_49;
  input [7:0] p_12_50;
  input [7:0] p_12_51;
  input [7:0] p_12_52;
  input [7:0] p_12_53;
  input [7:0] p_12_54;
  input [7:0] p_12_55;
  input [7:0] p_12_56;
  input [7:0] p_12_57;
  input [7:0] p_12_58;
  input [7:0] p_12_59;
  input [7:0] p_12_60;
  input [7:0] p_12_61;
  input [7:0] p_12_62;
  input [7:0] p_12_63;
  input [7:0] p_12_64;
  input [7:0] p_12_65;
  input [7:0] p_13_0;
  input [7:0] p_13_1;
  input [7:0] p_13_2;
  input [7:0] p_13_3;
  input [7:0] p_13_4;
  input [7:0] p_13_5;
  input [7:0] p_13_6;
  input [7:0] p_13_7;
  input [7:0] p_13_8;
  input [7:0] p_13_9;
  input [7:0] p_13_10;
  input [7:0] p_13_11;
  input [7:0] p_13_12;
  input [7:0] p_13_13;
  input [7:0] p_13_14;
  input [7:0] p_13_15;
  input [7:0] p_13_16;
  input [7:0] p_13_17;
  input [7:0] p_13_18;
  input [7:0] p_13_19;
  input [7:0] p_13_20;
  input [7:0] p_13_21;
  input [7:0] p_13_22;
  input [7:0] p_13_23;
  input [7:0] p_13_24;
  input [7:0] p_13_25;
  input [7:0] p_13_26;
  input [7:0] p_13_27;
  input [7:0] p_13_28;
  input [7:0] p_13_29;
  input [7:0] p_13_30;
  input [7:0] p_13_31;
  input [7:0] p_13_32;
  input [7:0] p_13_33;
  input [7:0] p_13_34;
  input [7:0] p_13_35;
  input [7:0] p_13_36;
  input [7:0] p_13_37;
  input [7:0] p_13_38;
  input [7:0] p_13_39;
  input [7:0] p_13_40;
  input [7:0] p_13_41;
  input [7:0] p_13_42;
  input [7:0] p_13_43;
  input [7:0] p_13_44;
  input [7:0] p_13_45;
  input [7:0] p_13_46;
  input [7:0] p_13_47;
  input [7:0] p_13_48;
  input [7:0] p_13_49;
  input [7:0] p_13_50;
  input [7:0] p_13_51;
  input [7:0] p_13_52;
  input [7:0] p_13_53;
  input [7:0] p_13_54;
  input [7:0] p_13_55;
  input [7:0] p_13_56;
  input [7:0] p_13_57;
  input [7:0] p_13_58;
  input [7:0] p_13_59;
  input [7:0] p_13_60;
  input [7:0] p_13_61;
  input [7:0] p_13_62;
  input [7:0] p_13_63;
  input [7:0] p_13_64;
  input [7:0] p_13_65;
  input [7:0] p_14_0;
  input [7:0] p_14_1;
  input [7:0] p_14_2;
  input [7:0] p_14_3;
  input [7:0] p_14_4;
  input [7:0] p_14_5;
  input [7:0] p_14_6;
  input [7:0] p_14_7;
  input [7:0] p_14_8;
  input [7:0] p_14_9;
  input [7:0] p_14_10;
  input [7:0] p_14_11;
  input [7:0] p_14_12;
  input [7:0] p_14_13;
  input [7:0] p_14_14;
  input [7:0] p_14_15;
  input [7:0] p_14_16;
  input [7:0] p_14_17;
  input [7:0] p_14_18;
  input [7:0] p_14_19;
  input [7:0] p_14_20;
  input [7:0] p_14_21;
  input [7:0] p_14_22;
  input [7:0] p_14_23;
  input [7:0] p_14_24;
  input [7:0] p_14_25;
  input [7:0] p_14_26;
  input [7:0] p_14_27;
  input [7:0] p_14_28;
  input [7:0] p_14_29;
  input [7:0] p_14_30;
  input [7:0] p_14_31;
  input [7:0] p_14_32;
  input [7:0] p_14_33;
  input [7:0] p_14_34;
  input [7:0] p_14_35;
  input [7:0] p_14_36;
  input [7:0] p_14_37;
  input [7:0] p_14_38;
  input [7:0] p_14_39;
  input [7:0] p_14_40;
  input [7:0] p_14_41;
  input [7:0] p_14_42;
  input [7:0] p_14_43;
  input [7:0] p_14_44;
  input [7:0] p_14_45;
  input [7:0] p_14_46;
  input [7:0] p_14_47;
  input [7:0] p_14_48;
  input [7:0] p_14_49;
  input [7:0] p_14_50;
  input [7:0] p_14_51;
  input [7:0] p_14_52;
  input [7:0] p_14_53;
  input [7:0] p_14_54;
  input [7:0] p_14_55;
  input [7:0] p_14_56;
  input [7:0] p_14_57;
  input [7:0] p_14_58;
  input [7:0] p_14_59;
  input [7:0] p_14_60;
  input [7:0] p_14_61;
  input [7:0] p_14_62;
  input [7:0] p_14_63;
  input [7:0] p_14_64;
  input [7:0] p_14_65;
  input [7:0] p_15_0;
  input [7:0] p_15_1;
  input [7:0] p_15_2;
  input [7:0] p_15_3;
  input [7:0] p_15_4;
  input [7:0] p_15_5;
  input [7:0] p_15_6;
  input [7:0] p_15_7;
  input [7:0] p_15_8;
  input [7:0] p_15_9;
  input [7:0] p_15_10;
  input [7:0] p_15_11;
  input [7:0] p_15_12;
  input [7:0] p_15_13;
  input [7:0] p_15_14;
  input [7:0] p_15_15;
  input [7:0] p_15_16;
  input [7:0] p_15_17;
  input [7:0] p_15_18;
  input [7:0] p_15_19;
  input [7:0] p_15_20;
  input [7:0] p_15_21;
  input [7:0] p_15_22;
  input [7:0] p_15_23;
  input [7:0] p_15_24;
  input [7:0] p_15_25;
  input [7:0] p_15_26;
  input [7:0] p_15_27;
  input [7:0] p_15_28;
  input [7:0] p_15_29;
  input [7:0] p_15_30;
  input [7:0] p_15_31;
  input [7:0] p_15_32;
  input [7:0] p_15_33;
  input [7:0] p_15_34;
  input [7:0] p_15_35;
  input [7:0] p_15_36;
  input [7:0] p_15_37;
  input [7:0] p_15_38;
  input [7:0] p_15_39;
  input [7:0] p_15_40;
  input [7:0] p_15_41;
  input [7:0] p_15_42;
  input [7:0] p_15_43;
  input [7:0] p_15_44;
  input [7:0] p_15_45;
  input [7:0] p_15_46;
  input [7:0] p_15_47;
  input [7:0] p_15_48;
  input [7:0] p_15_49;
  input [7:0] p_15_50;
  input [7:0] p_15_51;
  input [7:0] p_15_52;
  input [7:0] p_15_53;
  input [7:0] p_15_54;
  input [7:0] p_15_55;
  input [7:0] p_15_56;
  input [7:0] p_15_57;
  input [7:0] p_15_58;
  input [7:0] p_15_59;
  input [7:0] p_15_60;
  input [7:0] p_15_61;
  input [7:0] p_15_62;
  input [7:0] p_15_63;
  input [7:0] p_15_64;
  input [7:0] p_15_65;
  input [7:0] p_16_0;
  input [7:0] p_16_1;
  input [7:0] p_16_2;
  input [7:0] p_16_3;
  input [7:0] p_16_4;
  input [7:0] p_16_5;
  input [7:0] p_16_6;
  input [7:0] p_16_7;
  input [7:0] p_16_8;
  input [7:0] p_16_9;
  input [7:0] p_16_10;
  input [7:0] p_16_11;
  input [7:0] p_16_12;
  input [7:0] p_16_13;
  input [7:0] p_16_14;
  input [7:0] p_16_15;
  input [7:0] p_16_16;
  input [7:0] p_16_17;
  input [7:0] p_16_18;
  input [7:0] p_16_19;
  input [7:0] p_16_20;
  input [7:0] p_16_21;
  input [7:0] p_16_22;
  input [7:0] p_16_23;
  input [7:0] p_16_24;
  input [7:0] p_16_25;
  input [7:0] p_16_26;
  input [7:0] p_16_27;
  input [7:0] p_16_28;
  input [7:0] p_16_29;
  input [7:0] p_16_30;
  input [7:0] p_16_31;
  input [7:0] p_16_32;
  input [7:0] p_16_33;
  input [7:0] p_16_34;
  input [7:0] p_16_35;
  input [7:0] p_16_36;
  input [7:0] p_16_37;
  input [7:0] p_16_38;
  input [7:0] p_16_39;
  input [7:0] p_16_40;
  input [7:0] p_16_41;
  input [7:0] p_16_42;
  input [7:0] p_16_43;
  input [7:0] p_16_44;
  input [7:0] p_16_45;
  input [7:0] p_16_46;
  input [7:0] p_16_47;
  input [7:0] p_16_48;
  input [7:0] p_16_49;
  input [7:0] p_16_50;
  input [7:0] p_16_51;
  input [7:0] p_16_52;
  input [7:0] p_16_53;
  input [7:0] p_16_54;
  input [7:0] p_16_55;
  input [7:0] p_16_56;
  input [7:0] p_16_57;
  input [7:0] p_16_58;
  input [7:0] p_16_59;
  input [7:0] p_16_60;
  input [7:0] p_16_61;
  input [7:0] p_16_62;
  input [7:0] p_16_63;
  input [7:0] p_16_64;
  input [7:0] p_16_65;
  input [7:0] p_17_0;
  input [7:0] p_17_1;
  input [7:0] p_17_2;
  input [7:0] p_17_3;
  input [7:0] p_17_4;
  input [7:0] p_17_5;
  input [7:0] p_17_6;
  input [7:0] p_17_7;
  input [7:0] p_17_8;
  input [7:0] p_17_9;
  input [7:0] p_17_10;
  input [7:0] p_17_11;
  input [7:0] p_17_12;
  input [7:0] p_17_13;
  input [7:0] p_17_14;
  input [7:0] p_17_15;
  input [7:0] p_17_16;
  input [7:0] p_17_17;
  input [7:0] p_17_18;
  input [7:0] p_17_19;
  input [7:0] p_17_20;
  input [7:0] p_17_21;
  input [7:0] p_17_22;
  input [7:0] p_17_23;
  input [7:0] p_17_24;
  input [7:0] p_17_25;
  input [7:0] p_17_26;
  input [7:0] p_17_27;
  input [7:0] p_17_28;
  input [7:0] p_17_29;
  input [7:0] p_17_30;
  input [7:0] p_17_31;
  input [7:0] p_17_32;
  input [7:0] p_17_33;
  input [7:0] p_17_34;
  input [7:0] p_17_35;
  input [7:0] p_17_36;
  input [7:0] p_17_37;
  input [7:0] p_17_38;
  input [7:0] p_17_39;
  input [7:0] p_17_40;
  input [7:0] p_17_41;
  input [7:0] p_17_42;
  input [7:0] p_17_43;
  input [7:0] p_17_44;
  input [7:0] p_17_45;
  input [7:0] p_17_46;
  input [7:0] p_17_47;
  input [7:0] p_17_48;
  input [7:0] p_17_49;
  input [7:0] p_17_50;
  input [7:0] p_17_51;
  input [7:0] p_17_52;
  input [7:0] p_17_53;
  input [7:0] p_17_54;
  input [7:0] p_17_55;
  input [7:0] p_17_56;
  input [7:0] p_17_57;
  input [7:0] p_17_58;
  input [7:0] p_17_59;
  input [7:0] p_17_60;
  input [7:0] p_17_61;
  input [7:0] p_17_62;
  input [7:0] p_17_63;
  input [7:0] p_17_64;
  input [7:0] p_17_65;
  input [7:0] p_18_0;
  input [7:0] p_18_1;
  input [7:0] p_18_2;
  input [7:0] p_18_3;
  input [7:0] p_18_4;
  input [7:0] p_18_5;
  input [7:0] p_18_6;
  input [7:0] p_18_7;
  input [7:0] p_18_8;
  input [7:0] p_18_9;
  input [7:0] p_18_10;
  input [7:0] p_18_11;
  input [7:0] p_18_12;
  input [7:0] p_18_13;
  input [7:0] p_18_14;
  input [7:0] p_18_15;
  input [7:0] p_18_16;
  input [7:0] p_18_17;
  input [7:0] p_18_18;
  input [7:0] p_18_19;
  input [7:0] p_18_20;
  input [7:0] p_18_21;
  input [7:0] p_18_22;
  input [7:0] p_18_23;
  input [7:0] p_18_24;
  input [7:0] p_18_25;
  input [7:0] p_18_26;
  input [7:0] p_18_27;
  input [7:0] p_18_28;
  input [7:0] p_18_29;
  input [7:0] p_18_30;
  input [7:0] p_18_31;
  input [7:0] p_18_32;
  input [7:0] p_18_33;
  input [7:0] p_18_34;
  input [7:0] p_18_35;
  input [7:0] p_18_36;
  input [7:0] p_18_37;
  input [7:0] p_18_38;
  input [7:0] p_18_39;
  input [7:0] p_18_40;
  input [7:0] p_18_41;
  input [7:0] p_18_42;
  input [7:0] p_18_43;
  input [7:0] p_18_44;
  input [7:0] p_18_45;
  input [7:0] p_18_46;
  input [7:0] p_18_47;
  input [7:0] p_18_48;
  input [7:0] p_18_49;
  input [7:0] p_18_50;
  input [7:0] p_18_51;
  input [7:0] p_18_52;
  input [7:0] p_18_53;
  input [7:0] p_18_54;
  input [7:0] p_18_55;
  input [7:0] p_18_56;
  input [7:0] p_18_57;
  input [7:0] p_18_58;
  input [7:0] p_18_59;
  input [7:0] p_18_60;
  input [7:0] p_18_61;
  input [7:0] p_18_62;
  input [7:0] p_18_63;
  input [7:0] p_18_64;
  input [7:0] p_18_65;
  input [7:0] p_19_0;
  input [7:0] p_19_1;
  input [7:0] p_19_2;
  input [7:0] p_19_3;
  input [7:0] p_19_4;
  input [7:0] p_19_5;
  input [7:0] p_19_6;
  input [7:0] p_19_7;
  input [7:0] p_19_8;
  input [7:0] p_19_9;
  input [7:0] p_19_10;
  input [7:0] p_19_11;
  input [7:0] p_19_12;
  input [7:0] p_19_13;
  input [7:0] p_19_14;
  input [7:0] p_19_15;
  input [7:0] p_19_16;
  input [7:0] p_19_17;
  input [7:0] p_19_18;
  input [7:0] p_19_19;
  input [7:0] p_19_20;
  input [7:0] p_19_21;
  input [7:0] p_19_22;
  input [7:0] p_19_23;
  input [7:0] p_19_24;
  input [7:0] p_19_25;
  input [7:0] p_19_26;
  input [7:0] p_19_27;
  input [7:0] p_19_28;
  input [7:0] p_19_29;
  input [7:0] p_19_30;
  input [7:0] p_19_31;
  input [7:0] p_19_32;
  input [7:0] p_19_33;
  input [7:0] p_19_34;
  input [7:0] p_19_35;
  input [7:0] p_19_36;
  input [7:0] p_19_37;
  input [7:0] p_19_38;
  input [7:0] p_19_39;
  input [7:0] p_19_40;
  input [7:0] p_19_41;
  input [7:0] p_19_42;
  input [7:0] p_19_43;
  input [7:0] p_19_44;
  input [7:0] p_19_45;
  input [7:0] p_19_46;
  input [7:0] p_19_47;
  input [7:0] p_19_48;
  input [7:0] p_19_49;
  input [7:0] p_19_50;
  input [7:0] p_19_51;
  input [7:0] p_19_52;
  input [7:0] p_19_53;
  input [7:0] p_19_54;
  input [7:0] p_19_55;
  input [7:0] p_19_56;
  input [7:0] p_19_57;
  input [7:0] p_19_58;
  input [7:0] p_19_59;
  input [7:0] p_19_60;
  input [7:0] p_19_61;
  input [7:0] p_19_62;
  input [7:0] p_19_63;
  input [7:0] p_19_64;
  input [7:0] p_19_65;
  input [7:0] p_20_0;
  input [7:0] p_20_1;
  input [7:0] p_20_2;
  input [7:0] p_20_3;
  input [7:0] p_20_4;
  input [7:0] p_20_5;
  input [7:0] p_20_6;
  input [7:0] p_20_7;
  input [7:0] p_20_8;
  input [7:0] p_20_9;
  input [7:0] p_20_10;
  input [7:0] p_20_11;
  input [7:0] p_20_12;
  input [7:0] p_20_13;
  input [7:0] p_20_14;
  input [7:0] p_20_15;
  input [7:0] p_20_16;
  input [7:0] p_20_17;
  input [7:0] p_20_18;
  input [7:0] p_20_19;
  input [7:0] p_20_20;
  input [7:0] p_20_21;
  input [7:0] p_20_22;
  input [7:0] p_20_23;
  input [7:0] p_20_24;
  input [7:0] p_20_25;
  input [7:0] p_20_26;
  input [7:0] p_20_27;
  input [7:0] p_20_28;
  input [7:0] p_20_29;
  input [7:0] p_20_30;
  input [7:0] p_20_31;
  input [7:0] p_20_32;
  input [7:0] p_20_33;
  input [7:0] p_20_34;
  input [7:0] p_20_35;
  input [7:0] p_20_36;
  input [7:0] p_20_37;
  input [7:0] p_20_38;
  input [7:0] p_20_39;
  input [7:0] p_20_40;
  input [7:0] p_20_41;
  input [7:0] p_20_42;
  input [7:0] p_20_43;
  input [7:0] p_20_44;
  input [7:0] p_20_45;
  input [7:0] p_20_46;
  input [7:0] p_20_47;
  input [7:0] p_20_48;
  input [7:0] p_20_49;
  input [7:0] p_20_50;
  input [7:0] p_20_51;
  input [7:0] p_20_52;
  input [7:0] p_20_53;
  input [7:0] p_20_54;
  input [7:0] p_20_55;
  input [7:0] p_20_56;
  input [7:0] p_20_57;
  input [7:0] p_20_58;
  input [7:0] p_20_59;
  input [7:0] p_20_60;
  input [7:0] p_20_61;
  input [7:0] p_20_62;
  input [7:0] p_20_63;
  input [7:0] p_20_64;
  input [7:0] p_20_65;
  input [7:0] p_21_0;
  input [7:0] p_21_1;
  input [7:0] p_21_2;
  input [7:0] p_21_3;
  input [7:0] p_21_4;
  input [7:0] p_21_5;
  input [7:0] p_21_6;
  input [7:0] p_21_7;
  input [7:0] p_21_8;
  input [7:0] p_21_9;
  input [7:0] p_21_10;
  input [7:0] p_21_11;
  input [7:0] p_21_12;
  input [7:0] p_21_13;
  input [7:0] p_21_14;
  input [7:0] p_21_15;
  input [7:0] p_21_16;
  input [7:0] p_21_17;
  input [7:0] p_21_18;
  input [7:0] p_21_19;
  input [7:0] p_21_20;
  input [7:0] p_21_21;
  input [7:0] p_21_22;
  input [7:0] p_21_23;
  input [7:0] p_21_24;
  input [7:0] p_21_25;
  input [7:0] p_21_26;
  input [7:0] p_21_27;
  input [7:0] p_21_28;
  input [7:0] p_21_29;
  input [7:0] p_21_30;
  input [7:0] p_21_31;
  input [7:0] p_21_32;
  input [7:0] p_21_33;
  input [7:0] p_21_34;
  input [7:0] p_21_35;
  input [7:0] p_21_36;
  input [7:0] p_21_37;
  input [7:0] p_21_38;
  input [7:0] p_21_39;
  input [7:0] p_21_40;
  input [7:0] p_21_41;
  input [7:0] p_21_42;
  input [7:0] p_21_43;
  input [7:0] p_21_44;
  input [7:0] p_21_45;
  input [7:0] p_21_46;
  input [7:0] p_21_47;
  input [7:0] p_21_48;
  input [7:0] p_21_49;
  input [7:0] p_21_50;
  input [7:0] p_21_51;
  input [7:0] p_21_52;
  input [7:0] p_21_53;
  input [7:0] p_21_54;
  input [7:0] p_21_55;
  input [7:0] p_21_56;
  input [7:0] p_21_57;
  input [7:0] p_21_58;
  input [7:0] p_21_59;
  input [7:0] p_21_60;
  input [7:0] p_21_61;
  input [7:0] p_21_62;
  input [7:0] p_21_63;
  input [7:0] p_21_64;
  input [7:0] p_21_65;
  input [7:0] p_22_0;
  input [7:0] p_22_1;
  input [7:0] p_22_2;
  input [7:0] p_22_3;
  input [7:0] p_22_4;
  input [7:0] p_22_5;
  input [7:0] p_22_6;
  input [7:0] p_22_7;
  input [7:0] p_22_8;
  input [7:0] p_22_9;
  input [7:0] p_22_10;
  input [7:0] p_22_11;
  input [7:0] p_22_12;
  input [7:0] p_22_13;
  input [7:0] p_22_14;
  input [7:0] p_22_15;
  input [7:0] p_22_16;
  input [7:0] p_22_17;
  input [7:0] p_22_18;
  input [7:0] p_22_19;
  input [7:0] p_22_20;
  input [7:0] p_22_21;
  input [7:0] p_22_22;
  input [7:0] p_22_23;
  input [7:0] p_22_24;
  input [7:0] p_22_25;
  input [7:0] p_22_26;
  input [7:0] p_22_27;
  input [7:0] p_22_28;
  input [7:0] p_22_29;
  input [7:0] p_22_30;
  input [7:0] p_22_31;
  input [7:0] p_22_32;
  input [7:0] p_22_33;
  input [7:0] p_22_34;
  input [7:0] p_22_35;
  input [7:0] p_22_36;
  input [7:0] p_22_37;
  input [7:0] p_22_38;
  input [7:0] p_22_39;
  input [7:0] p_22_40;
  input [7:0] p_22_41;
  input [7:0] p_22_42;
  input [7:0] p_22_43;
  input [7:0] p_22_44;
  input [7:0] p_22_45;
  input [7:0] p_22_46;
  input [7:0] p_22_47;
  input [7:0] p_22_48;
  input [7:0] p_22_49;
  input [7:0] p_22_50;
  input [7:0] p_22_51;
  input [7:0] p_22_52;
  input [7:0] p_22_53;
  input [7:0] p_22_54;
  input [7:0] p_22_55;
  input [7:0] p_22_56;
  input [7:0] p_22_57;
  input [7:0] p_22_58;
  input [7:0] p_22_59;
  input [7:0] p_22_60;
  input [7:0] p_22_61;
  input [7:0] p_22_62;
  input [7:0] p_22_63;
  input [7:0] p_22_64;
  input [7:0] p_22_65;
  input [7:0] p_23_0;
  input [7:0] p_23_1;
  input [7:0] p_23_2;
  input [7:0] p_23_3;
  input [7:0] p_23_4;
  input [7:0] p_23_5;
  input [7:0] p_23_6;
  input [7:0] p_23_7;
  input [7:0] p_23_8;
  input [7:0] p_23_9;
  input [7:0] p_23_10;
  input [7:0] p_23_11;
  input [7:0] p_23_12;
  input [7:0] p_23_13;
  input [7:0] p_23_14;
  input [7:0] p_23_15;
  input [7:0] p_23_16;
  input [7:0] p_23_17;
  input [7:0] p_23_18;
  input [7:0] p_23_19;
  input [7:0] p_23_20;
  input [7:0] p_23_21;
  input [7:0] p_23_22;
  input [7:0] p_23_23;
  input [7:0] p_23_24;
  input [7:0] p_23_25;
  input [7:0] p_23_26;
  input [7:0] p_23_27;
  input [7:0] p_23_28;
  input [7:0] p_23_29;
  input [7:0] p_23_30;
  input [7:0] p_23_31;
  input [7:0] p_23_32;
  input [7:0] p_23_33;
  input [7:0] p_23_34;
  input [7:0] p_23_35;
  input [7:0] p_23_36;
  input [7:0] p_23_37;
  input [7:0] p_23_38;
  input [7:0] p_23_39;
  input [7:0] p_23_40;
  input [7:0] p_23_41;
  input [7:0] p_23_42;
  input [7:0] p_23_43;
  input [7:0] p_23_44;
  input [7:0] p_23_45;
  input [7:0] p_23_46;
  input [7:0] p_23_47;
  input [7:0] p_23_48;
  input [7:0] p_23_49;
  input [7:0] p_23_50;
  input [7:0] p_23_51;
  input [7:0] p_23_52;
  input [7:0] p_23_53;
  input [7:0] p_23_54;
  input [7:0] p_23_55;
  input [7:0] p_23_56;
  input [7:0] p_23_57;
  input [7:0] p_23_58;
  input [7:0] p_23_59;
  input [7:0] p_23_60;
  input [7:0] p_23_61;
  input [7:0] p_23_62;
  input [7:0] p_23_63;
  input [7:0] p_23_64;
  input [7:0] p_23_65;
  input [7:0] p_24_0;
  input [7:0] p_24_1;
  input [7:0] p_24_2;
  input [7:0] p_24_3;
  input [7:0] p_24_4;
  input [7:0] p_24_5;
  input [7:0] p_24_6;
  input [7:0] p_24_7;
  input [7:0] p_24_8;
  input [7:0] p_24_9;
  input [7:0] p_24_10;
  input [7:0] p_24_11;
  input [7:0] p_24_12;
  input [7:0] p_24_13;
  input [7:0] p_24_14;
  input [7:0] p_24_15;
  input [7:0] p_24_16;
  input [7:0] p_24_17;
  input [7:0] p_24_18;
  input [7:0] p_24_19;
  input [7:0] p_24_20;
  input [7:0] p_24_21;
  input [7:0] p_24_22;
  input [7:0] p_24_23;
  input [7:0] p_24_24;
  input [7:0] p_24_25;
  input [7:0] p_24_26;
  input [7:0] p_24_27;
  input [7:0] p_24_28;
  input [7:0] p_24_29;
  input [7:0] p_24_30;
  input [7:0] p_24_31;
  input [7:0] p_24_32;
  input [7:0] p_24_33;
  input [7:0] p_24_34;
  input [7:0] p_24_35;
  input [7:0] p_24_36;
  input [7:0] p_24_37;
  input [7:0] p_24_38;
  input [7:0] p_24_39;
  input [7:0] p_24_40;
  input [7:0] p_24_41;
  input [7:0] p_24_42;
  input [7:0] p_24_43;
  input [7:0] p_24_44;
  input [7:0] p_24_45;
  input [7:0] p_24_46;
  input [7:0] p_24_47;
  input [7:0] p_24_48;
  input [7:0] p_24_49;
  input [7:0] p_24_50;
  input [7:0] p_24_51;
  input [7:0] p_24_52;
  input [7:0] p_24_53;
  input [7:0] p_24_54;
  input [7:0] p_24_55;
  input [7:0] p_24_56;
  input [7:0] p_24_57;
  input [7:0] p_24_58;
  input [7:0] p_24_59;
  input [7:0] p_24_60;
  input [7:0] p_24_61;
  input [7:0] p_24_62;
  input [7:0] p_24_63;
  input [7:0] p_24_64;
  input [7:0] p_24_65;
  input [7:0] p_25_0;
  input [7:0] p_25_1;
  input [7:0] p_25_2;
  input [7:0] p_25_3;
  input [7:0] p_25_4;
  input [7:0] p_25_5;
  input [7:0] p_25_6;
  input [7:0] p_25_7;
  input [7:0] p_25_8;
  input [7:0] p_25_9;
  input [7:0] p_25_10;
  input [7:0] p_25_11;
  input [7:0] p_25_12;
  input [7:0] p_25_13;
  input [7:0] p_25_14;
  input [7:0] p_25_15;
  input [7:0] p_25_16;
  input [7:0] p_25_17;
  input [7:0] p_25_18;
  input [7:0] p_25_19;
  input [7:0] p_25_20;
  input [7:0] p_25_21;
  input [7:0] p_25_22;
  input [7:0] p_25_23;
  input [7:0] p_25_24;
  input [7:0] p_25_25;
  input [7:0] p_25_26;
  input [7:0] p_25_27;
  input [7:0] p_25_28;
  input [7:0] p_25_29;
  input [7:0] p_25_30;
  input [7:0] p_25_31;
  input [7:0] p_25_32;
  input [7:0] p_25_33;
  input [7:0] p_25_34;
  input [7:0] p_25_35;
  input [7:0] p_25_36;
  input [7:0] p_25_37;
  input [7:0] p_25_38;
  input [7:0] p_25_39;
  input [7:0] p_25_40;
  input [7:0] p_25_41;
  input [7:0] p_25_42;
  input [7:0] p_25_43;
  input [7:0] p_25_44;
  input [7:0] p_25_45;
  input [7:0] p_25_46;
  input [7:0] p_25_47;
  input [7:0] p_25_48;
  input [7:0] p_25_49;
  input [7:0] p_25_50;
  input [7:0] p_25_51;
  input [7:0] p_25_52;
  input [7:0] p_25_53;
  input [7:0] p_25_54;
  input [7:0] p_25_55;
  input [7:0] p_25_56;
  input [7:0] p_25_57;
  input [7:0] p_25_58;
  input [7:0] p_25_59;
  input [7:0] p_25_60;
  input [7:0] p_25_61;
  input [7:0] p_25_62;
  input [7:0] p_25_63;
  input [7:0] p_25_64;
  input [7:0] p_25_65;
  input [7:0] p_26_0;
  input [7:0] p_26_1;
  input [7:0] p_26_2;
  input [7:0] p_26_3;
  input [7:0] p_26_4;
  input [7:0] p_26_5;
  input [7:0] p_26_6;
  input [7:0] p_26_7;
  input [7:0] p_26_8;
  input [7:0] p_26_9;
  input [7:0] p_26_10;
  input [7:0] p_26_11;
  input [7:0] p_26_12;
  input [7:0] p_26_13;
  input [7:0] p_26_14;
  input [7:0] p_26_15;
  input [7:0] p_26_16;
  input [7:0] p_26_17;
  input [7:0] p_26_18;
  input [7:0] p_26_19;
  input [7:0] p_26_20;
  input [7:0] p_26_21;
  input [7:0] p_26_22;
  input [7:0] p_26_23;
  input [7:0] p_26_24;
  input [7:0] p_26_25;
  input [7:0] p_26_26;
  input [7:0] p_26_27;
  input [7:0] p_26_28;
  input [7:0] p_26_29;
  input [7:0] p_26_30;
  input [7:0] p_26_31;
  input [7:0] p_26_32;
  input [7:0] p_26_33;
  input [7:0] p_26_34;
  input [7:0] p_26_35;
  input [7:0] p_26_36;
  input [7:0] p_26_37;
  input [7:0] p_26_38;
  input [7:0] p_26_39;
  input [7:0] p_26_40;
  input [7:0] p_26_41;
  input [7:0] p_26_42;
  input [7:0] p_26_43;
  input [7:0] p_26_44;
  input [7:0] p_26_45;
  input [7:0] p_26_46;
  input [7:0] p_26_47;
  input [7:0] p_26_48;
  input [7:0] p_26_49;
  input [7:0] p_26_50;
  input [7:0] p_26_51;
  input [7:0] p_26_52;
  input [7:0] p_26_53;
  input [7:0] p_26_54;
  input [7:0] p_26_55;
  input [7:0] p_26_56;
  input [7:0] p_26_57;
  input [7:0] p_26_58;
  input [7:0] p_26_59;
  input [7:0] p_26_60;
  input [7:0] p_26_61;
  input [7:0] p_26_62;
  input [7:0] p_26_63;
  input [7:0] p_26_64;
  input [7:0] p_26_65;
  input [7:0] p_27_0;
  input [7:0] p_27_1;
  input [7:0] p_27_2;
  input [7:0] p_27_3;
  input [7:0] p_27_4;
  input [7:0] p_27_5;
  input [7:0] p_27_6;
  input [7:0] p_27_7;
  input [7:0] p_27_8;
  input [7:0] p_27_9;
  input [7:0] p_27_10;
  input [7:0] p_27_11;
  input [7:0] p_27_12;
  input [7:0] p_27_13;
  input [7:0] p_27_14;
  input [7:0] p_27_15;
  input [7:0] p_27_16;
  input [7:0] p_27_17;
  input [7:0] p_27_18;
  input [7:0] p_27_19;
  input [7:0] p_27_20;
  input [7:0] p_27_21;
  input [7:0] p_27_22;
  input [7:0] p_27_23;
  input [7:0] p_27_24;
  input [7:0] p_27_25;
  input [7:0] p_27_26;
  input [7:0] p_27_27;
  input [7:0] p_27_28;
  input [7:0] p_27_29;
  input [7:0] p_27_30;
  input [7:0] p_27_31;
  input [7:0] p_27_32;
  input [7:0] p_27_33;
  input [7:0] p_27_34;
  input [7:0] p_27_35;
  input [7:0] p_27_36;
  input [7:0] p_27_37;
  input [7:0] p_27_38;
  input [7:0] p_27_39;
  input [7:0] p_27_40;
  input [7:0] p_27_41;
  input [7:0] p_27_42;
  input [7:0] p_27_43;
  input [7:0] p_27_44;
  input [7:0] p_27_45;
  input [7:0] p_27_46;
  input [7:0] p_27_47;
  input [7:0] p_27_48;
  input [7:0] p_27_49;
  input [7:0] p_27_50;
  input [7:0] p_27_51;
  input [7:0] p_27_52;
  input [7:0] p_27_53;
  input [7:0] p_27_54;
  input [7:0] p_27_55;
  input [7:0] p_27_56;
  input [7:0] p_27_57;
  input [7:0] p_27_58;
  input [7:0] p_27_59;
  input [7:0] p_27_60;
  input [7:0] p_27_61;
  input [7:0] p_27_62;
  input [7:0] p_27_63;
  input [7:0] p_27_64;
  input [7:0] p_27_65;
  input [7:0] p_28_0;
  input [7:0] p_28_1;
  input [7:0] p_28_2;
  input [7:0] p_28_3;
  input [7:0] p_28_4;
  input [7:0] p_28_5;
  input [7:0] p_28_6;
  input [7:0] p_28_7;
  input [7:0] p_28_8;
  input [7:0] p_28_9;
  input [7:0] p_28_10;
  input [7:0] p_28_11;
  input [7:0] p_28_12;
  input [7:0] p_28_13;
  input [7:0] p_28_14;
  input [7:0] p_28_15;
  input [7:0] p_28_16;
  input [7:0] p_28_17;
  input [7:0] p_28_18;
  input [7:0] p_28_19;
  input [7:0] p_28_20;
  input [7:0] p_28_21;
  input [7:0] p_28_22;
  input [7:0] p_28_23;
  input [7:0] p_28_24;
  input [7:0] p_28_25;
  input [7:0] p_28_26;
  input [7:0] p_28_27;
  input [7:0] p_28_28;
  input [7:0] p_28_29;
  input [7:0] p_28_30;
  input [7:0] p_28_31;
  input [7:0] p_28_32;
  input [7:0] p_28_33;
  input [7:0] p_28_34;
  input [7:0] p_28_35;
  input [7:0] p_28_36;
  input [7:0] p_28_37;
  input [7:0] p_28_38;
  input [7:0] p_28_39;
  input [7:0] p_28_40;
  input [7:0] p_28_41;
  input [7:0] p_28_42;
  input [7:0] p_28_43;
  input [7:0] p_28_44;
  input [7:0] p_28_45;
  input [7:0] p_28_46;
  input [7:0] p_28_47;
  input [7:0] p_28_48;
  input [7:0] p_28_49;
  input [7:0] p_28_50;
  input [7:0] p_28_51;
  input [7:0] p_28_52;
  input [7:0] p_28_53;
  input [7:0] p_28_54;
  input [7:0] p_28_55;
  input [7:0] p_28_56;
  input [7:0] p_28_57;
  input [7:0] p_28_58;
  input [7:0] p_28_59;
  input [7:0] p_28_60;
  input [7:0] p_28_61;
  input [7:0] p_28_62;
  input [7:0] p_28_63;
  input [7:0] p_28_64;
  input [7:0] p_28_65;
  input [7:0] p_29_0;
  input [7:0] p_29_1;
  input [7:0] p_29_2;
  input [7:0] p_29_3;
  input [7:0] p_29_4;
  input [7:0] p_29_5;
  input [7:0] p_29_6;
  input [7:0] p_29_7;
  input [7:0] p_29_8;
  input [7:0] p_29_9;
  input [7:0] p_29_10;
  input [7:0] p_29_11;
  input [7:0] p_29_12;
  input [7:0] p_29_13;
  input [7:0] p_29_14;
  input [7:0] p_29_15;
  input [7:0] p_29_16;
  input [7:0] p_29_17;
  input [7:0] p_29_18;
  input [7:0] p_29_19;
  input [7:0] p_29_20;
  input [7:0] p_29_21;
  input [7:0] p_29_22;
  input [7:0] p_29_23;
  input [7:0] p_29_24;
  input [7:0] p_29_25;
  input [7:0] p_29_26;
  input [7:0] p_29_27;
  input [7:0] p_29_28;
  input [7:0] p_29_29;
  input [7:0] p_29_30;
  input [7:0] p_29_31;
  input [7:0] p_29_32;
  input [7:0] p_29_33;
  input [7:0] p_29_34;
  input [7:0] p_29_35;
  input [7:0] p_29_36;
  input [7:0] p_29_37;
  input [7:0] p_29_38;
  input [7:0] p_29_39;
  input [7:0] p_29_40;
  input [7:0] p_29_41;
  input [7:0] p_29_42;
  input [7:0] p_29_43;
  input [7:0] p_29_44;
  input [7:0] p_29_45;
  input [7:0] p_29_46;
  input [7:0] p_29_47;
  input [7:0] p_29_48;
  input [7:0] p_29_49;
  input [7:0] p_29_50;
  input [7:0] p_29_51;
  input [7:0] p_29_52;
  input [7:0] p_29_53;
  input [7:0] p_29_54;
  input [7:0] p_29_55;
  input [7:0] p_29_56;
  input [7:0] p_29_57;
  input [7:0] p_29_58;
  input [7:0] p_29_59;
  input [7:0] p_29_60;
  input [7:0] p_29_61;
  input [7:0] p_29_62;
  input [7:0] p_29_63;
  input [7:0] p_29_64;
  input [7:0] p_29_65;
  input [7:0] p_30_0;
  input [7:0] p_30_1;
  input [7:0] p_30_2;
  input [7:0] p_30_3;
  input [7:0] p_30_4;
  input [7:0] p_30_5;
  input [7:0] p_30_6;
  input [7:0] p_30_7;
  input [7:0] p_30_8;
  input [7:0] p_30_9;
  input [7:0] p_30_10;
  input [7:0] p_30_11;
  input [7:0] p_30_12;
  input [7:0] p_30_13;
  input [7:0] p_30_14;
  input [7:0] p_30_15;
  input [7:0] p_30_16;
  input [7:0] p_30_17;
  input [7:0] p_30_18;
  input [7:0] p_30_19;
  input [7:0] p_30_20;
  input [7:0] p_30_21;
  input [7:0] p_30_22;
  input [7:0] p_30_23;
  input [7:0] p_30_24;
  input [7:0] p_30_25;
  input [7:0] p_30_26;
  input [7:0] p_30_27;
  input [7:0] p_30_28;
  input [7:0] p_30_29;
  input [7:0] p_30_30;
  input [7:0] p_30_31;
  input [7:0] p_30_32;
  input [7:0] p_30_33;
  input [7:0] p_30_34;
  input [7:0] p_30_35;
  input [7:0] p_30_36;
  input [7:0] p_30_37;
  input [7:0] p_30_38;
  input [7:0] p_30_39;
  input [7:0] p_30_40;
  input [7:0] p_30_41;
  input [7:0] p_30_42;
  input [7:0] p_30_43;
  input [7:0] p_30_44;
  input [7:0] p_30_45;
  input [7:0] p_30_46;
  input [7:0] p_30_47;
  input [7:0] p_30_48;
  input [7:0] p_30_49;
  input [7:0] p_30_50;
  input [7:0] p_30_51;
  input [7:0] p_30_52;
  input [7:0] p_30_53;
  input [7:0] p_30_54;
  input [7:0] p_30_55;
  input [7:0] p_30_56;
  input [7:0] p_30_57;
  input [7:0] p_30_58;
  input [7:0] p_30_59;
  input [7:0] p_30_60;
  input [7:0] p_30_61;
  input [7:0] p_30_62;
  input [7:0] p_30_63;
  input [7:0] p_30_64;
  input [7:0] p_30_65;
  input [7:0] p_31_0;
  input [7:0] p_31_1;
  input [7:0] p_31_2;
  input [7:0] p_31_3;
  input [7:0] p_31_4;
  input [7:0] p_31_5;
  input [7:0] p_31_6;
  input [7:0] p_31_7;
  input [7:0] p_31_8;
  input [7:0] p_31_9;
  input [7:0] p_31_10;
  input [7:0] p_31_11;
  input [7:0] p_31_12;
  input [7:0] p_31_13;
  input [7:0] p_31_14;
  input [7:0] p_31_15;
  input [7:0] p_31_16;
  input [7:0] p_31_17;
  input [7:0] p_31_18;
  input [7:0] p_31_19;
  input [7:0] p_31_20;
  input [7:0] p_31_21;
  input [7:0] p_31_22;
  input [7:0] p_31_23;
  input [7:0] p_31_24;
  input [7:0] p_31_25;
  input [7:0] p_31_26;
  input [7:0] p_31_27;
  input [7:0] p_31_28;
  input [7:0] p_31_29;
  input [7:0] p_31_30;
  input [7:0] p_31_31;
  input [7:0] p_31_32;
  input [7:0] p_31_33;
  input [7:0] p_31_34;
  input [7:0] p_31_35;
  input [7:0] p_31_36;
  input [7:0] p_31_37;
  input [7:0] p_31_38;
  input [7:0] p_31_39;
  input [7:0] p_31_40;
  input [7:0] p_31_41;
  input [7:0] p_31_42;
  input [7:0] p_31_43;
  input [7:0] p_31_44;
  input [7:0] p_31_45;
  input [7:0] p_31_46;
  input [7:0] p_31_47;
  input [7:0] p_31_48;
  input [7:0] p_31_49;
  input [7:0] p_31_50;
  input [7:0] p_31_51;
  input [7:0] p_31_52;
  input [7:0] p_31_53;
  input [7:0] p_31_54;
  input [7:0] p_31_55;
  input [7:0] p_31_56;
  input [7:0] p_31_57;
  input [7:0] p_31_58;
  input [7:0] p_31_59;
  input [7:0] p_31_60;
  input [7:0] p_31_61;
  input [7:0] p_31_62;
  input [7:0] p_31_63;
  input [7:0] p_31_64;
  input [7:0] p_31_65;
  input [7:0] p_32_0;
  input [7:0] p_32_1;
  input [7:0] p_32_2;
  input [7:0] p_32_3;
  input [7:0] p_32_4;
  input [7:0] p_32_5;
  input [7:0] p_32_6;
  input [7:0] p_32_7;
  input [7:0] p_32_8;
  input [7:0] p_32_9;
  input [7:0] p_32_10;
  input [7:0] p_32_11;
  input [7:0] p_32_12;
  input [7:0] p_32_13;
  input [7:0] p_32_14;
  input [7:0] p_32_15;
  input [7:0] p_32_16;
  input [7:0] p_32_17;
  input [7:0] p_32_18;
  input [7:0] p_32_19;
  input [7:0] p_32_20;
  input [7:0] p_32_21;
  input [7:0] p_32_22;
  input [7:0] p_32_23;
  input [7:0] p_32_24;
  input [7:0] p_32_25;
  input [7:0] p_32_26;
  input [7:0] p_32_27;
  input [7:0] p_32_28;
  input [7:0] p_32_29;
  input [7:0] p_32_30;
  input [7:0] p_32_31;
  input [7:0] p_32_32;
  input [7:0] p_32_33;
  input [7:0] p_32_34;
  input [7:0] p_32_35;
  input [7:0] p_32_36;
  input [7:0] p_32_37;
  input [7:0] p_32_38;
  input [7:0] p_32_39;
  input [7:0] p_32_40;
  input [7:0] p_32_41;
  input [7:0] p_32_42;
  input [7:0] p_32_43;
  input [7:0] p_32_44;
  input [7:0] p_32_45;
  input [7:0] p_32_46;
  input [7:0] p_32_47;
  input [7:0] p_32_48;
  input [7:0] p_32_49;
  input [7:0] p_32_50;
  input [7:0] p_32_51;
  input [7:0] p_32_52;
  input [7:0] p_32_53;
  input [7:0] p_32_54;
  input [7:0] p_32_55;
  input [7:0] p_32_56;
  input [7:0] p_32_57;
  input [7:0] p_32_58;
  input [7:0] p_32_59;
  input [7:0] p_32_60;
  input [7:0] p_32_61;
  input [7:0] p_32_62;
  input [7:0] p_32_63;
  input [7:0] p_32_64;
  input [7:0] p_32_65;
  input [7:0] p_33_0;
  input [7:0] p_33_1;
  input [7:0] p_33_2;
  input [7:0] p_33_3;
  input [7:0] p_33_4;
  input [7:0] p_33_5;
  input [7:0] p_33_6;
  input [7:0] p_33_7;
  input [7:0] p_33_8;
  input [7:0] p_33_9;
  input [7:0] p_33_10;
  input [7:0] p_33_11;
  input [7:0] p_33_12;
  input [7:0] p_33_13;
  input [7:0] p_33_14;
  input [7:0] p_33_15;
  input [7:0] p_33_16;
  input [7:0] p_33_17;
  input [7:0] p_33_18;
  input [7:0] p_33_19;
  input [7:0] p_33_20;
  input [7:0] p_33_21;
  input [7:0] p_33_22;
  input [7:0] p_33_23;
  input [7:0] p_33_24;
  input [7:0] p_33_25;
  input [7:0] p_33_26;
  input [7:0] p_33_27;
  input [7:0] p_33_28;
  input [7:0] p_33_29;
  input [7:0] p_33_30;
  input [7:0] p_33_31;
  input [7:0] p_33_32;
  input [7:0] p_33_33;
  input [7:0] p_33_34;
  input [7:0] p_33_35;
  input [7:0] p_33_36;
  input [7:0] p_33_37;
  input [7:0] p_33_38;
  input [7:0] p_33_39;
  input [7:0] p_33_40;
  input [7:0] p_33_41;
  input [7:0] p_33_42;
  input [7:0] p_33_43;
  input [7:0] p_33_44;
  input [7:0] p_33_45;
  input [7:0] p_33_46;
  input [7:0] p_33_47;
  input [7:0] p_33_48;
  input [7:0] p_33_49;
  input [7:0] p_33_50;
  input [7:0] p_33_51;
  input [7:0] p_33_52;
  input [7:0] p_33_53;
  input [7:0] p_33_54;
  input [7:0] p_33_55;
  input [7:0] p_33_56;
  input [7:0] p_33_57;
  input [7:0] p_33_58;
  input [7:0] p_33_59;
  input [7:0] p_33_60;
  input [7:0] p_33_61;
  input [7:0] p_33_62;
  input [7:0] p_33_63;
  input [7:0] p_33_64;
  input [7:0] p_33_65;
  input [7:0] p_34_0;
  input [7:0] p_34_1;
  input [7:0] p_34_2;
  input [7:0] p_34_3;
  input [7:0] p_34_4;
  input [7:0] p_34_5;
  input [7:0] p_34_6;
  input [7:0] p_34_7;
  input [7:0] p_34_8;
  input [7:0] p_34_9;
  input [7:0] p_34_10;
  input [7:0] p_34_11;
  input [7:0] p_34_12;
  input [7:0] p_34_13;
  input [7:0] p_34_14;
  input [7:0] p_34_15;
  input [7:0] p_34_16;
  input [7:0] p_34_17;
  input [7:0] p_34_18;
  input [7:0] p_34_19;
  input [7:0] p_34_20;
  input [7:0] p_34_21;
  input [7:0] p_34_22;
  input [7:0] p_34_23;
  input [7:0] p_34_24;
  input [7:0] p_34_25;
  input [7:0] p_34_26;
  input [7:0] p_34_27;
  input [7:0] p_34_28;
  input [7:0] p_34_29;
  input [7:0] p_34_30;
  input [7:0] p_34_31;
  input [7:0] p_34_32;
  input [7:0] p_34_33;
  input [7:0] p_34_34;
  input [7:0] p_34_35;
  input [7:0] p_34_36;
  input [7:0] p_34_37;
  input [7:0] p_34_38;
  input [7:0] p_34_39;
  input [7:0] p_34_40;
  input [7:0] p_34_41;
  input [7:0] p_34_42;
  input [7:0] p_34_43;
  input [7:0] p_34_44;
  input [7:0] p_34_45;
  input [7:0] p_34_46;
  input [7:0] p_34_47;
  input [7:0] p_34_48;
  input [7:0] p_34_49;
  input [7:0] p_34_50;
  input [7:0] p_34_51;
  input [7:0] p_34_52;
  input [7:0] p_34_53;
  input [7:0] p_34_54;
  input [7:0] p_34_55;
  input [7:0] p_34_56;
  input [7:0] p_34_57;
  input [7:0] p_34_58;
  input [7:0] p_34_59;
  input [7:0] p_34_60;
  input [7:0] p_34_61;
  input [7:0] p_34_62;
  input [7:0] p_34_63;
  input [7:0] p_34_64;
  input [7:0] p_34_65;
  input [7:0] p_35_0;
  input [7:0] p_35_1;
  input [7:0] p_35_2;
  input [7:0] p_35_3;
  input [7:0] p_35_4;
  input [7:0] p_35_5;
  input [7:0] p_35_6;
  input [7:0] p_35_7;
  input [7:0] p_35_8;
  input [7:0] p_35_9;
  input [7:0] p_35_10;
  input [7:0] p_35_11;
  input [7:0] p_35_12;
  input [7:0] p_35_13;
  input [7:0] p_35_14;
  input [7:0] p_35_15;
  input [7:0] p_35_16;
  input [7:0] p_35_17;
  input [7:0] p_35_18;
  input [7:0] p_35_19;
  input [7:0] p_35_20;
  input [7:0] p_35_21;
  input [7:0] p_35_22;
  input [7:0] p_35_23;
  input [7:0] p_35_24;
  input [7:0] p_35_25;
  input [7:0] p_35_26;
  input [7:0] p_35_27;
  input [7:0] p_35_28;
  input [7:0] p_35_29;
  input [7:0] p_35_30;
  input [7:0] p_35_31;
  input [7:0] p_35_32;
  input [7:0] p_35_33;
  input [7:0] p_35_34;
  input [7:0] p_35_35;
  input [7:0] p_35_36;
  input [7:0] p_35_37;
  input [7:0] p_35_38;
  input [7:0] p_35_39;
  input [7:0] p_35_40;
  input [7:0] p_35_41;
  input [7:0] p_35_42;
  input [7:0] p_35_43;
  input [7:0] p_35_44;
  input [7:0] p_35_45;
  input [7:0] p_35_46;
  input [7:0] p_35_47;
  input [7:0] p_35_48;
  input [7:0] p_35_49;
  input [7:0] p_35_50;
  input [7:0] p_35_51;
  input [7:0] p_35_52;
  input [7:0] p_35_53;
  input [7:0] p_35_54;
  input [7:0] p_35_55;
  input [7:0] p_35_56;
  input [7:0] p_35_57;
  input [7:0] p_35_58;
  input [7:0] p_35_59;
  input [7:0] p_35_60;
  input [7:0] p_35_61;
  input [7:0] p_35_62;
  input [7:0] p_35_63;
  input [7:0] p_35_64;
  input [7:0] p_35_65;
  input [7:0] p_36_0;
  input [7:0] p_36_1;
  input [7:0] p_36_2;
  input [7:0] p_36_3;
  input [7:0] p_36_4;
  input [7:0] p_36_5;
  input [7:0] p_36_6;
  input [7:0] p_36_7;
  input [7:0] p_36_8;
  input [7:0] p_36_9;
  input [7:0] p_36_10;
  input [7:0] p_36_11;
  input [7:0] p_36_12;
  input [7:0] p_36_13;
  input [7:0] p_36_14;
  input [7:0] p_36_15;
  input [7:0] p_36_16;
  input [7:0] p_36_17;
  input [7:0] p_36_18;
  input [7:0] p_36_19;
  input [7:0] p_36_20;
  input [7:0] p_36_21;
  input [7:0] p_36_22;
  input [7:0] p_36_23;
  input [7:0] p_36_24;
  input [7:0] p_36_25;
  input [7:0] p_36_26;
  input [7:0] p_36_27;
  input [7:0] p_36_28;
  input [7:0] p_36_29;
  input [7:0] p_36_30;
  input [7:0] p_36_31;
  input [7:0] p_36_32;
  input [7:0] p_36_33;
  input [7:0] p_36_34;
  input [7:0] p_36_35;
  input [7:0] p_36_36;
  input [7:0] p_36_37;
  input [7:0] p_36_38;
  input [7:0] p_36_39;
  input [7:0] p_36_40;
  input [7:0] p_36_41;
  input [7:0] p_36_42;
  input [7:0] p_36_43;
  input [7:0] p_36_44;
  input [7:0] p_36_45;
  input [7:0] p_36_46;
  input [7:0] p_36_47;
  input [7:0] p_36_48;
  input [7:0] p_36_49;
  input [7:0] p_36_50;
  input [7:0] p_36_51;
  input [7:0] p_36_52;
  input [7:0] p_36_53;
  input [7:0] p_36_54;
  input [7:0] p_36_55;
  input [7:0] p_36_56;
  input [7:0] p_36_57;
  input [7:0] p_36_58;
  input [7:0] p_36_59;
  input [7:0] p_36_60;
  input [7:0] p_36_61;
  input [7:0] p_36_62;
  input [7:0] p_36_63;
  input [7:0] p_36_64;
  input [7:0] p_36_65;
  input [7:0] p_37_0;
  input [7:0] p_37_1;
  input [7:0] p_37_2;
  input [7:0] p_37_3;
  input [7:0] p_37_4;
  input [7:0] p_37_5;
  input [7:0] p_37_6;
  input [7:0] p_37_7;
  input [7:0] p_37_8;
  input [7:0] p_37_9;
  input [7:0] p_37_10;
  input [7:0] p_37_11;
  input [7:0] p_37_12;
  input [7:0] p_37_13;
  input [7:0] p_37_14;
  input [7:0] p_37_15;
  input [7:0] p_37_16;
  input [7:0] p_37_17;
  input [7:0] p_37_18;
  input [7:0] p_37_19;
  input [7:0] p_37_20;
  input [7:0] p_37_21;
  input [7:0] p_37_22;
  input [7:0] p_37_23;
  input [7:0] p_37_24;
  input [7:0] p_37_25;
  input [7:0] p_37_26;
  input [7:0] p_37_27;
  input [7:0] p_37_28;
  input [7:0] p_37_29;
  input [7:0] p_37_30;
  input [7:0] p_37_31;
  input [7:0] p_37_32;
  input [7:0] p_37_33;
  input [7:0] p_37_34;
  input [7:0] p_37_35;
  input [7:0] p_37_36;
  input [7:0] p_37_37;
  input [7:0] p_37_38;
  input [7:0] p_37_39;
  input [7:0] p_37_40;
  input [7:0] p_37_41;
  input [7:0] p_37_42;
  input [7:0] p_37_43;
  input [7:0] p_37_44;
  input [7:0] p_37_45;
  input [7:0] p_37_46;
  input [7:0] p_37_47;
  input [7:0] p_37_48;
  input [7:0] p_37_49;
  input [7:0] p_37_50;
  input [7:0] p_37_51;
  input [7:0] p_37_52;
  input [7:0] p_37_53;
  input [7:0] p_37_54;
  input [7:0] p_37_55;
  input [7:0] p_37_56;
  input [7:0] p_37_57;
  input [7:0] p_37_58;
  input [7:0] p_37_59;
  input [7:0] p_37_60;
  input [7:0] p_37_61;
  input [7:0] p_37_62;
  input [7:0] p_37_63;
  input [7:0] p_37_64;
  input [7:0] p_37_65;
  input [7:0] p_38_0;
  input [7:0] p_38_1;
  input [7:0] p_38_2;
  input [7:0] p_38_3;
  input [7:0] p_38_4;
  input [7:0] p_38_5;
  input [7:0] p_38_6;
  input [7:0] p_38_7;
  input [7:0] p_38_8;
  input [7:0] p_38_9;
  input [7:0] p_38_10;
  input [7:0] p_38_11;
  input [7:0] p_38_12;
  input [7:0] p_38_13;
  input [7:0] p_38_14;
  input [7:0] p_38_15;
  input [7:0] p_38_16;
  input [7:0] p_38_17;
  input [7:0] p_38_18;
  input [7:0] p_38_19;
  input [7:0] p_38_20;
  input [7:0] p_38_21;
  input [7:0] p_38_22;
  input [7:0] p_38_23;
  input [7:0] p_38_24;
  input [7:0] p_38_25;
  input [7:0] p_38_26;
  input [7:0] p_38_27;
  input [7:0] p_38_28;
  input [7:0] p_38_29;
  input [7:0] p_38_30;
  input [7:0] p_38_31;
  input [7:0] p_38_32;
  input [7:0] p_38_33;
  input [7:0] p_38_34;
  input [7:0] p_38_35;
  input [7:0] p_38_36;
  input [7:0] p_38_37;
  input [7:0] p_38_38;
  input [7:0] p_38_39;
  input [7:0] p_38_40;
  input [7:0] p_38_41;
  input [7:0] p_38_42;
  input [7:0] p_38_43;
  input [7:0] p_38_44;
  input [7:0] p_38_45;
  input [7:0] p_38_46;
  input [7:0] p_38_47;
  input [7:0] p_38_48;
  input [7:0] p_38_49;
  input [7:0] p_38_50;
  input [7:0] p_38_51;
  input [7:0] p_38_52;
  input [7:0] p_38_53;
  input [7:0] p_38_54;
  input [7:0] p_38_55;
  input [7:0] p_38_56;
  input [7:0] p_38_57;
  input [7:0] p_38_58;
  input [7:0] p_38_59;
  input [7:0] p_38_60;
  input [7:0] p_38_61;
  input [7:0] p_38_62;
  input [7:0] p_38_63;
  input [7:0] p_38_64;
  input [7:0] p_38_65;
  input [7:0] p_39_0;
  input [7:0] p_39_1;
  input [7:0] p_39_2;
  input [7:0] p_39_3;
  input [7:0] p_39_4;
  input [7:0] p_39_5;
  input [7:0] p_39_6;
  input [7:0] p_39_7;
  input [7:0] p_39_8;
  input [7:0] p_39_9;
  input [7:0] p_39_10;
  input [7:0] p_39_11;
  input [7:0] p_39_12;
  input [7:0] p_39_13;
  input [7:0] p_39_14;
  input [7:0] p_39_15;
  input [7:0] p_39_16;
  input [7:0] p_39_17;
  input [7:0] p_39_18;
  input [7:0] p_39_19;
  input [7:0] p_39_20;
  input [7:0] p_39_21;
  input [7:0] p_39_22;
  input [7:0] p_39_23;
  input [7:0] p_39_24;
  input [7:0] p_39_25;
  input [7:0] p_39_26;
  input [7:0] p_39_27;
  input [7:0] p_39_28;
  input [7:0] p_39_29;
  input [7:0] p_39_30;
  input [7:0] p_39_31;
  input [7:0] p_39_32;
  input [7:0] p_39_33;
  input [7:0] p_39_34;
  input [7:0] p_39_35;
  input [7:0] p_39_36;
  input [7:0] p_39_37;
  input [7:0] p_39_38;
  input [7:0] p_39_39;
  input [7:0] p_39_40;
  input [7:0] p_39_41;
  input [7:0] p_39_42;
  input [7:0] p_39_43;
  input [7:0] p_39_44;
  input [7:0] p_39_45;
  input [7:0] p_39_46;
  input [7:0] p_39_47;
  input [7:0] p_39_48;
  input [7:0] p_39_49;
  input [7:0] p_39_50;
  input [7:0] p_39_51;
  input [7:0] p_39_52;
  input [7:0] p_39_53;
  input [7:0] p_39_54;
  input [7:0] p_39_55;
  input [7:0] p_39_56;
  input [7:0] p_39_57;
  input [7:0] p_39_58;
  input [7:0] p_39_59;
  input [7:0] p_39_60;
  input [7:0] p_39_61;
  input [7:0] p_39_62;
  input [7:0] p_39_63;
  input [7:0] p_39_64;
  input [7:0] p_39_65;
  input [7:0] p_40_0;
  input [7:0] p_40_1;
  input [7:0] p_40_2;
  input [7:0] p_40_3;
  input [7:0] p_40_4;
  input [7:0] p_40_5;
  input [7:0] p_40_6;
  input [7:0] p_40_7;
  input [7:0] p_40_8;
  input [7:0] p_40_9;
  input [7:0] p_40_10;
  input [7:0] p_40_11;
  input [7:0] p_40_12;
  input [7:0] p_40_13;
  input [7:0] p_40_14;
  input [7:0] p_40_15;
  input [7:0] p_40_16;
  input [7:0] p_40_17;
  input [7:0] p_40_18;
  input [7:0] p_40_19;
  input [7:0] p_40_20;
  input [7:0] p_40_21;
  input [7:0] p_40_22;
  input [7:0] p_40_23;
  input [7:0] p_40_24;
  input [7:0] p_40_25;
  input [7:0] p_40_26;
  input [7:0] p_40_27;
  input [7:0] p_40_28;
  input [7:0] p_40_29;
  input [7:0] p_40_30;
  input [7:0] p_40_31;
  input [7:0] p_40_32;
  input [7:0] p_40_33;
  input [7:0] p_40_34;
  input [7:0] p_40_35;
  input [7:0] p_40_36;
  input [7:0] p_40_37;
  input [7:0] p_40_38;
  input [7:0] p_40_39;
  input [7:0] p_40_40;
  input [7:0] p_40_41;
  input [7:0] p_40_42;
  input [7:0] p_40_43;
  input [7:0] p_40_44;
  input [7:0] p_40_45;
  input [7:0] p_40_46;
  input [7:0] p_40_47;
  input [7:0] p_40_48;
  input [7:0] p_40_49;
  input [7:0] p_40_50;
  input [7:0] p_40_51;
  input [7:0] p_40_52;
  input [7:0] p_40_53;
  input [7:0] p_40_54;
  input [7:0] p_40_55;
  input [7:0] p_40_56;
  input [7:0] p_40_57;
  input [7:0] p_40_58;
  input [7:0] p_40_59;
  input [7:0] p_40_60;
  input [7:0] p_40_61;
  input [7:0] p_40_62;
  input [7:0] p_40_63;
  input [7:0] p_40_64;
  input [7:0] p_40_65;
  input [7:0] p_41_0;
  input [7:0] p_41_1;
  input [7:0] p_41_2;
  input [7:0] p_41_3;
  input [7:0] p_41_4;
  input [7:0] p_41_5;
  input [7:0] p_41_6;
  input [7:0] p_41_7;
  input [7:0] p_41_8;
  input [7:0] p_41_9;
  input [7:0] p_41_10;
  input [7:0] p_41_11;
  input [7:0] p_41_12;
  input [7:0] p_41_13;
  input [7:0] p_41_14;
  input [7:0] p_41_15;
  input [7:0] p_41_16;
  input [7:0] p_41_17;
  input [7:0] p_41_18;
  input [7:0] p_41_19;
  input [7:0] p_41_20;
  input [7:0] p_41_21;
  input [7:0] p_41_22;
  input [7:0] p_41_23;
  input [7:0] p_41_24;
  input [7:0] p_41_25;
  input [7:0] p_41_26;
  input [7:0] p_41_27;
  input [7:0] p_41_28;
  input [7:0] p_41_29;
  input [7:0] p_41_30;
  input [7:0] p_41_31;
  input [7:0] p_41_32;
  input [7:0] p_41_33;
  input [7:0] p_41_34;
  input [7:0] p_41_35;
  input [7:0] p_41_36;
  input [7:0] p_41_37;
  input [7:0] p_41_38;
  input [7:0] p_41_39;
  input [7:0] p_41_40;
  input [7:0] p_41_41;
  input [7:0] p_41_42;
  input [7:0] p_41_43;
  input [7:0] p_41_44;
  input [7:0] p_41_45;
  input [7:0] p_41_46;
  input [7:0] p_41_47;
  input [7:0] p_41_48;
  input [7:0] p_41_49;
  input [7:0] p_41_50;
  input [7:0] p_41_51;
  input [7:0] p_41_52;
  input [7:0] p_41_53;
  input [7:0] p_41_54;
  input [7:0] p_41_55;
  input [7:0] p_41_56;
  input [7:0] p_41_57;
  input [7:0] p_41_58;
  input [7:0] p_41_59;
  input [7:0] p_41_60;
  input [7:0] p_41_61;
  input [7:0] p_41_62;
  input [7:0] p_41_63;
  input [7:0] p_41_64;
  input [7:0] p_41_65;
  input [7:0] p_42_0;
  input [7:0] p_42_1;
  input [7:0] p_42_2;
  input [7:0] p_42_3;
  input [7:0] p_42_4;
  input [7:0] p_42_5;
  input [7:0] p_42_6;
  input [7:0] p_42_7;
  input [7:0] p_42_8;
  input [7:0] p_42_9;
  input [7:0] p_42_10;
  input [7:0] p_42_11;
  input [7:0] p_42_12;
  input [7:0] p_42_13;
  input [7:0] p_42_14;
  input [7:0] p_42_15;
  input [7:0] p_42_16;
  input [7:0] p_42_17;
  input [7:0] p_42_18;
  input [7:0] p_42_19;
  input [7:0] p_42_20;
  input [7:0] p_42_21;
  input [7:0] p_42_22;
  input [7:0] p_42_23;
  input [7:0] p_42_24;
  input [7:0] p_42_25;
  input [7:0] p_42_26;
  input [7:0] p_42_27;
  input [7:0] p_42_28;
  input [7:0] p_42_29;
  input [7:0] p_42_30;
  input [7:0] p_42_31;
  input [7:0] p_42_32;
  input [7:0] p_42_33;
  input [7:0] p_42_34;
  input [7:0] p_42_35;
  input [7:0] p_42_36;
  input [7:0] p_42_37;
  input [7:0] p_42_38;
  input [7:0] p_42_39;
  input [7:0] p_42_40;
  input [7:0] p_42_41;
  input [7:0] p_42_42;
  input [7:0] p_42_43;
  input [7:0] p_42_44;
  input [7:0] p_42_45;
  input [7:0] p_42_46;
  input [7:0] p_42_47;
  input [7:0] p_42_48;
  input [7:0] p_42_49;
  input [7:0] p_42_50;
  input [7:0] p_42_51;
  input [7:0] p_42_52;
  input [7:0] p_42_53;
  input [7:0] p_42_54;
  input [7:0] p_42_55;
  input [7:0] p_42_56;
  input [7:0] p_42_57;
  input [7:0] p_42_58;
  input [7:0] p_42_59;
  input [7:0] p_42_60;
  input [7:0] p_42_61;
  input [7:0] p_42_62;
  input [7:0] p_42_63;
  input [7:0] p_42_64;
  input [7:0] p_42_65;
  input [7:0] p_43_0;
  input [7:0] p_43_1;
  input [7:0] p_43_2;
  input [7:0] p_43_3;
  input [7:0] p_43_4;
  input [7:0] p_43_5;
  input [7:0] p_43_6;
  input [7:0] p_43_7;
  input [7:0] p_43_8;
  input [7:0] p_43_9;
  input [7:0] p_43_10;
  input [7:0] p_43_11;
  input [7:0] p_43_12;
  input [7:0] p_43_13;
  input [7:0] p_43_14;
  input [7:0] p_43_15;
  input [7:0] p_43_16;
  input [7:0] p_43_17;
  input [7:0] p_43_18;
  input [7:0] p_43_19;
  input [7:0] p_43_20;
  input [7:0] p_43_21;
  input [7:0] p_43_22;
  input [7:0] p_43_23;
  input [7:0] p_43_24;
  input [7:0] p_43_25;
  input [7:0] p_43_26;
  input [7:0] p_43_27;
  input [7:0] p_43_28;
  input [7:0] p_43_29;
  input [7:0] p_43_30;
  input [7:0] p_43_31;
  input [7:0] p_43_32;
  input [7:0] p_43_33;
  input [7:0] p_43_34;
  input [7:0] p_43_35;
  input [7:0] p_43_36;
  input [7:0] p_43_37;
  input [7:0] p_43_38;
  input [7:0] p_43_39;
  input [7:0] p_43_40;
  input [7:0] p_43_41;
  input [7:0] p_43_42;
  input [7:0] p_43_43;
  input [7:0] p_43_44;
  input [7:0] p_43_45;
  input [7:0] p_43_46;
  input [7:0] p_43_47;
  input [7:0] p_43_48;
  input [7:0] p_43_49;
  input [7:0] p_43_50;
  input [7:0] p_43_51;
  input [7:0] p_43_52;
  input [7:0] p_43_53;
  input [7:0] p_43_54;
  input [7:0] p_43_55;
  input [7:0] p_43_56;
  input [7:0] p_43_57;
  input [7:0] p_43_58;
  input [7:0] p_43_59;
  input [7:0] p_43_60;
  input [7:0] p_43_61;
  input [7:0] p_43_62;
  input [7:0] p_43_63;
  input [7:0] p_43_64;
  input [7:0] p_43_65;
  input [7:0] p_44_0;
  input [7:0] p_44_1;
  input [7:0] p_44_2;
  input [7:0] p_44_3;
  input [7:0] p_44_4;
  input [7:0] p_44_5;
  input [7:0] p_44_6;
  input [7:0] p_44_7;
  input [7:0] p_44_8;
  input [7:0] p_44_9;
  input [7:0] p_44_10;
  input [7:0] p_44_11;
  input [7:0] p_44_12;
  input [7:0] p_44_13;
  input [7:0] p_44_14;
  input [7:0] p_44_15;
  input [7:0] p_44_16;
  input [7:0] p_44_17;
  input [7:0] p_44_18;
  input [7:0] p_44_19;
  input [7:0] p_44_20;
  input [7:0] p_44_21;
  input [7:0] p_44_22;
  input [7:0] p_44_23;
  input [7:0] p_44_24;
  input [7:0] p_44_25;
  input [7:0] p_44_26;
  input [7:0] p_44_27;
  input [7:0] p_44_28;
  input [7:0] p_44_29;
  input [7:0] p_44_30;
  input [7:0] p_44_31;
  input [7:0] p_44_32;
  input [7:0] p_44_33;
  input [7:0] p_44_34;
  input [7:0] p_44_35;
  input [7:0] p_44_36;
  input [7:0] p_44_37;
  input [7:0] p_44_38;
  input [7:0] p_44_39;
  input [7:0] p_44_40;
  input [7:0] p_44_41;
  input [7:0] p_44_42;
  input [7:0] p_44_43;
  input [7:0] p_44_44;
  input [7:0] p_44_45;
  input [7:0] p_44_46;
  input [7:0] p_44_47;
  input [7:0] p_44_48;
  input [7:0] p_44_49;
  input [7:0] p_44_50;
  input [7:0] p_44_51;
  input [7:0] p_44_52;
  input [7:0] p_44_53;
  input [7:0] p_44_54;
  input [7:0] p_44_55;
  input [7:0] p_44_56;
  input [7:0] p_44_57;
  input [7:0] p_44_58;
  input [7:0] p_44_59;
  input [7:0] p_44_60;
  input [7:0] p_44_61;
  input [7:0] p_44_62;
  input [7:0] p_44_63;
  input [7:0] p_44_64;
  input [7:0] p_44_65;

  output [7:0] out_1_1;
  output [7:0] out_1_2;
  output [7:0] out_1_3;
  output [7:0] out_1_4;
  output [7:0] out_1_5;
  output [7:0] out_1_6;
  output [7:0] out_1_7;
  output [7:0] out_1_8;
  output [7:0] out_1_9;
  output [7:0] out_1_10;
  output [7:0] out_1_11;
  output [7:0] out_1_12;
  output [7:0] out_1_13;
  output [7:0] out_1_14;
  output [7:0] out_1_15;
  output [7:0] out_1_16;
  output [7:0] out_1_17;
  output [7:0] out_1_18;
  output [7:0] out_1_19;
  output [7:0] out_1_20;
  output [7:0] out_1_21;
  output [7:0] out_1_22;
  output [7:0] out_1_23;
  output [7:0] out_1_24;
  output [7:0] out_1_25;
  output [7:0] out_1_26;
  output [7:0] out_1_27;
  output [7:0] out_1_28;
  output [7:0] out_1_29;
  output [7:0] out_1_30;
  output [7:0] out_1_31;
  output [7:0] out_1_32;
  output [7:0] out_1_33;
  output [7:0] out_1_34;
  output [7:0] out_1_35;
  output [7:0] out_1_36;
  output [7:0] out_1_37;
  output [7:0] out_1_38;
  output [7:0] out_1_39;
  output [7:0] out_1_40;
  output [7:0] out_1_41;
  output [7:0] out_1_42;
  output [7:0] out_1_43;
  output [7:0] out_1_44;
  output [7:0] out_1_45;
  output [7:0] out_1_46;
  output [7:0] out_1_47;
  output [7:0] out_1_48;
  output [7:0] out_1_49;
  output [7:0] out_1_50;
  output [7:0] out_1_51;
  output [7:0] out_1_52;
  output [7:0] out_1_53;
  output [7:0] out_1_54;
  output [7:0] out_1_55;
  output [7:0] out_1_56;
  output [7:0] out_1_57;
  output [7:0] out_1_58;
  output [7:0] out_1_59;
  output [7:0] out_1_60;
  output [7:0] out_1_61;
  output [7:0] out_1_62;
  output [7:0] out_1_63;
  output [7:0] out_1_64;
  output [7:0] out_2_1;
  output [7:0] out_2_2;
  output [7:0] out_2_3;
  output [7:0] out_2_4;
  output [7:0] out_2_5;
  output [7:0] out_2_6;
  output [7:0] out_2_7;
  output [7:0] out_2_8;
  output [7:0] out_2_9;
  output [7:0] out_2_10;
  output [7:0] out_2_11;
  output [7:0] out_2_12;
  output [7:0] out_2_13;
  output [7:0] out_2_14;
  output [7:0] out_2_15;
  output [7:0] out_2_16;
  output [7:0] out_2_17;
  output [7:0] out_2_18;
  output [7:0] out_2_19;
  output [7:0] out_2_20;
  output [7:0] out_2_21;
  output [7:0] out_2_22;
  output [7:0] out_2_23;
  output [7:0] out_2_24;
  output [7:0] out_2_25;
  output [7:0] out_2_26;
  output [7:0] out_2_27;
  output [7:0] out_2_28;
  output [7:0] out_2_29;
  output [7:0] out_2_30;
  output [7:0] out_2_31;
  output [7:0] out_2_32;
  output [7:0] out_2_33;
  output [7:0] out_2_34;
  output [7:0] out_2_35;
  output [7:0] out_2_36;
  output [7:0] out_2_37;
  output [7:0] out_2_38;
  output [7:0] out_2_39;
  output [7:0] out_2_40;
  output [7:0] out_2_41;
  output [7:0] out_2_42;
  output [7:0] out_2_43;
  output [7:0] out_2_44;
  output [7:0] out_2_45;
  output [7:0] out_2_46;
  output [7:0] out_2_47;
  output [7:0] out_2_48;
  output [7:0] out_2_49;
  output [7:0] out_2_50;
  output [7:0] out_2_51;
  output [7:0] out_2_52;
  output [7:0] out_2_53;
  output [7:0] out_2_54;
  output [7:0] out_2_55;
  output [7:0] out_2_56;
  output [7:0] out_2_57;
  output [7:0] out_2_58;
  output [7:0] out_2_59;
  output [7:0] out_2_60;
  output [7:0] out_2_61;
  output [7:0] out_2_62;
  output [7:0] out_2_63;
  output [7:0] out_2_64;
  output [7:0] out_3_1;
  output [7:0] out_3_2;
  output [7:0] out_3_3;
  output [7:0] out_3_4;
  output [7:0] out_3_5;
  output [7:0] out_3_6;
  output [7:0] out_3_7;
  output [7:0] out_3_8;
  output [7:0] out_3_9;
  output [7:0] out_3_10;
  output [7:0] out_3_11;
  output [7:0] out_3_12;
  output [7:0] out_3_13;
  output [7:0] out_3_14;
  output [7:0] out_3_15;
  output [7:0] out_3_16;
  output [7:0] out_3_17;
  output [7:0] out_3_18;
  output [7:0] out_3_19;
  output [7:0] out_3_20;
  output [7:0] out_3_21;
  output [7:0] out_3_22;
  output [7:0] out_3_23;
  output [7:0] out_3_24;
  output [7:0] out_3_25;
  output [7:0] out_3_26;
  output [7:0] out_3_27;
  output [7:0] out_3_28;
  output [7:0] out_3_29;
  output [7:0] out_3_30;
  output [7:0] out_3_31;
  output [7:0] out_3_32;
  output [7:0] out_3_33;
  output [7:0] out_3_34;
  output [7:0] out_3_35;
  output [7:0] out_3_36;
  output [7:0] out_3_37;
  output [7:0] out_3_38;
  output [7:0] out_3_39;
  output [7:0] out_3_40;
  output [7:0] out_3_41;
  output [7:0] out_3_42;
  output [7:0] out_3_43;
  output [7:0] out_3_44;
  output [7:0] out_3_45;
  output [7:0] out_3_46;
  output [7:0] out_3_47;
  output [7:0] out_3_48;
  output [7:0] out_3_49;
  output [7:0] out_3_50;
  output [7:0] out_3_51;
  output [7:0] out_3_52;
  output [7:0] out_3_53;
  output [7:0] out_3_54;
  output [7:0] out_3_55;
  output [7:0] out_3_56;
  output [7:0] out_3_57;
  output [7:0] out_3_58;
  output [7:0] out_3_59;
  output [7:0] out_3_60;
  output [7:0] out_3_61;
  output [7:0] out_3_62;
  output [7:0] out_3_63;
  output [7:0] out_3_64;
  output [7:0] out_4_1;
  output [7:0] out_4_2;
  output [7:0] out_4_3;
  output [7:0] out_4_4;
  output [7:0] out_4_5;
  output [7:0] out_4_6;
  output [7:0] out_4_7;
  output [7:0] out_4_8;
  output [7:0] out_4_9;
  output [7:0] out_4_10;
  output [7:0] out_4_11;
  output [7:0] out_4_12;
  output [7:0] out_4_13;
  output [7:0] out_4_14;
  output [7:0] out_4_15;
  output [7:0] out_4_16;
  output [7:0] out_4_17;
  output [7:0] out_4_18;
  output [7:0] out_4_19;
  output [7:0] out_4_20;
  output [7:0] out_4_21;
  output [7:0] out_4_22;
  output [7:0] out_4_23;
  output [7:0] out_4_24;
  output [7:0] out_4_25;
  output [7:0] out_4_26;
  output [7:0] out_4_27;
  output [7:0] out_4_28;
  output [7:0] out_4_29;
  output [7:0] out_4_30;
  output [7:0] out_4_31;
  output [7:0] out_4_32;
  output [7:0] out_4_33;
  output [7:0] out_4_34;
  output [7:0] out_4_35;
  output [7:0] out_4_36;
  output [7:0] out_4_37;
  output [7:0] out_4_38;
  output [7:0] out_4_39;
  output [7:0] out_4_40;
  output [7:0] out_4_41;
  output [7:0] out_4_42;
  output [7:0] out_4_43;
  output [7:0] out_4_44;
  output [7:0] out_4_45;
  output [7:0] out_4_46;
  output [7:0] out_4_47;
  output [7:0] out_4_48;
  output [7:0] out_4_49;
  output [7:0] out_4_50;
  output [7:0] out_4_51;
  output [7:0] out_4_52;
  output [7:0] out_4_53;
  output [7:0] out_4_54;
  output [7:0] out_4_55;
  output [7:0] out_4_56;
  output [7:0] out_4_57;
  output [7:0] out_4_58;
  output [7:0] out_4_59;
  output [7:0] out_4_60;
  output [7:0] out_4_61;
  output [7:0] out_4_62;
  output [7:0] out_4_63;
  output [7:0] out_4_64;
  output [7:0] out_5_1;
  output [7:0] out_5_2;
  output [7:0] out_5_3;
  output [7:0] out_5_4;
  output [7:0] out_5_5;
  output [7:0] out_5_6;
  output [7:0] out_5_7;
  output [7:0] out_5_8;
  output [7:0] out_5_9;
  output [7:0] out_5_10;
  output [7:0] out_5_11;
  output [7:0] out_5_12;
  output [7:0] out_5_13;
  output [7:0] out_5_14;
  output [7:0] out_5_15;
  output [7:0] out_5_16;
  output [7:0] out_5_17;
  output [7:0] out_5_18;
  output [7:0] out_5_19;
  output [7:0] out_5_20;
  output [7:0] out_5_21;
  output [7:0] out_5_22;
  output [7:0] out_5_23;
  output [7:0] out_5_24;
  output [7:0] out_5_25;
  output [7:0] out_5_26;
  output [7:0] out_5_27;
  output [7:0] out_5_28;
  output [7:0] out_5_29;
  output [7:0] out_5_30;
  output [7:0] out_5_31;
  output [7:0] out_5_32;
  output [7:0] out_5_33;
  output [7:0] out_5_34;
  output [7:0] out_5_35;
  output [7:0] out_5_36;
  output [7:0] out_5_37;
  output [7:0] out_5_38;
  output [7:0] out_5_39;
  output [7:0] out_5_40;
  output [7:0] out_5_41;
  output [7:0] out_5_42;
  output [7:0] out_5_43;
  output [7:0] out_5_44;
  output [7:0] out_5_45;
  output [7:0] out_5_46;
  output [7:0] out_5_47;
  output [7:0] out_5_48;
  output [7:0] out_5_49;
  output [7:0] out_5_50;
  output [7:0] out_5_51;
  output [7:0] out_5_52;
  output [7:0] out_5_53;
  output [7:0] out_5_54;
  output [7:0] out_5_55;
  output [7:0] out_5_56;
  output [7:0] out_5_57;
  output [7:0] out_5_58;
  output [7:0] out_5_59;
  output [7:0] out_5_60;
  output [7:0] out_5_61;
  output [7:0] out_5_62;
  output [7:0] out_5_63;
  output [7:0] out_5_64;
  output [7:0] out_6_1;
  output [7:0] out_6_2;
  output [7:0] out_6_3;
  output [7:0] out_6_4;
  output [7:0] out_6_5;
  output [7:0] out_6_6;
  output [7:0] out_6_7;
  output [7:0] out_6_8;
  output [7:0] out_6_9;
  output [7:0] out_6_10;
  output [7:0] out_6_11;
  output [7:0] out_6_12;
  output [7:0] out_6_13;
  output [7:0] out_6_14;
  output [7:0] out_6_15;
  output [7:0] out_6_16;
  output [7:0] out_6_17;
  output [7:0] out_6_18;
  output [7:0] out_6_19;
  output [7:0] out_6_20;
  output [7:0] out_6_21;
  output [7:0] out_6_22;
  output [7:0] out_6_23;
  output [7:0] out_6_24;
  output [7:0] out_6_25;
  output [7:0] out_6_26;
  output [7:0] out_6_27;
  output [7:0] out_6_28;
  output [7:0] out_6_29;
  output [7:0] out_6_30;
  output [7:0] out_6_31;
  output [7:0] out_6_32;
  output [7:0] out_6_33;
  output [7:0] out_6_34;
  output [7:0] out_6_35;
  output [7:0] out_6_36;
  output [7:0] out_6_37;
  output [7:0] out_6_38;
  output [7:0] out_6_39;
  output [7:0] out_6_40;
  output [7:0] out_6_41;
  output [7:0] out_6_42;
  output [7:0] out_6_43;
  output [7:0] out_6_44;
  output [7:0] out_6_45;
  output [7:0] out_6_46;
  output [7:0] out_6_47;
  output [7:0] out_6_48;
  output [7:0] out_6_49;
  output [7:0] out_6_50;
  output [7:0] out_6_51;
  output [7:0] out_6_52;
  output [7:0] out_6_53;
  output [7:0] out_6_54;
  output [7:0] out_6_55;
  output [7:0] out_6_56;
  output [7:0] out_6_57;
  output [7:0] out_6_58;
  output [7:0] out_6_59;
  output [7:0] out_6_60;
  output [7:0] out_6_61;
  output [7:0] out_6_62;
  output [7:0] out_6_63;
  output [7:0] out_6_64;
  output [7:0] out_7_1;
  output [7:0] out_7_2;
  output [7:0] out_7_3;
  output [7:0] out_7_4;
  output [7:0] out_7_5;
  output [7:0] out_7_6;
  output [7:0] out_7_7;
  output [7:0] out_7_8;
  output [7:0] out_7_9;
  output [7:0] out_7_10;
  output [7:0] out_7_11;
  output [7:0] out_7_12;
  output [7:0] out_7_13;
  output [7:0] out_7_14;
  output [7:0] out_7_15;
  output [7:0] out_7_16;
  output [7:0] out_7_17;
  output [7:0] out_7_18;
  output [7:0] out_7_19;
  output [7:0] out_7_20;
  output [7:0] out_7_21;
  output [7:0] out_7_22;
  output [7:0] out_7_23;
  output [7:0] out_7_24;
  output [7:0] out_7_25;
  output [7:0] out_7_26;
  output [7:0] out_7_27;
  output [7:0] out_7_28;
  output [7:0] out_7_29;
  output [7:0] out_7_30;
  output [7:0] out_7_31;
  output [7:0] out_7_32;
  output [7:0] out_7_33;
  output [7:0] out_7_34;
  output [7:0] out_7_35;
  output [7:0] out_7_36;
  output [7:0] out_7_37;
  output [7:0] out_7_38;
  output [7:0] out_7_39;
  output [7:0] out_7_40;
  output [7:0] out_7_41;
  output [7:0] out_7_42;
  output [7:0] out_7_43;
  output [7:0] out_7_44;
  output [7:0] out_7_45;
  output [7:0] out_7_46;
  output [7:0] out_7_47;
  output [7:0] out_7_48;
  output [7:0] out_7_49;
  output [7:0] out_7_50;
  output [7:0] out_7_51;
  output [7:0] out_7_52;
  output [7:0] out_7_53;
  output [7:0] out_7_54;
  output [7:0] out_7_55;
  output [7:0] out_7_56;
  output [7:0] out_7_57;
  output [7:0] out_7_58;
  output [7:0] out_7_59;
  output [7:0] out_7_60;
  output [7:0] out_7_61;
  output [7:0] out_7_62;
  output [7:0] out_7_63;
  output [7:0] out_7_64;
  output [7:0] out_8_1;
  output [7:0] out_8_2;
  output [7:0] out_8_3;
  output [7:0] out_8_4;
  output [7:0] out_8_5;
  output [7:0] out_8_6;
  output [7:0] out_8_7;
  output [7:0] out_8_8;
  output [7:0] out_8_9;
  output [7:0] out_8_10;
  output [7:0] out_8_11;
  output [7:0] out_8_12;
  output [7:0] out_8_13;
  output [7:0] out_8_14;
  output [7:0] out_8_15;
  output [7:0] out_8_16;
  output [7:0] out_8_17;
  output [7:0] out_8_18;
  output [7:0] out_8_19;
  output [7:0] out_8_20;
  output [7:0] out_8_21;
  output [7:0] out_8_22;
  output [7:0] out_8_23;
  output [7:0] out_8_24;
  output [7:0] out_8_25;
  output [7:0] out_8_26;
  output [7:0] out_8_27;
  output [7:0] out_8_28;
  output [7:0] out_8_29;
  output [7:0] out_8_30;
  output [7:0] out_8_31;
  output [7:0] out_8_32;
  output [7:0] out_8_33;
  output [7:0] out_8_34;
  output [7:0] out_8_35;
  output [7:0] out_8_36;
  output [7:0] out_8_37;
  output [7:0] out_8_38;
  output [7:0] out_8_39;
  output [7:0] out_8_40;
  output [7:0] out_8_41;
  output [7:0] out_8_42;
  output [7:0] out_8_43;
  output [7:0] out_8_44;
  output [7:0] out_8_45;
  output [7:0] out_8_46;
  output [7:0] out_8_47;
  output [7:0] out_8_48;
  output [7:0] out_8_49;
  output [7:0] out_8_50;
  output [7:0] out_8_51;
  output [7:0] out_8_52;
  output [7:0] out_8_53;
  output [7:0] out_8_54;
  output [7:0] out_8_55;
  output [7:0] out_8_56;
  output [7:0] out_8_57;
  output [7:0] out_8_58;
  output [7:0] out_8_59;
  output [7:0] out_8_60;
  output [7:0] out_8_61;
  output [7:0] out_8_62;
  output [7:0] out_8_63;
  output [7:0] out_8_64;
  output [7:0] out_9_1;
  output [7:0] out_9_2;
  output [7:0] out_9_3;
  output [7:0] out_9_4;
  output [7:0] out_9_5;
  output [7:0] out_9_6;
  output [7:0] out_9_7;
  output [7:0] out_9_8;
  output [7:0] out_9_9;
  output [7:0] out_9_10;
  output [7:0] out_9_11;
  output [7:0] out_9_12;
  output [7:0] out_9_13;
  output [7:0] out_9_14;
  output [7:0] out_9_15;
  output [7:0] out_9_16;
  output [7:0] out_9_17;
  output [7:0] out_9_18;
  output [7:0] out_9_19;
  output [7:0] out_9_20;
  output [7:0] out_9_21;
  output [7:0] out_9_22;
  output [7:0] out_9_23;
  output [7:0] out_9_24;
  output [7:0] out_9_25;
  output [7:0] out_9_26;
  output [7:0] out_9_27;
  output [7:0] out_9_28;
  output [7:0] out_9_29;
  output [7:0] out_9_30;
  output [7:0] out_9_31;
  output [7:0] out_9_32;
  output [7:0] out_9_33;
  output [7:0] out_9_34;
  output [7:0] out_9_35;
  output [7:0] out_9_36;
  output [7:0] out_9_37;
  output [7:0] out_9_38;
  output [7:0] out_9_39;
  output [7:0] out_9_40;
  output [7:0] out_9_41;
  output [7:0] out_9_42;
  output [7:0] out_9_43;
  output [7:0] out_9_44;
  output [7:0] out_9_45;
  output [7:0] out_9_46;
  output [7:0] out_9_47;
  output [7:0] out_9_48;
  output [7:0] out_9_49;
  output [7:0] out_9_50;
  output [7:0] out_9_51;
  output [7:0] out_9_52;
  output [7:0] out_9_53;
  output [7:0] out_9_54;
  output [7:0] out_9_55;
  output [7:0] out_9_56;
  output [7:0] out_9_57;
  output [7:0] out_9_58;
  output [7:0] out_9_59;
  output [7:0] out_9_60;
  output [7:0] out_9_61;
  output [7:0] out_9_62;
  output [7:0] out_9_63;
  output [7:0] out_9_64;
  output [7:0] out_10_1;
  output [7:0] out_10_2;
  output [7:0] out_10_3;
  output [7:0] out_10_4;
  output [7:0] out_10_5;
  output [7:0] out_10_6;
  output [7:0] out_10_7;
  output [7:0] out_10_8;
  output [7:0] out_10_9;
  output [7:0] out_10_10;
  output [7:0] out_10_11;
  output [7:0] out_10_12;
  output [7:0] out_10_13;
  output [7:0] out_10_14;
  output [7:0] out_10_15;
  output [7:0] out_10_16;
  output [7:0] out_10_17;
  output [7:0] out_10_18;
  output [7:0] out_10_19;
  output [7:0] out_10_20;
  output [7:0] out_10_21;
  output [7:0] out_10_22;
  output [7:0] out_10_23;
  output [7:0] out_10_24;
  output [7:0] out_10_25;
  output [7:0] out_10_26;
  output [7:0] out_10_27;
  output [7:0] out_10_28;
  output [7:0] out_10_29;
  output [7:0] out_10_30;
  output [7:0] out_10_31;
  output [7:0] out_10_32;
  output [7:0] out_10_33;
  output [7:0] out_10_34;
  output [7:0] out_10_35;
  output [7:0] out_10_36;
  output [7:0] out_10_37;
  output [7:0] out_10_38;
  output [7:0] out_10_39;
  output [7:0] out_10_40;
  output [7:0] out_10_41;
  output [7:0] out_10_42;
  output [7:0] out_10_43;
  output [7:0] out_10_44;
  output [7:0] out_10_45;
  output [7:0] out_10_46;
  output [7:0] out_10_47;
  output [7:0] out_10_48;
  output [7:0] out_10_49;
  output [7:0] out_10_50;
  output [7:0] out_10_51;
  output [7:0] out_10_52;
  output [7:0] out_10_53;
  output [7:0] out_10_54;
  output [7:0] out_10_55;
  output [7:0] out_10_56;
  output [7:0] out_10_57;
  output [7:0] out_10_58;
  output [7:0] out_10_59;
  output [7:0] out_10_60;
  output [7:0] out_10_61;
  output [7:0] out_10_62;
  output [7:0] out_10_63;
  output [7:0] out_10_64;
  output [7:0] out_11_1;
  output [7:0] out_11_2;
  output [7:0] out_11_3;
  output [7:0] out_11_4;
  output [7:0] out_11_5;
  output [7:0] out_11_6;
  output [7:0] out_11_7;
  output [7:0] out_11_8;
  output [7:0] out_11_9;
  output [7:0] out_11_10;
  output [7:0] out_11_11;
  output [7:0] out_11_12;
  output [7:0] out_11_13;
  output [7:0] out_11_14;
  output [7:0] out_11_15;
  output [7:0] out_11_16;
  output [7:0] out_11_17;
  output [7:0] out_11_18;
  output [7:0] out_11_19;
  output [7:0] out_11_20;
  output [7:0] out_11_21;
  output [7:0] out_11_22;
  output [7:0] out_11_23;
  output [7:0] out_11_24;
  output [7:0] out_11_25;
  output [7:0] out_11_26;
  output [7:0] out_11_27;
  output [7:0] out_11_28;
  output [7:0] out_11_29;
  output [7:0] out_11_30;
  output [7:0] out_11_31;
  output [7:0] out_11_32;
  output [7:0] out_11_33;
  output [7:0] out_11_34;
  output [7:0] out_11_35;
  output [7:0] out_11_36;
  output [7:0] out_11_37;
  output [7:0] out_11_38;
  output [7:0] out_11_39;
  output [7:0] out_11_40;
  output [7:0] out_11_41;
  output [7:0] out_11_42;
  output [7:0] out_11_43;
  output [7:0] out_11_44;
  output [7:0] out_11_45;
  output [7:0] out_11_46;
  output [7:0] out_11_47;
  output [7:0] out_11_48;
  output [7:0] out_11_49;
  output [7:0] out_11_50;
  output [7:0] out_11_51;
  output [7:0] out_11_52;
  output [7:0] out_11_53;
  output [7:0] out_11_54;
  output [7:0] out_11_55;
  output [7:0] out_11_56;
  output [7:0] out_11_57;
  output [7:0] out_11_58;
  output [7:0] out_11_59;
  output [7:0] out_11_60;
  output [7:0] out_11_61;
  output [7:0] out_11_62;
  output [7:0] out_11_63;
  output [7:0] out_11_64;
  output [7:0] out_12_1;
  output [7:0] out_12_2;
  output [7:0] out_12_3;
  output [7:0] out_12_4;
  output [7:0] out_12_5;
  output [7:0] out_12_6;
  output [7:0] out_12_7;
  output [7:0] out_12_8;
  output [7:0] out_12_9;
  output [7:0] out_12_10;
  output [7:0] out_12_11;
  output [7:0] out_12_12;
  output [7:0] out_12_13;
  output [7:0] out_12_14;
  output [7:0] out_12_15;
  output [7:0] out_12_16;
  output [7:0] out_12_17;
  output [7:0] out_12_18;
  output [7:0] out_12_19;
  output [7:0] out_12_20;
  output [7:0] out_12_21;
  output [7:0] out_12_22;
  output [7:0] out_12_23;
  output [7:0] out_12_24;
  output [7:0] out_12_25;
  output [7:0] out_12_26;
  output [7:0] out_12_27;
  output [7:0] out_12_28;
  output [7:0] out_12_29;
  output [7:0] out_12_30;
  output [7:0] out_12_31;
  output [7:0] out_12_32;
  output [7:0] out_12_33;
  output [7:0] out_12_34;
  output [7:0] out_12_35;
  output [7:0] out_12_36;
  output [7:0] out_12_37;
  output [7:0] out_12_38;
  output [7:0] out_12_39;
  output [7:0] out_12_40;
  output [7:0] out_12_41;
  output [7:0] out_12_42;
  output [7:0] out_12_43;
  output [7:0] out_12_44;
  output [7:0] out_12_45;
  output [7:0] out_12_46;
  output [7:0] out_12_47;
  output [7:0] out_12_48;
  output [7:0] out_12_49;
  output [7:0] out_12_50;
  output [7:0] out_12_51;
  output [7:0] out_12_52;
  output [7:0] out_12_53;
  output [7:0] out_12_54;
  output [7:0] out_12_55;
  output [7:0] out_12_56;
  output [7:0] out_12_57;
  output [7:0] out_12_58;
  output [7:0] out_12_59;
  output [7:0] out_12_60;
  output [7:0] out_12_61;
  output [7:0] out_12_62;
  output [7:0] out_12_63;
  output [7:0] out_12_64;
  output [7:0] out_13_1;
  output [7:0] out_13_2;
  output [7:0] out_13_3;
  output [7:0] out_13_4;
  output [7:0] out_13_5;
  output [7:0] out_13_6;
  output [7:0] out_13_7;
  output [7:0] out_13_8;
  output [7:0] out_13_9;
  output [7:0] out_13_10;
  output [7:0] out_13_11;
  output [7:0] out_13_12;
  output [7:0] out_13_13;
  output [7:0] out_13_14;
  output [7:0] out_13_15;
  output [7:0] out_13_16;
  output [7:0] out_13_17;
  output [7:0] out_13_18;
  output [7:0] out_13_19;
  output [7:0] out_13_20;
  output [7:0] out_13_21;
  output [7:0] out_13_22;
  output [7:0] out_13_23;
  output [7:0] out_13_24;
  output [7:0] out_13_25;
  output [7:0] out_13_26;
  output [7:0] out_13_27;
  output [7:0] out_13_28;
  output [7:0] out_13_29;
  output [7:0] out_13_30;
  output [7:0] out_13_31;
  output [7:0] out_13_32;
  output [7:0] out_13_33;
  output [7:0] out_13_34;
  output [7:0] out_13_35;
  output [7:0] out_13_36;
  output [7:0] out_13_37;
  output [7:0] out_13_38;
  output [7:0] out_13_39;
  output [7:0] out_13_40;
  output [7:0] out_13_41;
  output [7:0] out_13_42;
  output [7:0] out_13_43;
  output [7:0] out_13_44;
  output [7:0] out_13_45;
  output [7:0] out_13_46;
  output [7:0] out_13_47;
  output [7:0] out_13_48;
  output [7:0] out_13_49;
  output [7:0] out_13_50;
  output [7:0] out_13_51;
  output [7:0] out_13_52;
  output [7:0] out_13_53;
  output [7:0] out_13_54;
  output [7:0] out_13_55;
  output [7:0] out_13_56;
  output [7:0] out_13_57;
  output [7:0] out_13_58;
  output [7:0] out_13_59;
  output [7:0] out_13_60;
  output [7:0] out_13_61;
  output [7:0] out_13_62;
  output [7:0] out_13_63;
  output [7:0] out_13_64;
  output [7:0] out_14_1;
  output [7:0] out_14_2;
  output [7:0] out_14_3;
  output [7:0] out_14_4;
  output [7:0] out_14_5;
  output [7:0] out_14_6;
  output [7:0] out_14_7;
  output [7:0] out_14_8;
  output [7:0] out_14_9;
  output [7:0] out_14_10;
  output [7:0] out_14_11;
  output [7:0] out_14_12;
  output [7:0] out_14_13;
  output [7:0] out_14_14;
  output [7:0] out_14_15;
  output [7:0] out_14_16;
  output [7:0] out_14_17;
  output [7:0] out_14_18;
  output [7:0] out_14_19;
  output [7:0] out_14_20;
  output [7:0] out_14_21;
  output [7:0] out_14_22;
  output [7:0] out_14_23;
  output [7:0] out_14_24;
  output [7:0] out_14_25;
  output [7:0] out_14_26;
  output [7:0] out_14_27;
  output [7:0] out_14_28;
  output [7:0] out_14_29;
  output [7:0] out_14_30;
  output [7:0] out_14_31;
  output [7:0] out_14_32;
  output [7:0] out_14_33;
  output [7:0] out_14_34;
  output [7:0] out_14_35;
  output [7:0] out_14_36;
  output [7:0] out_14_37;
  output [7:0] out_14_38;
  output [7:0] out_14_39;
  output [7:0] out_14_40;
  output [7:0] out_14_41;
  output [7:0] out_14_42;
  output [7:0] out_14_43;
  output [7:0] out_14_44;
  output [7:0] out_14_45;
  output [7:0] out_14_46;
  output [7:0] out_14_47;
  output [7:0] out_14_48;
  output [7:0] out_14_49;
  output [7:0] out_14_50;
  output [7:0] out_14_51;
  output [7:0] out_14_52;
  output [7:0] out_14_53;
  output [7:0] out_14_54;
  output [7:0] out_14_55;
  output [7:0] out_14_56;
  output [7:0] out_14_57;
  output [7:0] out_14_58;
  output [7:0] out_14_59;
  output [7:0] out_14_60;
  output [7:0] out_14_61;
  output [7:0] out_14_62;
  output [7:0] out_14_63;
  output [7:0] out_14_64;
  output [7:0] out_15_1;
  output [7:0] out_15_2;
  output [7:0] out_15_3;
  output [7:0] out_15_4;
  output [7:0] out_15_5;
  output [7:0] out_15_6;
  output [7:0] out_15_7;
  output [7:0] out_15_8;
  output [7:0] out_15_9;
  output [7:0] out_15_10;
  output [7:0] out_15_11;
  output [7:0] out_15_12;
  output [7:0] out_15_13;
  output [7:0] out_15_14;
  output [7:0] out_15_15;
  output [7:0] out_15_16;
  output [7:0] out_15_17;
  output [7:0] out_15_18;
  output [7:0] out_15_19;
  output [7:0] out_15_20;
  output [7:0] out_15_21;
  output [7:0] out_15_22;
  output [7:0] out_15_23;
  output [7:0] out_15_24;
  output [7:0] out_15_25;
  output [7:0] out_15_26;
  output [7:0] out_15_27;
  output [7:0] out_15_28;
  output [7:0] out_15_29;
  output [7:0] out_15_30;
  output [7:0] out_15_31;
  output [7:0] out_15_32;
  output [7:0] out_15_33;
  output [7:0] out_15_34;
  output [7:0] out_15_35;
  output [7:0] out_15_36;
  output [7:0] out_15_37;
  output [7:0] out_15_38;
  output [7:0] out_15_39;
  output [7:0] out_15_40;
  output [7:0] out_15_41;
  output [7:0] out_15_42;
  output [7:0] out_15_43;
  output [7:0] out_15_44;
  output [7:0] out_15_45;
  output [7:0] out_15_46;
  output [7:0] out_15_47;
  output [7:0] out_15_48;
  output [7:0] out_15_49;
  output [7:0] out_15_50;
  output [7:0] out_15_51;
  output [7:0] out_15_52;
  output [7:0] out_15_53;
  output [7:0] out_15_54;
  output [7:0] out_15_55;
  output [7:0] out_15_56;
  output [7:0] out_15_57;
  output [7:0] out_15_58;
  output [7:0] out_15_59;
  output [7:0] out_15_60;
  output [7:0] out_15_61;
  output [7:0] out_15_62;
  output [7:0] out_15_63;
  output [7:0] out_15_64;
  output [7:0] out_16_1;
  output [7:0] out_16_2;
  output [7:0] out_16_3;
  output [7:0] out_16_4;
  output [7:0] out_16_5;
  output [7:0] out_16_6;
  output [7:0] out_16_7;
  output [7:0] out_16_8;
  output [7:0] out_16_9;
  output [7:0] out_16_10;
  output [7:0] out_16_11;
  output [7:0] out_16_12;
  output [7:0] out_16_13;
  output [7:0] out_16_14;
  output [7:0] out_16_15;
  output [7:0] out_16_16;
  output [7:0] out_16_17;
  output [7:0] out_16_18;
  output [7:0] out_16_19;
  output [7:0] out_16_20;
  output [7:0] out_16_21;
  output [7:0] out_16_22;
  output [7:0] out_16_23;
  output [7:0] out_16_24;
  output [7:0] out_16_25;
  output [7:0] out_16_26;
  output [7:0] out_16_27;
  output [7:0] out_16_28;
  output [7:0] out_16_29;
  output [7:0] out_16_30;
  output [7:0] out_16_31;
  output [7:0] out_16_32;
  output [7:0] out_16_33;
  output [7:0] out_16_34;
  output [7:0] out_16_35;
  output [7:0] out_16_36;
  output [7:0] out_16_37;
  output [7:0] out_16_38;
  output [7:0] out_16_39;
  output [7:0] out_16_40;
  output [7:0] out_16_41;
  output [7:0] out_16_42;
  output [7:0] out_16_43;
  output [7:0] out_16_44;
  output [7:0] out_16_45;
  output [7:0] out_16_46;
  output [7:0] out_16_47;
  output [7:0] out_16_48;
  output [7:0] out_16_49;
  output [7:0] out_16_50;
  output [7:0] out_16_51;
  output [7:0] out_16_52;
  output [7:0] out_16_53;
  output [7:0] out_16_54;
  output [7:0] out_16_55;
  output [7:0] out_16_56;
  output [7:0] out_16_57;
  output [7:0] out_16_58;
  output [7:0] out_16_59;
  output [7:0] out_16_60;
  output [7:0] out_16_61;
  output [7:0] out_16_62;
  output [7:0] out_16_63;
  output [7:0] out_16_64;
  output [7:0] out_17_1;
  output [7:0] out_17_2;
  output [7:0] out_17_3;
  output [7:0] out_17_4;
  output [7:0] out_17_5;
  output [7:0] out_17_6;
  output [7:0] out_17_7;
  output [7:0] out_17_8;
  output [7:0] out_17_9;
  output [7:0] out_17_10;
  output [7:0] out_17_11;
  output [7:0] out_17_12;
  output [7:0] out_17_13;
  output [7:0] out_17_14;
  output [7:0] out_17_15;
  output [7:0] out_17_16;
  output [7:0] out_17_17;
  output [7:0] out_17_18;
  output [7:0] out_17_19;
  output [7:0] out_17_20;
  output [7:0] out_17_21;
  output [7:0] out_17_22;
  output [7:0] out_17_23;
  output [7:0] out_17_24;
  output [7:0] out_17_25;
  output [7:0] out_17_26;
  output [7:0] out_17_27;
  output [7:0] out_17_28;
  output [7:0] out_17_29;
  output [7:0] out_17_30;
  output [7:0] out_17_31;
  output [7:0] out_17_32;
  output [7:0] out_17_33;
  output [7:0] out_17_34;
  output [7:0] out_17_35;
  output [7:0] out_17_36;
  output [7:0] out_17_37;
  output [7:0] out_17_38;
  output [7:0] out_17_39;
  output [7:0] out_17_40;
  output [7:0] out_17_41;
  output [7:0] out_17_42;
  output [7:0] out_17_43;
  output [7:0] out_17_44;
  output [7:0] out_17_45;
  output [7:0] out_17_46;
  output [7:0] out_17_47;
  output [7:0] out_17_48;
  output [7:0] out_17_49;
  output [7:0] out_17_50;
  output [7:0] out_17_51;
  output [7:0] out_17_52;
  output [7:0] out_17_53;
  output [7:0] out_17_54;
  output [7:0] out_17_55;
  output [7:0] out_17_56;
  output [7:0] out_17_57;
  output [7:0] out_17_58;
  output [7:0] out_17_59;
  output [7:0] out_17_60;
  output [7:0] out_17_61;
  output [7:0] out_17_62;
  output [7:0] out_17_63;
  output [7:0] out_17_64;
  output [7:0] out_18_1;
  output [7:0] out_18_2;
  output [7:0] out_18_3;
  output [7:0] out_18_4;
  output [7:0] out_18_5;
  output [7:0] out_18_6;
  output [7:0] out_18_7;
  output [7:0] out_18_8;
  output [7:0] out_18_9;
  output [7:0] out_18_10;
  output [7:0] out_18_11;
  output [7:0] out_18_12;
  output [7:0] out_18_13;
  output [7:0] out_18_14;
  output [7:0] out_18_15;
  output [7:0] out_18_16;
  output [7:0] out_18_17;
  output [7:0] out_18_18;
  output [7:0] out_18_19;
  output [7:0] out_18_20;
  output [7:0] out_18_21;
  output [7:0] out_18_22;
  output [7:0] out_18_23;
  output [7:0] out_18_24;
  output [7:0] out_18_25;
  output [7:0] out_18_26;
  output [7:0] out_18_27;
  output [7:0] out_18_28;
  output [7:0] out_18_29;
  output [7:0] out_18_30;
  output [7:0] out_18_31;
  output [7:0] out_18_32;
  output [7:0] out_18_33;
  output [7:0] out_18_34;
  output [7:0] out_18_35;
  output [7:0] out_18_36;
  output [7:0] out_18_37;
  output [7:0] out_18_38;
  output [7:0] out_18_39;
  output [7:0] out_18_40;
  output [7:0] out_18_41;
  output [7:0] out_18_42;
  output [7:0] out_18_43;
  output [7:0] out_18_44;
  output [7:0] out_18_45;
  output [7:0] out_18_46;
  output [7:0] out_18_47;
  output [7:0] out_18_48;
  output [7:0] out_18_49;
  output [7:0] out_18_50;
  output [7:0] out_18_51;
  output [7:0] out_18_52;
  output [7:0] out_18_53;
  output [7:0] out_18_54;
  output [7:0] out_18_55;
  output [7:0] out_18_56;
  output [7:0] out_18_57;
  output [7:0] out_18_58;
  output [7:0] out_18_59;
  output [7:0] out_18_60;
  output [7:0] out_18_61;
  output [7:0] out_18_62;
  output [7:0] out_18_63;
  output [7:0] out_18_64;
  output [7:0] out_19_1;
  output [7:0] out_19_2;
  output [7:0] out_19_3;
  output [7:0] out_19_4;
  output [7:0] out_19_5;
  output [7:0] out_19_6;
  output [7:0] out_19_7;
  output [7:0] out_19_8;
  output [7:0] out_19_9;
  output [7:0] out_19_10;
  output [7:0] out_19_11;
  output [7:0] out_19_12;
  output [7:0] out_19_13;
  output [7:0] out_19_14;
  output [7:0] out_19_15;
  output [7:0] out_19_16;
  output [7:0] out_19_17;
  output [7:0] out_19_18;
  output [7:0] out_19_19;
  output [7:0] out_19_20;
  output [7:0] out_19_21;
  output [7:0] out_19_22;
  output [7:0] out_19_23;
  output [7:0] out_19_24;
  output [7:0] out_19_25;
  output [7:0] out_19_26;
  output [7:0] out_19_27;
  output [7:0] out_19_28;
  output [7:0] out_19_29;
  output [7:0] out_19_30;
  output [7:0] out_19_31;
  output [7:0] out_19_32;
  output [7:0] out_19_33;
  output [7:0] out_19_34;
  output [7:0] out_19_35;
  output [7:0] out_19_36;
  output [7:0] out_19_37;
  output [7:0] out_19_38;
  output [7:0] out_19_39;
  output [7:0] out_19_40;
  output [7:0] out_19_41;
  output [7:0] out_19_42;
  output [7:0] out_19_43;
  output [7:0] out_19_44;
  output [7:0] out_19_45;
  output [7:0] out_19_46;
  output [7:0] out_19_47;
  output [7:0] out_19_48;
  output [7:0] out_19_49;
  output [7:0] out_19_50;
  output [7:0] out_19_51;
  output [7:0] out_19_52;
  output [7:0] out_19_53;
  output [7:0] out_19_54;
  output [7:0] out_19_55;
  output [7:0] out_19_56;
  output [7:0] out_19_57;
  output [7:0] out_19_58;
  output [7:0] out_19_59;
  output [7:0] out_19_60;
  output [7:0] out_19_61;
  output [7:0] out_19_62;
  output [7:0] out_19_63;
  output [7:0] out_19_64;
  output [7:0] out_20_1;
  output [7:0] out_20_2;
  output [7:0] out_20_3;
  output [7:0] out_20_4;
  output [7:0] out_20_5;
  output [7:0] out_20_6;
  output [7:0] out_20_7;
  output [7:0] out_20_8;
  output [7:0] out_20_9;
  output [7:0] out_20_10;
  output [7:0] out_20_11;
  output [7:0] out_20_12;
  output [7:0] out_20_13;
  output [7:0] out_20_14;
  output [7:0] out_20_15;
  output [7:0] out_20_16;
  output [7:0] out_20_17;
  output [7:0] out_20_18;
  output [7:0] out_20_19;
  output [7:0] out_20_20;
  output [7:0] out_20_21;
  output [7:0] out_20_22;
  output [7:0] out_20_23;
  output [7:0] out_20_24;
  output [7:0] out_20_25;
  output [7:0] out_20_26;
  output [7:0] out_20_27;
  output [7:0] out_20_28;
  output [7:0] out_20_29;
  output [7:0] out_20_30;
  output [7:0] out_20_31;
  output [7:0] out_20_32;
  output [7:0] out_20_33;
  output [7:0] out_20_34;
  output [7:0] out_20_35;
  output [7:0] out_20_36;
  output [7:0] out_20_37;
  output [7:0] out_20_38;
  output [7:0] out_20_39;
  output [7:0] out_20_40;
  output [7:0] out_20_41;
  output [7:0] out_20_42;
  output [7:0] out_20_43;
  output [7:0] out_20_44;
  output [7:0] out_20_45;
  output [7:0] out_20_46;
  output [7:0] out_20_47;
  output [7:0] out_20_48;
  output [7:0] out_20_49;
  output [7:0] out_20_50;
  output [7:0] out_20_51;
  output [7:0] out_20_52;
  output [7:0] out_20_53;
  output [7:0] out_20_54;
  output [7:0] out_20_55;
  output [7:0] out_20_56;
  output [7:0] out_20_57;
  output [7:0] out_20_58;
  output [7:0] out_20_59;
  output [7:0] out_20_60;
  output [7:0] out_20_61;
  output [7:0] out_20_62;
  output [7:0] out_20_63;
  output [7:0] out_20_64;
  output [7:0] out_21_1;
  output [7:0] out_21_2;
  output [7:0] out_21_3;
  output [7:0] out_21_4;
  output [7:0] out_21_5;
  output [7:0] out_21_6;
  output [7:0] out_21_7;
  output [7:0] out_21_8;
  output [7:0] out_21_9;
  output [7:0] out_21_10;
  output [7:0] out_21_11;
  output [7:0] out_21_12;
  output [7:0] out_21_13;
  output [7:0] out_21_14;
  output [7:0] out_21_15;
  output [7:0] out_21_16;
  output [7:0] out_21_17;
  output [7:0] out_21_18;
  output [7:0] out_21_19;
  output [7:0] out_21_20;
  output [7:0] out_21_21;
  output [7:0] out_21_22;
  output [7:0] out_21_23;
  output [7:0] out_21_24;
  output [7:0] out_21_25;
  output [7:0] out_21_26;
  output [7:0] out_21_27;
  output [7:0] out_21_28;
  output [7:0] out_21_29;
  output [7:0] out_21_30;
  output [7:0] out_21_31;
  output [7:0] out_21_32;
  output [7:0] out_21_33;
  output [7:0] out_21_34;
  output [7:0] out_21_35;
  output [7:0] out_21_36;
  output [7:0] out_21_37;
  output [7:0] out_21_38;
  output [7:0] out_21_39;
  output [7:0] out_21_40;
  output [7:0] out_21_41;
  output [7:0] out_21_42;
  output [7:0] out_21_43;
  output [7:0] out_21_44;
  output [7:0] out_21_45;
  output [7:0] out_21_46;
  output [7:0] out_21_47;
  output [7:0] out_21_48;
  output [7:0] out_21_49;
  output [7:0] out_21_50;
  output [7:0] out_21_51;
  output [7:0] out_21_52;
  output [7:0] out_21_53;
  output [7:0] out_21_54;
  output [7:0] out_21_55;
  output [7:0] out_21_56;
  output [7:0] out_21_57;
  output [7:0] out_21_58;
  output [7:0] out_21_59;
  output [7:0] out_21_60;
  output [7:0] out_21_61;
  output [7:0] out_21_62;
  output [7:0] out_21_63;
  output [7:0] out_21_64;
  output [7:0] out_22_1;
  output [7:0] out_22_2;
  output [7:0] out_22_3;
  output [7:0] out_22_4;
  output [7:0] out_22_5;
  output [7:0] out_22_6;
  output [7:0] out_22_7;
  output [7:0] out_22_8;
  output [7:0] out_22_9;
  output [7:0] out_22_10;
  output [7:0] out_22_11;
  output [7:0] out_22_12;
  output [7:0] out_22_13;
  output [7:0] out_22_14;
  output [7:0] out_22_15;
  output [7:0] out_22_16;
  output [7:0] out_22_17;
  output [7:0] out_22_18;
  output [7:0] out_22_19;
  output [7:0] out_22_20;
  output [7:0] out_22_21;
  output [7:0] out_22_22;
  output [7:0] out_22_23;
  output [7:0] out_22_24;
  output [7:0] out_22_25;
  output [7:0] out_22_26;
  output [7:0] out_22_27;
  output [7:0] out_22_28;
  output [7:0] out_22_29;
  output [7:0] out_22_30;
  output [7:0] out_22_31;
  output [7:0] out_22_32;
  output [7:0] out_22_33;
  output [7:0] out_22_34;
  output [7:0] out_22_35;
  output [7:0] out_22_36;
  output [7:0] out_22_37;
  output [7:0] out_22_38;
  output [7:0] out_22_39;
  output [7:0] out_22_40;
  output [7:0] out_22_41;
  output [7:0] out_22_42;
  output [7:0] out_22_43;
  output [7:0] out_22_44;
  output [7:0] out_22_45;
  output [7:0] out_22_46;
  output [7:0] out_22_47;
  output [7:0] out_22_48;
  output [7:0] out_22_49;
  output [7:0] out_22_50;
  output [7:0] out_22_51;
  output [7:0] out_22_52;
  output [7:0] out_22_53;
  output [7:0] out_22_54;
  output [7:0] out_22_55;
  output [7:0] out_22_56;
  output [7:0] out_22_57;
  output [7:0] out_22_58;
  output [7:0] out_22_59;
  output [7:0] out_22_60;
  output [7:0] out_22_61;
  output [7:0] out_22_62;
  output [7:0] out_22_63;
  output [7:0] out_22_64;
  output [7:0] out_23_1;
  output [7:0] out_23_2;
  output [7:0] out_23_3;
  output [7:0] out_23_4;
  output [7:0] out_23_5;
  output [7:0] out_23_6;
  output [7:0] out_23_7;
  output [7:0] out_23_8;
  output [7:0] out_23_9;
  output [7:0] out_23_10;
  output [7:0] out_23_11;
  output [7:0] out_23_12;
  output [7:0] out_23_13;
  output [7:0] out_23_14;
  output [7:0] out_23_15;
  output [7:0] out_23_16;
  output [7:0] out_23_17;
  output [7:0] out_23_18;
  output [7:0] out_23_19;
  output [7:0] out_23_20;
  output [7:0] out_23_21;
  output [7:0] out_23_22;
  output [7:0] out_23_23;
  output [7:0] out_23_24;
  output [7:0] out_23_25;
  output [7:0] out_23_26;
  output [7:0] out_23_27;
  output [7:0] out_23_28;
  output [7:0] out_23_29;
  output [7:0] out_23_30;
  output [7:0] out_23_31;
  output [7:0] out_23_32;
  output [7:0] out_23_33;
  output [7:0] out_23_34;
  output [7:0] out_23_35;
  output [7:0] out_23_36;
  output [7:0] out_23_37;
  output [7:0] out_23_38;
  output [7:0] out_23_39;
  output [7:0] out_23_40;
  output [7:0] out_23_41;
  output [7:0] out_23_42;
  output [7:0] out_23_43;
  output [7:0] out_23_44;
  output [7:0] out_23_45;
  output [7:0] out_23_46;
  output [7:0] out_23_47;
  output [7:0] out_23_48;
  output [7:0] out_23_49;
  output [7:0] out_23_50;
  output [7:0] out_23_51;
  output [7:0] out_23_52;
  output [7:0] out_23_53;
  output [7:0] out_23_54;
  output [7:0] out_23_55;
  output [7:0] out_23_56;
  output [7:0] out_23_57;
  output [7:0] out_23_58;
  output [7:0] out_23_59;
  output [7:0] out_23_60;
  output [7:0] out_23_61;
  output [7:0] out_23_62;
  output [7:0] out_23_63;
  output [7:0] out_23_64;
  output [7:0] out_24_1;
  output [7:0] out_24_2;
  output [7:0] out_24_3;
  output [7:0] out_24_4;
  output [7:0] out_24_5;
  output [7:0] out_24_6;
  output [7:0] out_24_7;
  output [7:0] out_24_8;
  output [7:0] out_24_9;
  output [7:0] out_24_10;
  output [7:0] out_24_11;
  output [7:0] out_24_12;
  output [7:0] out_24_13;
  output [7:0] out_24_14;
  output [7:0] out_24_15;
  output [7:0] out_24_16;
  output [7:0] out_24_17;
  output [7:0] out_24_18;
  output [7:0] out_24_19;
  output [7:0] out_24_20;
  output [7:0] out_24_21;
  output [7:0] out_24_22;
  output [7:0] out_24_23;
  output [7:0] out_24_24;
  output [7:0] out_24_25;
  output [7:0] out_24_26;
  output [7:0] out_24_27;
  output [7:0] out_24_28;
  output [7:0] out_24_29;
  output [7:0] out_24_30;
  output [7:0] out_24_31;
  output [7:0] out_24_32;
  output [7:0] out_24_33;
  output [7:0] out_24_34;
  output [7:0] out_24_35;
  output [7:0] out_24_36;
  output [7:0] out_24_37;
  output [7:0] out_24_38;
  output [7:0] out_24_39;
  output [7:0] out_24_40;
  output [7:0] out_24_41;
  output [7:0] out_24_42;
  output [7:0] out_24_43;
  output [7:0] out_24_44;
  output [7:0] out_24_45;
  output [7:0] out_24_46;
  output [7:0] out_24_47;
  output [7:0] out_24_48;
  output [7:0] out_24_49;
  output [7:0] out_24_50;
  output [7:0] out_24_51;
  output [7:0] out_24_52;
  output [7:0] out_24_53;
  output [7:0] out_24_54;
  output [7:0] out_24_55;
  output [7:0] out_24_56;
  output [7:0] out_24_57;
  output [7:0] out_24_58;
  output [7:0] out_24_59;
  output [7:0] out_24_60;
  output [7:0] out_24_61;
  output [7:0] out_24_62;
  output [7:0] out_24_63;
  output [7:0] out_24_64;
  output [7:0] out_25_1;
  output [7:0] out_25_2;
  output [7:0] out_25_3;
  output [7:0] out_25_4;
  output [7:0] out_25_5;
  output [7:0] out_25_6;
  output [7:0] out_25_7;
  output [7:0] out_25_8;
  output [7:0] out_25_9;
  output [7:0] out_25_10;
  output [7:0] out_25_11;
  output [7:0] out_25_12;
  output [7:0] out_25_13;
  output [7:0] out_25_14;
  output [7:0] out_25_15;
  output [7:0] out_25_16;
  output [7:0] out_25_17;
  output [7:0] out_25_18;
  output [7:0] out_25_19;
  output [7:0] out_25_20;
  output [7:0] out_25_21;
  output [7:0] out_25_22;
  output [7:0] out_25_23;
  output [7:0] out_25_24;
  output [7:0] out_25_25;
  output [7:0] out_25_26;
  output [7:0] out_25_27;
  output [7:0] out_25_28;
  output [7:0] out_25_29;
  output [7:0] out_25_30;
  output [7:0] out_25_31;
  output [7:0] out_25_32;
  output [7:0] out_25_33;
  output [7:0] out_25_34;
  output [7:0] out_25_35;
  output [7:0] out_25_36;
  output [7:0] out_25_37;
  output [7:0] out_25_38;
  output [7:0] out_25_39;
  output [7:0] out_25_40;
  output [7:0] out_25_41;
  output [7:0] out_25_42;
  output [7:0] out_25_43;
  output [7:0] out_25_44;
  output [7:0] out_25_45;
  output [7:0] out_25_46;
  output [7:0] out_25_47;
  output [7:0] out_25_48;
  output [7:0] out_25_49;
  output [7:0] out_25_50;
  output [7:0] out_25_51;
  output [7:0] out_25_52;
  output [7:0] out_25_53;
  output [7:0] out_25_54;
  output [7:0] out_25_55;
  output [7:0] out_25_56;
  output [7:0] out_25_57;
  output [7:0] out_25_58;
  output [7:0] out_25_59;
  output [7:0] out_25_60;
  output [7:0] out_25_61;
  output [7:0] out_25_62;
  output [7:0] out_25_63;
  output [7:0] out_25_64;
  output [7:0] out_26_1;
  output [7:0] out_26_2;
  output [7:0] out_26_3;
  output [7:0] out_26_4;
  output [7:0] out_26_5;
  output [7:0] out_26_6;
  output [7:0] out_26_7;
  output [7:0] out_26_8;
  output [7:0] out_26_9;
  output [7:0] out_26_10;
  output [7:0] out_26_11;
  output [7:0] out_26_12;
  output [7:0] out_26_13;
  output [7:0] out_26_14;
  output [7:0] out_26_15;
  output [7:0] out_26_16;
  output [7:0] out_26_17;
  output [7:0] out_26_18;
  output [7:0] out_26_19;
  output [7:0] out_26_20;
  output [7:0] out_26_21;
  output [7:0] out_26_22;
  output [7:0] out_26_23;
  output [7:0] out_26_24;
  output [7:0] out_26_25;
  output [7:0] out_26_26;
  output [7:0] out_26_27;
  output [7:0] out_26_28;
  output [7:0] out_26_29;
  output [7:0] out_26_30;
  output [7:0] out_26_31;
  output [7:0] out_26_32;
  output [7:0] out_26_33;
  output [7:0] out_26_34;
  output [7:0] out_26_35;
  output [7:0] out_26_36;
  output [7:0] out_26_37;
  output [7:0] out_26_38;
  output [7:0] out_26_39;
  output [7:0] out_26_40;
  output [7:0] out_26_41;
  output [7:0] out_26_42;
  output [7:0] out_26_43;
  output [7:0] out_26_44;
  output [7:0] out_26_45;
  output [7:0] out_26_46;
  output [7:0] out_26_47;
  output [7:0] out_26_48;
  output [7:0] out_26_49;
  output [7:0] out_26_50;
  output [7:0] out_26_51;
  output [7:0] out_26_52;
  output [7:0] out_26_53;
  output [7:0] out_26_54;
  output [7:0] out_26_55;
  output [7:0] out_26_56;
  output [7:0] out_26_57;
  output [7:0] out_26_58;
  output [7:0] out_26_59;
  output [7:0] out_26_60;
  output [7:0] out_26_61;
  output [7:0] out_26_62;
  output [7:0] out_26_63;
  output [7:0] out_26_64;
  output [7:0] out_27_1;
  output [7:0] out_27_2;
  output [7:0] out_27_3;
  output [7:0] out_27_4;
  output [7:0] out_27_5;
  output [7:0] out_27_6;
  output [7:0] out_27_7;
  output [7:0] out_27_8;
  output [7:0] out_27_9;
  output [7:0] out_27_10;
  output [7:0] out_27_11;
  output [7:0] out_27_12;
  output [7:0] out_27_13;
  output [7:0] out_27_14;
  output [7:0] out_27_15;
  output [7:0] out_27_16;
  output [7:0] out_27_17;
  output [7:0] out_27_18;
  output [7:0] out_27_19;
  output [7:0] out_27_20;
  output [7:0] out_27_21;
  output [7:0] out_27_22;
  output [7:0] out_27_23;
  output [7:0] out_27_24;
  output [7:0] out_27_25;
  output [7:0] out_27_26;
  output [7:0] out_27_27;
  output [7:0] out_27_28;
  output [7:0] out_27_29;
  output [7:0] out_27_30;
  output [7:0] out_27_31;
  output [7:0] out_27_32;
  output [7:0] out_27_33;
  output [7:0] out_27_34;
  output [7:0] out_27_35;
  output [7:0] out_27_36;
  output [7:0] out_27_37;
  output [7:0] out_27_38;
  output [7:0] out_27_39;
  output [7:0] out_27_40;
  output [7:0] out_27_41;
  output [7:0] out_27_42;
  output [7:0] out_27_43;
  output [7:0] out_27_44;
  output [7:0] out_27_45;
  output [7:0] out_27_46;
  output [7:0] out_27_47;
  output [7:0] out_27_48;
  output [7:0] out_27_49;
  output [7:0] out_27_50;
  output [7:0] out_27_51;
  output [7:0] out_27_52;
  output [7:0] out_27_53;
  output [7:0] out_27_54;
  output [7:0] out_27_55;
  output [7:0] out_27_56;
  output [7:0] out_27_57;
  output [7:0] out_27_58;
  output [7:0] out_27_59;
  output [7:0] out_27_60;
  output [7:0] out_27_61;
  output [7:0] out_27_62;
  output [7:0] out_27_63;
  output [7:0] out_27_64;
  output [7:0] out_28_1;
  output [7:0] out_28_2;
  output [7:0] out_28_3;
  output [7:0] out_28_4;
  output [7:0] out_28_5;
  output [7:0] out_28_6;
  output [7:0] out_28_7;
  output [7:0] out_28_8;
  output [7:0] out_28_9;
  output [7:0] out_28_10;
  output [7:0] out_28_11;
  output [7:0] out_28_12;
  output [7:0] out_28_13;
  output [7:0] out_28_14;
  output [7:0] out_28_15;
  output [7:0] out_28_16;
  output [7:0] out_28_17;
  output [7:0] out_28_18;
  output [7:0] out_28_19;
  output [7:0] out_28_20;
  output [7:0] out_28_21;
  output [7:0] out_28_22;
  output [7:0] out_28_23;
  output [7:0] out_28_24;
  output [7:0] out_28_25;
  output [7:0] out_28_26;
  output [7:0] out_28_27;
  output [7:0] out_28_28;
  output [7:0] out_28_29;
  output [7:0] out_28_30;
  output [7:0] out_28_31;
  output [7:0] out_28_32;
  output [7:0] out_28_33;
  output [7:0] out_28_34;
  output [7:0] out_28_35;
  output [7:0] out_28_36;
  output [7:0] out_28_37;
  output [7:0] out_28_38;
  output [7:0] out_28_39;
  output [7:0] out_28_40;
  output [7:0] out_28_41;
  output [7:0] out_28_42;
  output [7:0] out_28_43;
  output [7:0] out_28_44;
  output [7:0] out_28_45;
  output [7:0] out_28_46;
  output [7:0] out_28_47;
  output [7:0] out_28_48;
  output [7:0] out_28_49;
  output [7:0] out_28_50;
  output [7:0] out_28_51;
  output [7:0] out_28_52;
  output [7:0] out_28_53;
  output [7:0] out_28_54;
  output [7:0] out_28_55;
  output [7:0] out_28_56;
  output [7:0] out_28_57;
  output [7:0] out_28_58;
  output [7:0] out_28_59;
  output [7:0] out_28_60;
  output [7:0] out_28_61;
  output [7:0] out_28_62;
  output [7:0] out_28_63;
  output [7:0] out_28_64;
  output [7:0] out_29_1;
  output [7:0] out_29_2;
  output [7:0] out_29_3;
  output [7:0] out_29_4;
  output [7:0] out_29_5;
  output [7:0] out_29_6;
  output [7:0] out_29_7;
  output [7:0] out_29_8;
  output [7:0] out_29_9;
  output [7:0] out_29_10;
  output [7:0] out_29_11;
  output [7:0] out_29_12;
  output [7:0] out_29_13;
  output [7:0] out_29_14;
  output [7:0] out_29_15;
  output [7:0] out_29_16;
  output [7:0] out_29_17;
  output [7:0] out_29_18;
  output [7:0] out_29_19;
  output [7:0] out_29_20;
  output [7:0] out_29_21;
  output [7:0] out_29_22;
  output [7:0] out_29_23;
  output [7:0] out_29_24;
  output [7:0] out_29_25;
  output [7:0] out_29_26;
  output [7:0] out_29_27;
  output [7:0] out_29_28;
  output [7:0] out_29_29;
  output [7:0] out_29_30;
  output [7:0] out_29_31;
  output [7:0] out_29_32;
  output [7:0] out_29_33;
  output [7:0] out_29_34;
  output [7:0] out_29_35;
  output [7:0] out_29_36;
  output [7:0] out_29_37;
  output [7:0] out_29_38;
  output [7:0] out_29_39;
  output [7:0] out_29_40;
  output [7:0] out_29_41;
  output [7:0] out_29_42;
  output [7:0] out_29_43;
  output [7:0] out_29_44;
  output [7:0] out_29_45;
  output [7:0] out_29_46;
  output [7:0] out_29_47;
  output [7:0] out_29_48;
  output [7:0] out_29_49;
  output [7:0] out_29_50;
  output [7:0] out_29_51;
  output [7:0] out_29_52;
  output [7:0] out_29_53;
  output [7:0] out_29_54;
  output [7:0] out_29_55;
  output [7:0] out_29_56;
  output [7:0] out_29_57;
  output [7:0] out_29_58;
  output [7:0] out_29_59;
  output [7:0] out_29_60;
  output [7:0] out_29_61;
  output [7:0] out_29_62;
  output [7:0] out_29_63;
  output [7:0] out_29_64;
  output [7:0] out_30_1;
  output [7:0] out_30_2;
  output [7:0] out_30_3;
  output [7:0] out_30_4;
  output [7:0] out_30_5;
  output [7:0] out_30_6;
  output [7:0] out_30_7;
  output [7:0] out_30_8;
  output [7:0] out_30_9;
  output [7:0] out_30_10;
  output [7:0] out_30_11;
  output [7:0] out_30_12;
  output [7:0] out_30_13;
  output [7:0] out_30_14;
  output [7:0] out_30_15;
  output [7:0] out_30_16;
  output [7:0] out_30_17;
  output [7:0] out_30_18;
  output [7:0] out_30_19;
  output [7:0] out_30_20;
  output [7:0] out_30_21;
  output [7:0] out_30_22;
  output [7:0] out_30_23;
  output [7:0] out_30_24;
  output [7:0] out_30_25;
  output [7:0] out_30_26;
  output [7:0] out_30_27;
  output [7:0] out_30_28;
  output [7:0] out_30_29;
  output [7:0] out_30_30;
  output [7:0] out_30_31;
  output [7:0] out_30_32;
  output [7:0] out_30_33;
  output [7:0] out_30_34;
  output [7:0] out_30_35;
  output [7:0] out_30_36;
  output [7:0] out_30_37;
  output [7:0] out_30_38;
  output [7:0] out_30_39;
  output [7:0] out_30_40;
  output [7:0] out_30_41;
  output [7:0] out_30_42;
  output [7:0] out_30_43;
  output [7:0] out_30_44;
  output [7:0] out_30_45;
  output [7:0] out_30_46;
  output [7:0] out_30_47;
  output [7:0] out_30_48;
  output [7:0] out_30_49;
  output [7:0] out_30_50;
  output [7:0] out_30_51;
  output [7:0] out_30_52;
  output [7:0] out_30_53;
  output [7:0] out_30_54;
  output [7:0] out_30_55;
  output [7:0] out_30_56;
  output [7:0] out_30_57;
  output [7:0] out_30_58;
  output [7:0] out_30_59;
  output [7:0] out_30_60;
  output [7:0] out_30_61;
  output [7:0] out_30_62;
  output [7:0] out_30_63;
  output [7:0] out_30_64;
  output [7:0] out_31_1;
  output [7:0] out_31_2;
  output [7:0] out_31_3;
  output [7:0] out_31_4;
  output [7:0] out_31_5;
  output [7:0] out_31_6;
  output [7:0] out_31_7;
  output [7:0] out_31_8;
  output [7:0] out_31_9;
  output [7:0] out_31_10;
  output [7:0] out_31_11;
  output [7:0] out_31_12;
  output [7:0] out_31_13;
  output [7:0] out_31_14;
  output [7:0] out_31_15;
  output [7:0] out_31_16;
  output [7:0] out_31_17;
  output [7:0] out_31_18;
  output [7:0] out_31_19;
  output [7:0] out_31_20;
  output [7:0] out_31_21;
  output [7:0] out_31_22;
  output [7:0] out_31_23;
  output [7:0] out_31_24;
  output [7:0] out_31_25;
  output [7:0] out_31_26;
  output [7:0] out_31_27;
  output [7:0] out_31_28;
  output [7:0] out_31_29;
  output [7:0] out_31_30;
  output [7:0] out_31_31;
  output [7:0] out_31_32;
  output [7:0] out_31_33;
  output [7:0] out_31_34;
  output [7:0] out_31_35;
  output [7:0] out_31_36;
  output [7:0] out_31_37;
  output [7:0] out_31_38;
  output [7:0] out_31_39;
  output [7:0] out_31_40;
  output [7:0] out_31_41;
  output [7:0] out_31_42;
  output [7:0] out_31_43;
  output [7:0] out_31_44;
  output [7:0] out_31_45;
  output [7:0] out_31_46;
  output [7:0] out_31_47;
  output [7:0] out_31_48;
  output [7:0] out_31_49;
  output [7:0] out_31_50;
  output [7:0] out_31_51;
  output [7:0] out_31_52;
  output [7:0] out_31_53;
  output [7:0] out_31_54;
  output [7:0] out_31_55;
  output [7:0] out_31_56;
  output [7:0] out_31_57;
  output [7:0] out_31_58;
  output [7:0] out_31_59;
  output [7:0] out_31_60;
  output [7:0] out_31_61;
  output [7:0] out_31_62;
  output [7:0] out_31_63;
  output [7:0] out_31_64;
  output [7:0] out_32_1;
  output [7:0] out_32_2;
  output [7:0] out_32_3;
  output [7:0] out_32_4;
  output [7:0] out_32_5;
  output [7:0] out_32_6;
  output [7:0] out_32_7;
  output [7:0] out_32_8;
  output [7:0] out_32_9;
  output [7:0] out_32_10;
  output [7:0] out_32_11;
  output [7:0] out_32_12;
  output [7:0] out_32_13;
  output [7:0] out_32_14;
  output [7:0] out_32_15;
  output [7:0] out_32_16;
  output [7:0] out_32_17;
  output [7:0] out_32_18;
  output [7:0] out_32_19;
  output [7:0] out_32_20;
  output [7:0] out_32_21;
  output [7:0] out_32_22;
  output [7:0] out_32_23;
  output [7:0] out_32_24;
  output [7:0] out_32_25;
  output [7:0] out_32_26;
  output [7:0] out_32_27;
  output [7:0] out_32_28;
  output [7:0] out_32_29;
  output [7:0] out_32_30;
  output [7:0] out_32_31;
  output [7:0] out_32_32;
  output [7:0] out_32_33;
  output [7:0] out_32_34;
  output [7:0] out_32_35;
  output [7:0] out_32_36;
  output [7:0] out_32_37;
  output [7:0] out_32_38;
  output [7:0] out_32_39;
  output [7:0] out_32_40;
  output [7:0] out_32_41;
  output [7:0] out_32_42;
  output [7:0] out_32_43;
  output [7:0] out_32_44;
  output [7:0] out_32_45;
  output [7:0] out_32_46;
  output [7:0] out_32_47;
  output [7:0] out_32_48;
  output [7:0] out_32_49;
  output [7:0] out_32_50;
  output [7:0] out_32_51;
  output [7:0] out_32_52;
  output [7:0] out_32_53;
  output [7:0] out_32_54;
  output [7:0] out_32_55;
  output [7:0] out_32_56;
  output [7:0] out_32_57;
  output [7:0] out_32_58;
  output [7:0] out_32_59;
  output [7:0] out_32_60;
  output [7:0] out_32_61;
  output [7:0] out_32_62;
  output [7:0] out_32_63;
  output [7:0] out_32_64;
  output [7:0] out_33_1;
  output [7:0] out_33_2;
  output [7:0] out_33_3;
  output [7:0] out_33_4;
  output [7:0] out_33_5;
  output [7:0] out_33_6;
  output [7:0] out_33_7;
  output [7:0] out_33_8;
  output [7:0] out_33_9;
  output [7:0] out_33_10;
  output [7:0] out_33_11;
  output [7:0] out_33_12;
  output [7:0] out_33_13;
  output [7:0] out_33_14;
  output [7:0] out_33_15;
  output [7:0] out_33_16;
  output [7:0] out_33_17;
  output [7:0] out_33_18;
  output [7:0] out_33_19;
  output [7:0] out_33_20;
  output [7:0] out_33_21;
  output [7:0] out_33_22;
  output [7:0] out_33_23;
  output [7:0] out_33_24;
  output [7:0] out_33_25;
  output [7:0] out_33_26;
  output [7:0] out_33_27;
  output [7:0] out_33_28;
  output [7:0] out_33_29;
  output [7:0] out_33_30;
  output [7:0] out_33_31;
  output [7:0] out_33_32;
  output [7:0] out_33_33;
  output [7:0] out_33_34;
  output [7:0] out_33_35;
  output [7:0] out_33_36;
  output [7:0] out_33_37;
  output [7:0] out_33_38;
  output [7:0] out_33_39;
  output [7:0] out_33_40;
  output [7:0] out_33_41;
  output [7:0] out_33_42;
  output [7:0] out_33_43;
  output [7:0] out_33_44;
  output [7:0] out_33_45;
  output [7:0] out_33_46;
  output [7:0] out_33_47;
  output [7:0] out_33_48;
  output [7:0] out_33_49;
  output [7:0] out_33_50;
  output [7:0] out_33_51;
  output [7:0] out_33_52;
  output [7:0] out_33_53;
  output [7:0] out_33_54;
  output [7:0] out_33_55;
  output [7:0] out_33_56;
  output [7:0] out_33_57;
  output [7:0] out_33_58;
  output [7:0] out_33_59;
  output [7:0] out_33_60;
  output [7:0] out_33_61;
  output [7:0] out_33_62;
  output [7:0] out_33_63;
  output [7:0] out_33_64;
  output [7:0] out_34_1;
  output [7:0] out_34_2;
  output [7:0] out_34_3;
  output [7:0] out_34_4;
  output [7:0] out_34_5;
  output [7:0] out_34_6;
  output [7:0] out_34_7;
  output [7:0] out_34_8;
  output [7:0] out_34_9;
  output [7:0] out_34_10;
  output [7:0] out_34_11;
  output [7:0] out_34_12;
  output [7:0] out_34_13;
  output [7:0] out_34_14;
  output [7:0] out_34_15;
  output [7:0] out_34_16;
  output [7:0] out_34_17;
  output [7:0] out_34_18;
  output [7:0] out_34_19;
  output [7:0] out_34_20;
  output [7:0] out_34_21;
  output [7:0] out_34_22;
  output [7:0] out_34_23;
  output [7:0] out_34_24;
  output [7:0] out_34_25;
  output [7:0] out_34_26;
  output [7:0] out_34_27;
  output [7:0] out_34_28;
  output [7:0] out_34_29;
  output [7:0] out_34_30;
  output [7:0] out_34_31;
  output [7:0] out_34_32;
  output [7:0] out_34_33;
  output [7:0] out_34_34;
  output [7:0] out_34_35;
  output [7:0] out_34_36;
  output [7:0] out_34_37;
  output [7:0] out_34_38;
  output [7:0] out_34_39;
  output [7:0] out_34_40;
  output [7:0] out_34_41;
  output [7:0] out_34_42;
  output [7:0] out_34_43;
  output [7:0] out_34_44;
  output [7:0] out_34_45;
  output [7:0] out_34_46;
  output [7:0] out_34_47;
  output [7:0] out_34_48;
  output [7:0] out_34_49;
  output [7:0] out_34_50;
  output [7:0] out_34_51;
  output [7:0] out_34_52;
  output [7:0] out_34_53;
  output [7:0] out_34_54;
  output [7:0] out_34_55;
  output [7:0] out_34_56;
  output [7:0] out_34_57;
  output [7:0] out_34_58;
  output [7:0] out_34_59;
  output [7:0] out_34_60;
  output [7:0] out_34_61;
  output [7:0] out_34_62;
  output [7:0] out_34_63;
  output [7:0] out_34_64;
  output [7:0] out_35_1;
  output [7:0] out_35_2;
  output [7:0] out_35_3;
  output [7:0] out_35_4;
  output [7:0] out_35_5;
  output [7:0] out_35_6;
  output [7:0] out_35_7;
  output [7:0] out_35_8;
  output [7:0] out_35_9;
  output [7:0] out_35_10;
  output [7:0] out_35_11;
  output [7:0] out_35_12;
  output [7:0] out_35_13;
  output [7:0] out_35_14;
  output [7:0] out_35_15;
  output [7:0] out_35_16;
  output [7:0] out_35_17;
  output [7:0] out_35_18;
  output [7:0] out_35_19;
  output [7:0] out_35_20;
  output [7:0] out_35_21;
  output [7:0] out_35_22;
  output [7:0] out_35_23;
  output [7:0] out_35_24;
  output [7:0] out_35_25;
  output [7:0] out_35_26;
  output [7:0] out_35_27;
  output [7:0] out_35_28;
  output [7:0] out_35_29;
  output [7:0] out_35_30;
  output [7:0] out_35_31;
  output [7:0] out_35_32;
  output [7:0] out_35_33;
  output [7:0] out_35_34;
  output [7:0] out_35_35;
  output [7:0] out_35_36;
  output [7:0] out_35_37;
  output [7:0] out_35_38;
  output [7:0] out_35_39;
  output [7:0] out_35_40;
  output [7:0] out_35_41;
  output [7:0] out_35_42;
  output [7:0] out_35_43;
  output [7:0] out_35_44;
  output [7:0] out_35_45;
  output [7:0] out_35_46;
  output [7:0] out_35_47;
  output [7:0] out_35_48;
  output [7:0] out_35_49;
  output [7:0] out_35_50;
  output [7:0] out_35_51;
  output [7:0] out_35_52;
  output [7:0] out_35_53;
  output [7:0] out_35_54;
  output [7:0] out_35_55;
  output [7:0] out_35_56;
  output [7:0] out_35_57;
  output [7:0] out_35_58;
  output [7:0] out_35_59;
  output [7:0] out_35_60;
  output [7:0] out_35_61;
  output [7:0] out_35_62;
  output [7:0] out_35_63;
  output [7:0] out_35_64;
  output [7:0] out_36_1;
  output [7:0] out_36_2;
  output [7:0] out_36_3;
  output [7:0] out_36_4;
  output [7:0] out_36_5;
  output [7:0] out_36_6;
  output [7:0] out_36_7;
  output [7:0] out_36_8;
  output [7:0] out_36_9;
  output [7:0] out_36_10;
  output [7:0] out_36_11;
  output [7:0] out_36_12;
  output [7:0] out_36_13;
  output [7:0] out_36_14;
  output [7:0] out_36_15;
  output [7:0] out_36_16;
  output [7:0] out_36_17;
  output [7:0] out_36_18;
  output [7:0] out_36_19;
  output [7:0] out_36_20;
  output [7:0] out_36_21;
  output [7:0] out_36_22;
  output [7:0] out_36_23;
  output [7:0] out_36_24;
  output [7:0] out_36_25;
  output [7:0] out_36_26;
  output [7:0] out_36_27;
  output [7:0] out_36_28;
  output [7:0] out_36_29;
  output [7:0] out_36_30;
  output [7:0] out_36_31;
  output [7:0] out_36_32;
  output [7:0] out_36_33;
  output [7:0] out_36_34;
  output [7:0] out_36_35;
  output [7:0] out_36_36;
  output [7:0] out_36_37;
  output [7:0] out_36_38;
  output [7:0] out_36_39;
  output [7:0] out_36_40;
  output [7:0] out_36_41;
  output [7:0] out_36_42;
  output [7:0] out_36_43;
  output [7:0] out_36_44;
  output [7:0] out_36_45;
  output [7:0] out_36_46;
  output [7:0] out_36_47;
  output [7:0] out_36_48;
  output [7:0] out_36_49;
  output [7:0] out_36_50;
  output [7:0] out_36_51;
  output [7:0] out_36_52;
  output [7:0] out_36_53;
  output [7:0] out_36_54;
  output [7:0] out_36_55;
  output [7:0] out_36_56;
  output [7:0] out_36_57;
  output [7:0] out_36_58;
  output [7:0] out_36_59;
  output [7:0] out_36_60;
  output [7:0] out_36_61;
  output [7:0] out_36_62;
  output [7:0] out_36_63;
  output [7:0] out_36_64;
  output [7:0] out_37_1;
  output [7:0] out_37_2;
  output [7:0] out_37_3;
  output [7:0] out_37_4;
  output [7:0] out_37_5;
  output [7:0] out_37_6;
  output [7:0] out_37_7;
  output [7:0] out_37_8;
  output [7:0] out_37_9;
  output [7:0] out_37_10;
  output [7:0] out_37_11;
  output [7:0] out_37_12;
  output [7:0] out_37_13;
  output [7:0] out_37_14;
  output [7:0] out_37_15;
  output [7:0] out_37_16;
  output [7:0] out_37_17;
  output [7:0] out_37_18;
  output [7:0] out_37_19;
  output [7:0] out_37_20;
  output [7:0] out_37_21;
  output [7:0] out_37_22;
  output [7:0] out_37_23;
  output [7:0] out_37_24;
  output [7:0] out_37_25;
  output [7:0] out_37_26;
  output [7:0] out_37_27;
  output [7:0] out_37_28;
  output [7:0] out_37_29;
  output [7:0] out_37_30;
  output [7:0] out_37_31;
  output [7:0] out_37_32;
  output [7:0] out_37_33;
  output [7:0] out_37_34;
  output [7:0] out_37_35;
  output [7:0] out_37_36;
  output [7:0] out_37_37;
  output [7:0] out_37_38;
  output [7:0] out_37_39;
  output [7:0] out_37_40;
  output [7:0] out_37_41;
  output [7:0] out_37_42;
  output [7:0] out_37_43;
  output [7:0] out_37_44;
  output [7:0] out_37_45;
  output [7:0] out_37_46;
  output [7:0] out_37_47;
  output [7:0] out_37_48;
  output [7:0] out_37_49;
  output [7:0] out_37_50;
  output [7:0] out_37_51;
  output [7:0] out_37_52;
  output [7:0] out_37_53;
  output [7:0] out_37_54;
  output [7:0] out_37_55;
  output [7:0] out_37_56;
  output [7:0] out_37_57;
  output [7:0] out_37_58;
  output [7:0] out_37_59;
  output [7:0] out_37_60;
  output [7:0] out_37_61;
  output [7:0] out_37_62;
  output [7:0] out_37_63;
  output [7:0] out_37_64;
  output [7:0] out_38_1;
  output [7:0] out_38_2;
  output [7:0] out_38_3;
  output [7:0] out_38_4;
  output [7:0] out_38_5;
  output [7:0] out_38_6;
  output [7:0] out_38_7;
  output [7:0] out_38_8;
  output [7:0] out_38_9;
  output [7:0] out_38_10;
  output [7:0] out_38_11;
  output [7:0] out_38_12;
  output [7:0] out_38_13;
  output [7:0] out_38_14;
  output [7:0] out_38_15;
  output [7:0] out_38_16;
  output [7:0] out_38_17;
  output [7:0] out_38_18;
  output [7:0] out_38_19;
  output [7:0] out_38_20;
  output [7:0] out_38_21;
  output [7:0] out_38_22;
  output [7:0] out_38_23;
  output [7:0] out_38_24;
  output [7:0] out_38_25;
  output [7:0] out_38_26;
  output [7:0] out_38_27;
  output [7:0] out_38_28;
  output [7:0] out_38_29;
  output [7:0] out_38_30;
  output [7:0] out_38_31;
  output [7:0] out_38_32;
  output [7:0] out_38_33;
  output [7:0] out_38_34;
  output [7:0] out_38_35;
  output [7:0] out_38_36;
  output [7:0] out_38_37;
  output [7:0] out_38_38;
  output [7:0] out_38_39;
  output [7:0] out_38_40;
  output [7:0] out_38_41;
  output [7:0] out_38_42;
  output [7:0] out_38_43;
  output [7:0] out_38_44;
  output [7:0] out_38_45;
  output [7:0] out_38_46;
  output [7:0] out_38_47;
  output [7:0] out_38_48;
  output [7:0] out_38_49;
  output [7:0] out_38_50;
  output [7:0] out_38_51;
  output [7:0] out_38_52;
  output [7:0] out_38_53;
  output [7:0] out_38_54;
  output [7:0] out_38_55;
  output [7:0] out_38_56;
  output [7:0] out_38_57;
  output [7:0] out_38_58;
  output [7:0] out_38_59;
  output [7:0] out_38_60;
  output [7:0] out_38_61;
  output [7:0] out_38_62;
  output [7:0] out_38_63;
  output [7:0] out_38_64;
  output [7:0] out_39_1;
  output [7:0] out_39_2;
  output [7:0] out_39_3;
  output [7:0] out_39_4;
  output [7:0] out_39_5;
  output [7:0] out_39_6;
  output [7:0] out_39_7;
  output [7:0] out_39_8;
  output [7:0] out_39_9;
  output [7:0] out_39_10;
  output [7:0] out_39_11;
  output [7:0] out_39_12;
  output [7:0] out_39_13;
  output [7:0] out_39_14;
  output [7:0] out_39_15;
  output [7:0] out_39_16;
  output [7:0] out_39_17;
  output [7:0] out_39_18;
  output [7:0] out_39_19;
  output [7:0] out_39_20;
  output [7:0] out_39_21;
  output [7:0] out_39_22;
  output [7:0] out_39_23;
  output [7:0] out_39_24;
  output [7:0] out_39_25;
  output [7:0] out_39_26;
  output [7:0] out_39_27;
  output [7:0] out_39_28;
  output [7:0] out_39_29;
  output [7:0] out_39_30;
  output [7:0] out_39_31;
  output [7:0] out_39_32;
  output [7:0] out_39_33;
  output [7:0] out_39_34;
  output [7:0] out_39_35;
  output [7:0] out_39_36;
  output [7:0] out_39_37;
  output [7:0] out_39_38;
  output [7:0] out_39_39;
  output [7:0] out_39_40;
  output [7:0] out_39_41;
  output [7:0] out_39_42;
  output [7:0] out_39_43;
  output [7:0] out_39_44;
  output [7:0] out_39_45;
  output [7:0] out_39_46;
  output [7:0] out_39_47;
  output [7:0] out_39_48;
  output [7:0] out_39_49;
  output [7:0] out_39_50;
  output [7:0] out_39_51;
  output [7:0] out_39_52;
  output [7:0] out_39_53;
  output [7:0] out_39_54;
  output [7:0] out_39_55;
  output [7:0] out_39_56;
  output [7:0] out_39_57;
  output [7:0] out_39_58;
  output [7:0] out_39_59;
  output [7:0] out_39_60;
  output [7:0] out_39_61;
  output [7:0] out_39_62;
  output [7:0] out_39_63;
  output [7:0] out_39_64;
  output [7:0] out_40_1;
  output [7:0] out_40_2;
  output [7:0] out_40_3;
  output [7:0] out_40_4;
  output [7:0] out_40_5;
  output [7:0] out_40_6;
  output [7:0] out_40_7;
  output [7:0] out_40_8;
  output [7:0] out_40_9;
  output [7:0] out_40_10;
  output [7:0] out_40_11;
  output [7:0] out_40_12;
  output [7:0] out_40_13;
  output [7:0] out_40_14;
  output [7:0] out_40_15;
  output [7:0] out_40_16;
  output [7:0] out_40_17;
  output [7:0] out_40_18;
  output [7:0] out_40_19;
  output [7:0] out_40_20;
  output [7:0] out_40_21;
  output [7:0] out_40_22;
  output [7:0] out_40_23;
  output [7:0] out_40_24;
  output [7:0] out_40_25;
  output [7:0] out_40_26;
  output [7:0] out_40_27;
  output [7:0] out_40_28;
  output [7:0] out_40_29;
  output [7:0] out_40_30;
  output [7:0] out_40_31;
  output [7:0] out_40_32;
  output [7:0] out_40_33;
  output [7:0] out_40_34;
  output [7:0] out_40_35;
  output [7:0] out_40_36;
  output [7:0] out_40_37;
  output [7:0] out_40_38;
  output [7:0] out_40_39;
  output [7:0] out_40_40;
  output [7:0] out_40_41;
  output [7:0] out_40_42;
  output [7:0] out_40_43;
  output [7:0] out_40_44;
  output [7:0] out_40_45;
  output [7:0] out_40_46;
  output [7:0] out_40_47;
  output [7:0] out_40_48;
  output [7:0] out_40_49;
  output [7:0] out_40_50;
  output [7:0] out_40_51;
  output [7:0] out_40_52;
  output [7:0] out_40_53;
  output [7:0] out_40_54;
  output [7:0] out_40_55;
  output [7:0] out_40_56;
  output [7:0] out_40_57;
  output [7:0] out_40_58;
  output [7:0] out_40_59;
  output [7:0] out_40_60;
  output [7:0] out_40_61;
  output [7:0] out_40_62;
  output [7:0] out_40_63;
  output [7:0] out_40_64;
  output [7:0] out_41_1;
  output [7:0] out_41_2;
  output [7:0] out_41_3;
  output [7:0] out_41_4;
  output [7:0] out_41_5;
  output [7:0] out_41_6;
  output [7:0] out_41_7;
  output [7:0] out_41_8;
  output [7:0] out_41_9;
  output [7:0] out_41_10;
  output [7:0] out_41_11;
  output [7:0] out_41_12;
  output [7:0] out_41_13;
  output [7:0] out_41_14;
  output [7:0] out_41_15;
  output [7:0] out_41_16;
  output [7:0] out_41_17;
  output [7:0] out_41_18;
  output [7:0] out_41_19;
  output [7:0] out_41_20;
  output [7:0] out_41_21;
  output [7:0] out_41_22;
  output [7:0] out_41_23;
  output [7:0] out_41_24;
  output [7:0] out_41_25;
  output [7:0] out_41_26;
  output [7:0] out_41_27;
  output [7:0] out_41_28;
  output [7:0] out_41_29;
  output [7:0] out_41_30;
  output [7:0] out_41_31;
  output [7:0] out_41_32;
  output [7:0] out_41_33;
  output [7:0] out_41_34;
  output [7:0] out_41_35;
  output [7:0] out_41_36;
  output [7:0] out_41_37;
  output [7:0] out_41_38;
  output [7:0] out_41_39;
  output [7:0] out_41_40;
  output [7:0] out_41_41;
  output [7:0] out_41_42;
  output [7:0] out_41_43;
  output [7:0] out_41_44;
  output [7:0] out_41_45;
  output [7:0] out_41_46;
  output [7:0] out_41_47;
  output [7:0] out_41_48;
  output [7:0] out_41_49;
  output [7:0] out_41_50;
  output [7:0] out_41_51;
  output [7:0] out_41_52;
  output [7:0] out_41_53;
  output [7:0] out_41_54;
  output [7:0] out_41_55;
  output [7:0] out_41_56;
  output [7:0] out_41_57;
  output [7:0] out_41_58;
  output [7:0] out_41_59;
  output [7:0] out_41_60;
  output [7:0] out_41_61;
  output [7:0] out_41_62;
  output [7:0] out_41_63;
  output [7:0] out_41_64;
  output [7:0] out_42_1;
  output [7:0] out_42_2;
  output [7:0] out_42_3;
  output [7:0] out_42_4;
  output [7:0] out_42_5;
  output [7:0] out_42_6;
  output [7:0] out_42_7;
  output [7:0] out_42_8;
  output [7:0] out_42_9;
  output [7:0] out_42_10;
  output [7:0] out_42_11;
  output [7:0] out_42_12;
  output [7:0] out_42_13;
  output [7:0] out_42_14;
  output [7:0] out_42_15;
  output [7:0] out_42_16;
  output [7:0] out_42_17;
  output [7:0] out_42_18;
  output [7:0] out_42_19;
  output [7:0] out_42_20;
  output [7:0] out_42_21;
  output [7:0] out_42_22;
  output [7:0] out_42_23;
  output [7:0] out_42_24;
  output [7:0] out_42_25;
  output [7:0] out_42_26;
  output [7:0] out_42_27;
  output [7:0] out_42_28;
  output [7:0] out_42_29;
  output [7:0] out_42_30;
  output [7:0] out_42_31;
  output [7:0] out_42_32;
  output [7:0] out_42_33;
  output [7:0] out_42_34;
  output [7:0] out_42_35;
  output [7:0] out_42_36;
  output [7:0] out_42_37;
  output [7:0] out_42_38;
  output [7:0] out_42_39;
  output [7:0] out_42_40;
  output [7:0] out_42_41;
  output [7:0] out_42_42;
  output [7:0] out_42_43;
  output [7:0] out_42_44;
  output [7:0] out_42_45;
  output [7:0] out_42_46;
  output [7:0] out_42_47;
  output [7:0] out_42_48;
  output [7:0] out_42_49;
  output [7:0] out_42_50;
  output [7:0] out_42_51;
  output [7:0] out_42_52;
  output [7:0] out_42_53;
  output [7:0] out_42_54;
  output [7:0] out_42_55;
  output [7:0] out_42_56;
  output [7:0] out_42_57;
  output [7:0] out_42_58;
  output [7:0] out_42_59;
  output [7:0] out_42_60;
  output [7:0] out_42_61;
  output [7:0] out_42_62;
  output [7:0] out_42_63;
  output [7:0] out_42_64;
  output [7:0] out_43_1;
  output [7:0] out_43_2;
  output [7:0] out_43_3;
  output [7:0] out_43_4;
  output [7:0] out_43_5;
  output [7:0] out_43_6;
  output [7:0] out_43_7;
  output [7:0] out_43_8;
  output [7:0] out_43_9;
  output [7:0] out_43_10;
  output [7:0] out_43_11;
  output [7:0] out_43_12;
  output [7:0] out_43_13;
  output [7:0] out_43_14;
  output [7:0] out_43_15;
  output [7:0] out_43_16;
  output [7:0] out_43_17;
  output [7:0] out_43_18;
  output [7:0] out_43_19;
  output [7:0] out_43_20;
  output [7:0] out_43_21;
  output [7:0] out_43_22;
  output [7:0] out_43_23;
  output [7:0] out_43_24;
  output [7:0] out_43_25;
  output [7:0] out_43_26;
  output [7:0] out_43_27;
  output [7:0] out_43_28;
  output [7:0] out_43_29;
  output [7:0] out_43_30;
  output [7:0] out_43_31;
  output [7:0] out_43_32;
  output [7:0] out_43_33;
  output [7:0] out_43_34;
  output [7:0] out_43_35;
  output [7:0] out_43_36;
  output [7:0] out_43_37;
  output [7:0] out_43_38;
  output [7:0] out_43_39;
  output [7:0] out_43_40;
  output [7:0] out_43_41;
  output [7:0] out_43_42;
  output [7:0] out_43_43;
  output [7:0] out_43_44;
  output [7:0] out_43_45;
  output [7:0] out_43_46;
  output [7:0] out_43_47;
  output [7:0] out_43_48;
  output [7:0] out_43_49;
  output [7:0] out_43_50;
  output [7:0] out_43_51;
  output [7:0] out_43_52;
  output [7:0] out_43_53;
  output [7:0] out_43_54;
  output [7:0] out_43_55;
  output [7:0] out_43_56;
  output [7:0] out_43_57;
  output [7:0] out_43_58;
  output [7:0] out_43_59;
  output [7:0] out_43_60;
  output [7:0] out_43_61;
  output [7:0] out_43_62;
  output [7:0] out_43_63;
  output [7:0] out_43_64;

  wire [7:0] t_r0_c0_0;
  wire [7:0] t_r0_c0_1;
  wire [7:0] t_r0_c0_2;
  wire [7:0] t_r0_c0_3;
  wire [7:0] t_r0_c0_4;
  wire [7:0] t_r0_c0_5;
  wire [7:0] t_r0_c0_6;
  wire [7:0] t_r0_c0_7;
  wire [7:0] t_r0_c0_8;
  wire [7:0] t_r0_c0_9;
  wire [7:0] t_r0_c0_10;
  wire [7:0] t_r0_c0_11;
  wire [7:0] t_r0_c0_12;
  wire [7:0] t_r0_c1_0;
  wire [7:0] t_r0_c1_1;
  wire [7:0] t_r0_c1_2;
  wire [7:0] t_r0_c1_3;
  wire [7:0] t_r0_c1_4;
  wire [7:0] t_r0_c1_5;
  wire [7:0] t_r0_c1_6;
  wire [7:0] t_r0_c1_7;
  wire [7:0] t_r0_c1_8;
  wire [7:0] t_r0_c1_9;
  wire [7:0] t_r0_c1_10;
  wire [7:0] t_r0_c1_11;
  wire [7:0] t_r0_c1_12;
  wire [7:0] t_r0_c2_0;
  wire [7:0] t_r0_c2_1;
  wire [7:0] t_r0_c2_2;
  wire [7:0] t_r0_c2_3;
  wire [7:0] t_r0_c2_4;
  wire [7:0] t_r0_c2_5;
  wire [7:0] t_r0_c2_6;
  wire [7:0] t_r0_c2_7;
  wire [7:0] t_r0_c2_8;
  wire [7:0] t_r0_c2_9;
  wire [7:0] t_r0_c2_10;
  wire [7:0] t_r0_c2_11;
  wire [7:0] t_r0_c2_12;
  wire [7:0] t_r0_c3_0;
  wire [7:0] t_r0_c3_1;
  wire [7:0] t_r0_c3_2;
  wire [7:0] t_r0_c3_3;
  wire [7:0] t_r0_c3_4;
  wire [7:0] t_r0_c3_5;
  wire [7:0] t_r0_c3_6;
  wire [7:0] t_r0_c3_7;
  wire [7:0] t_r0_c3_8;
  wire [7:0] t_r0_c3_9;
  wire [7:0] t_r0_c3_10;
  wire [7:0] t_r0_c3_11;
  wire [7:0] t_r0_c3_12;
  wire [7:0] t_r0_c4_0;
  wire [7:0] t_r0_c4_1;
  wire [7:0] t_r0_c4_2;
  wire [7:0] t_r0_c4_3;
  wire [7:0] t_r0_c4_4;
  wire [7:0] t_r0_c4_5;
  wire [7:0] t_r0_c4_6;
  wire [7:0] t_r0_c4_7;
  wire [7:0] t_r0_c4_8;
  wire [7:0] t_r0_c4_9;
  wire [7:0] t_r0_c4_10;
  wire [7:0] t_r0_c4_11;
  wire [7:0] t_r0_c4_12;
  wire [7:0] t_r0_c5_0;
  wire [7:0] t_r0_c5_1;
  wire [7:0] t_r0_c5_2;
  wire [7:0] t_r0_c5_3;
  wire [7:0] t_r0_c5_4;
  wire [7:0] t_r0_c5_5;
  wire [7:0] t_r0_c5_6;
  wire [7:0] t_r0_c5_7;
  wire [7:0] t_r0_c5_8;
  wire [7:0] t_r0_c5_9;
  wire [7:0] t_r0_c5_10;
  wire [7:0] t_r0_c5_11;
  wire [7:0] t_r0_c5_12;
  wire [7:0] t_r0_c6_0;
  wire [7:0] t_r0_c6_1;
  wire [7:0] t_r0_c6_2;
  wire [7:0] t_r0_c6_3;
  wire [7:0] t_r0_c6_4;
  wire [7:0] t_r0_c6_5;
  wire [7:0] t_r0_c6_6;
  wire [7:0] t_r0_c6_7;
  wire [7:0] t_r0_c6_8;
  wire [7:0] t_r0_c6_9;
  wire [7:0] t_r0_c6_10;
  wire [7:0] t_r0_c6_11;
  wire [7:0] t_r0_c6_12;
  wire [7:0] t_r0_c7_0;
  wire [7:0] t_r0_c7_1;
  wire [7:0] t_r0_c7_2;
  wire [7:0] t_r0_c7_3;
  wire [7:0] t_r0_c7_4;
  wire [7:0] t_r0_c7_5;
  wire [7:0] t_r0_c7_6;
  wire [7:0] t_r0_c7_7;
  wire [7:0] t_r0_c7_8;
  wire [7:0] t_r0_c7_9;
  wire [7:0] t_r0_c7_10;
  wire [7:0] t_r0_c7_11;
  wire [7:0] t_r0_c7_12;
  wire [7:0] t_r0_c8_0;
  wire [7:0] t_r0_c8_1;
  wire [7:0] t_r0_c8_2;
  wire [7:0] t_r0_c8_3;
  wire [7:0] t_r0_c8_4;
  wire [7:0] t_r0_c8_5;
  wire [7:0] t_r0_c8_6;
  wire [7:0] t_r0_c8_7;
  wire [7:0] t_r0_c8_8;
  wire [7:0] t_r0_c8_9;
  wire [7:0] t_r0_c8_10;
  wire [7:0] t_r0_c8_11;
  wire [7:0] t_r0_c8_12;
  wire [7:0] t_r0_c9_0;
  wire [7:0] t_r0_c9_1;
  wire [7:0] t_r0_c9_2;
  wire [7:0] t_r0_c9_3;
  wire [7:0] t_r0_c9_4;
  wire [7:0] t_r0_c9_5;
  wire [7:0] t_r0_c9_6;
  wire [7:0] t_r0_c9_7;
  wire [7:0] t_r0_c9_8;
  wire [7:0] t_r0_c9_9;
  wire [7:0] t_r0_c9_10;
  wire [7:0] t_r0_c9_11;
  wire [7:0] t_r0_c9_12;
  wire [7:0] t_r0_c10_0;
  wire [7:0] t_r0_c10_1;
  wire [7:0] t_r0_c10_2;
  wire [7:0] t_r0_c10_3;
  wire [7:0] t_r0_c10_4;
  wire [7:0] t_r0_c10_5;
  wire [7:0] t_r0_c10_6;
  wire [7:0] t_r0_c10_7;
  wire [7:0] t_r0_c10_8;
  wire [7:0] t_r0_c10_9;
  wire [7:0] t_r0_c10_10;
  wire [7:0] t_r0_c10_11;
  wire [7:0] t_r0_c10_12;
  wire [7:0] t_r0_c11_0;
  wire [7:0] t_r0_c11_1;
  wire [7:0] t_r0_c11_2;
  wire [7:0] t_r0_c11_3;
  wire [7:0] t_r0_c11_4;
  wire [7:0] t_r0_c11_5;
  wire [7:0] t_r0_c11_6;
  wire [7:0] t_r0_c11_7;
  wire [7:0] t_r0_c11_8;
  wire [7:0] t_r0_c11_9;
  wire [7:0] t_r0_c11_10;
  wire [7:0] t_r0_c11_11;
  wire [7:0] t_r0_c11_12;
  wire [7:0] t_r0_c12_0;
  wire [7:0] t_r0_c12_1;
  wire [7:0] t_r0_c12_2;
  wire [7:0] t_r0_c12_3;
  wire [7:0] t_r0_c12_4;
  wire [7:0] t_r0_c12_5;
  wire [7:0] t_r0_c12_6;
  wire [7:0] t_r0_c12_7;
  wire [7:0] t_r0_c12_8;
  wire [7:0] t_r0_c12_9;
  wire [7:0] t_r0_c12_10;
  wire [7:0] t_r0_c12_11;
  wire [7:0] t_r0_c12_12;
  wire [7:0] t_r0_c13_0;
  wire [7:0] t_r0_c13_1;
  wire [7:0] t_r0_c13_2;
  wire [7:0] t_r0_c13_3;
  wire [7:0] t_r0_c13_4;
  wire [7:0] t_r0_c13_5;
  wire [7:0] t_r0_c13_6;
  wire [7:0] t_r0_c13_7;
  wire [7:0] t_r0_c13_8;
  wire [7:0] t_r0_c13_9;
  wire [7:0] t_r0_c13_10;
  wire [7:0] t_r0_c13_11;
  wire [7:0] t_r0_c13_12;
  wire [7:0] t_r0_c14_0;
  wire [7:0] t_r0_c14_1;
  wire [7:0] t_r0_c14_2;
  wire [7:0] t_r0_c14_3;
  wire [7:0] t_r0_c14_4;
  wire [7:0] t_r0_c14_5;
  wire [7:0] t_r0_c14_6;
  wire [7:0] t_r0_c14_7;
  wire [7:0] t_r0_c14_8;
  wire [7:0] t_r0_c14_9;
  wire [7:0] t_r0_c14_10;
  wire [7:0] t_r0_c14_11;
  wire [7:0] t_r0_c14_12;
  wire [7:0] t_r0_c15_0;
  wire [7:0] t_r0_c15_1;
  wire [7:0] t_r0_c15_2;
  wire [7:0] t_r0_c15_3;
  wire [7:0] t_r0_c15_4;
  wire [7:0] t_r0_c15_5;
  wire [7:0] t_r0_c15_6;
  wire [7:0] t_r0_c15_7;
  wire [7:0] t_r0_c15_8;
  wire [7:0] t_r0_c15_9;
  wire [7:0] t_r0_c15_10;
  wire [7:0] t_r0_c15_11;
  wire [7:0] t_r0_c15_12;
  wire [7:0] t_r0_c16_0;
  wire [7:0] t_r0_c16_1;
  wire [7:0] t_r0_c16_2;
  wire [7:0] t_r0_c16_3;
  wire [7:0] t_r0_c16_4;
  wire [7:0] t_r0_c16_5;
  wire [7:0] t_r0_c16_6;
  wire [7:0] t_r0_c16_7;
  wire [7:0] t_r0_c16_8;
  wire [7:0] t_r0_c16_9;
  wire [7:0] t_r0_c16_10;
  wire [7:0] t_r0_c16_11;
  wire [7:0] t_r0_c16_12;
  wire [7:0] t_r0_c17_0;
  wire [7:0] t_r0_c17_1;
  wire [7:0] t_r0_c17_2;
  wire [7:0] t_r0_c17_3;
  wire [7:0] t_r0_c17_4;
  wire [7:0] t_r0_c17_5;
  wire [7:0] t_r0_c17_6;
  wire [7:0] t_r0_c17_7;
  wire [7:0] t_r0_c17_8;
  wire [7:0] t_r0_c17_9;
  wire [7:0] t_r0_c17_10;
  wire [7:0] t_r0_c17_11;
  wire [7:0] t_r0_c17_12;
  wire [7:0] t_r0_c18_0;
  wire [7:0] t_r0_c18_1;
  wire [7:0] t_r0_c18_2;
  wire [7:0] t_r0_c18_3;
  wire [7:0] t_r0_c18_4;
  wire [7:0] t_r0_c18_5;
  wire [7:0] t_r0_c18_6;
  wire [7:0] t_r0_c18_7;
  wire [7:0] t_r0_c18_8;
  wire [7:0] t_r0_c18_9;
  wire [7:0] t_r0_c18_10;
  wire [7:0] t_r0_c18_11;
  wire [7:0] t_r0_c18_12;
  wire [7:0] t_r0_c19_0;
  wire [7:0] t_r0_c19_1;
  wire [7:0] t_r0_c19_2;
  wire [7:0] t_r0_c19_3;
  wire [7:0] t_r0_c19_4;
  wire [7:0] t_r0_c19_5;
  wire [7:0] t_r0_c19_6;
  wire [7:0] t_r0_c19_7;
  wire [7:0] t_r0_c19_8;
  wire [7:0] t_r0_c19_9;
  wire [7:0] t_r0_c19_10;
  wire [7:0] t_r0_c19_11;
  wire [7:0] t_r0_c19_12;
  wire [7:0] t_r0_c20_0;
  wire [7:0] t_r0_c20_1;
  wire [7:0] t_r0_c20_2;
  wire [7:0] t_r0_c20_3;
  wire [7:0] t_r0_c20_4;
  wire [7:0] t_r0_c20_5;
  wire [7:0] t_r0_c20_6;
  wire [7:0] t_r0_c20_7;
  wire [7:0] t_r0_c20_8;
  wire [7:0] t_r0_c20_9;
  wire [7:0] t_r0_c20_10;
  wire [7:0] t_r0_c20_11;
  wire [7:0] t_r0_c20_12;
  wire [7:0] t_r0_c21_0;
  wire [7:0] t_r0_c21_1;
  wire [7:0] t_r0_c21_2;
  wire [7:0] t_r0_c21_3;
  wire [7:0] t_r0_c21_4;
  wire [7:0] t_r0_c21_5;
  wire [7:0] t_r0_c21_6;
  wire [7:0] t_r0_c21_7;
  wire [7:0] t_r0_c21_8;
  wire [7:0] t_r0_c21_9;
  wire [7:0] t_r0_c21_10;
  wire [7:0] t_r0_c21_11;
  wire [7:0] t_r0_c21_12;
  wire [7:0] t_r0_c22_0;
  wire [7:0] t_r0_c22_1;
  wire [7:0] t_r0_c22_2;
  wire [7:0] t_r0_c22_3;
  wire [7:0] t_r0_c22_4;
  wire [7:0] t_r0_c22_5;
  wire [7:0] t_r0_c22_6;
  wire [7:0] t_r0_c22_7;
  wire [7:0] t_r0_c22_8;
  wire [7:0] t_r0_c22_9;
  wire [7:0] t_r0_c22_10;
  wire [7:0] t_r0_c22_11;
  wire [7:0] t_r0_c22_12;
  wire [7:0] t_r0_c23_0;
  wire [7:0] t_r0_c23_1;
  wire [7:0] t_r0_c23_2;
  wire [7:0] t_r0_c23_3;
  wire [7:0] t_r0_c23_4;
  wire [7:0] t_r0_c23_5;
  wire [7:0] t_r0_c23_6;
  wire [7:0] t_r0_c23_7;
  wire [7:0] t_r0_c23_8;
  wire [7:0] t_r0_c23_9;
  wire [7:0] t_r0_c23_10;
  wire [7:0] t_r0_c23_11;
  wire [7:0] t_r0_c23_12;
  wire [7:0] t_r0_c24_0;
  wire [7:0] t_r0_c24_1;
  wire [7:0] t_r0_c24_2;
  wire [7:0] t_r0_c24_3;
  wire [7:0] t_r0_c24_4;
  wire [7:0] t_r0_c24_5;
  wire [7:0] t_r0_c24_6;
  wire [7:0] t_r0_c24_7;
  wire [7:0] t_r0_c24_8;
  wire [7:0] t_r0_c24_9;
  wire [7:0] t_r0_c24_10;
  wire [7:0] t_r0_c24_11;
  wire [7:0] t_r0_c24_12;
  wire [7:0] t_r0_c25_0;
  wire [7:0] t_r0_c25_1;
  wire [7:0] t_r0_c25_2;
  wire [7:0] t_r0_c25_3;
  wire [7:0] t_r0_c25_4;
  wire [7:0] t_r0_c25_5;
  wire [7:0] t_r0_c25_6;
  wire [7:0] t_r0_c25_7;
  wire [7:0] t_r0_c25_8;
  wire [7:0] t_r0_c25_9;
  wire [7:0] t_r0_c25_10;
  wire [7:0] t_r0_c25_11;
  wire [7:0] t_r0_c25_12;
  wire [7:0] t_r0_c26_0;
  wire [7:0] t_r0_c26_1;
  wire [7:0] t_r0_c26_2;
  wire [7:0] t_r0_c26_3;
  wire [7:0] t_r0_c26_4;
  wire [7:0] t_r0_c26_5;
  wire [7:0] t_r0_c26_6;
  wire [7:0] t_r0_c26_7;
  wire [7:0] t_r0_c26_8;
  wire [7:0] t_r0_c26_9;
  wire [7:0] t_r0_c26_10;
  wire [7:0] t_r0_c26_11;
  wire [7:0] t_r0_c26_12;
  wire [7:0] t_r0_c27_0;
  wire [7:0] t_r0_c27_1;
  wire [7:0] t_r0_c27_2;
  wire [7:0] t_r0_c27_3;
  wire [7:0] t_r0_c27_4;
  wire [7:0] t_r0_c27_5;
  wire [7:0] t_r0_c27_6;
  wire [7:0] t_r0_c27_7;
  wire [7:0] t_r0_c27_8;
  wire [7:0] t_r0_c27_9;
  wire [7:0] t_r0_c27_10;
  wire [7:0] t_r0_c27_11;
  wire [7:0] t_r0_c27_12;
  wire [7:0] t_r0_c28_0;
  wire [7:0] t_r0_c28_1;
  wire [7:0] t_r0_c28_2;
  wire [7:0] t_r0_c28_3;
  wire [7:0] t_r0_c28_4;
  wire [7:0] t_r0_c28_5;
  wire [7:0] t_r0_c28_6;
  wire [7:0] t_r0_c28_7;
  wire [7:0] t_r0_c28_8;
  wire [7:0] t_r0_c28_9;
  wire [7:0] t_r0_c28_10;
  wire [7:0] t_r0_c28_11;
  wire [7:0] t_r0_c28_12;
  wire [7:0] t_r0_c29_0;
  wire [7:0] t_r0_c29_1;
  wire [7:0] t_r0_c29_2;
  wire [7:0] t_r0_c29_3;
  wire [7:0] t_r0_c29_4;
  wire [7:0] t_r0_c29_5;
  wire [7:0] t_r0_c29_6;
  wire [7:0] t_r0_c29_7;
  wire [7:0] t_r0_c29_8;
  wire [7:0] t_r0_c29_9;
  wire [7:0] t_r0_c29_10;
  wire [7:0] t_r0_c29_11;
  wire [7:0] t_r0_c29_12;
  wire [7:0] t_r0_c30_0;
  wire [7:0] t_r0_c30_1;
  wire [7:0] t_r0_c30_2;
  wire [7:0] t_r0_c30_3;
  wire [7:0] t_r0_c30_4;
  wire [7:0] t_r0_c30_5;
  wire [7:0] t_r0_c30_6;
  wire [7:0] t_r0_c30_7;
  wire [7:0] t_r0_c30_8;
  wire [7:0] t_r0_c30_9;
  wire [7:0] t_r0_c30_10;
  wire [7:0] t_r0_c30_11;
  wire [7:0] t_r0_c30_12;
  wire [7:0] t_r0_c31_0;
  wire [7:0] t_r0_c31_1;
  wire [7:0] t_r0_c31_2;
  wire [7:0] t_r0_c31_3;
  wire [7:0] t_r0_c31_4;
  wire [7:0] t_r0_c31_5;
  wire [7:0] t_r0_c31_6;
  wire [7:0] t_r0_c31_7;
  wire [7:0] t_r0_c31_8;
  wire [7:0] t_r0_c31_9;
  wire [7:0] t_r0_c31_10;
  wire [7:0] t_r0_c31_11;
  wire [7:0] t_r0_c31_12;
  wire [7:0] t_r0_c32_0;
  wire [7:0] t_r0_c32_1;
  wire [7:0] t_r0_c32_2;
  wire [7:0] t_r0_c32_3;
  wire [7:0] t_r0_c32_4;
  wire [7:0] t_r0_c32_5;
  wire [7:0] t_r0_c32_6;
  wire [7:0] t_r0_c32_7;
  wire [7:0] t_r0_c32_8;
  wire [7:0] t_r0_c32_9;
  wire [7:0] t_r0_c32_10;
  wire [7:0] t_r0_c32_11;
  wire [7:0] t_r0_c32_12;
  wire [7:0] t_r0_c33_0;
  wire [7:0] t_r0_c33_1;
  wire [7:0] t_r0_c33_2;
  wire [7:0] t_r0_c33_3;
  wire [7:0] t_r0_c33_4;
  wire [7:0] t_r0_c33_5;
  wire [7:0] t_r0_c33_6;
  wire [7:0] t_r0_c33_7;
  wire [7:0] t_r0_c33_8;
  wire [7:0] t_r0_c33_9;
  wire [7:0] t_r0_c33_10;
  wire [7:0] t_r0_c33_11;
  wire [7:0] t_r0_c33_12;
  wire [7:0] t_r0_c34_0;
  wire [7:0] t_r0_c34_1;
  wire [7:0] t_r0_c34_2;
  wire [7:0] t_r0_c34_3;
  wire [7:0] t_r0_c34_4;
  wire [7:0] t_r0_c34_5;
  wire [7:0] t_r0_c34_6;
  wire [7:0] t_r0_c34_7;
  wire [7:0] t_r0_c34_8;
  wire [7:0] t_r0_c34_9;
  wire [7:0] t_r0_c34_10;
  wire [7:0] t_r0_c34_11;
  wire [7:0] t_r0_c34_12;
  wire [7:0] t_r0_c35_0;
  wire [7:0] t_r0_c35_1;
  wire [7:0] t_r0_c35_2;
  wire [7:0] t_r0_c35_3;
  wire [7:0] t_r0_c35_4;
  wire [7:0] t_r0_c35_5;
  wire [7:0] t_r0_c35_6;
  wire [7:0] t_r0_c35_7;
  wire [7:0] t_r0_c35_8;
  wire [7:0] t_r0_c35_9;
  wire [7:0] t_r0_c35_10;
  wire [7:0] t_r0_c35_11;
  wire [7:0] t_r0_c35_12;
  wire [7:0] t_r0_c36_0;
  wire [7:0] t_r0_c36_1;
  wire [7:0] t_r0_c36_2;
  wire [7:0] t_r0_c36_3;
  wire [7:0] t_r0_c36_4;
  wire [7:0] t_r0_c36_5;
  wire [7:0] t_r0_c36_6;
  wire [7:0] t_r0_c36_7;
  wire [7:0] t_r0_c36_8;
  wire [7:0] t_r0_c36_9;
  wire [7:0] t_r0_c36_10;
  wire [7:0] t_r0_c36_11;
  wire [7:0] t_r0_c36_12;
  wire [7:0] t_r0_c37_0;
  wire [7:0] t_r0_c37_1;
  wire [7:0] t_r0_c37_2;
  wire [7:0] t_r0_c37_3;
  wire [7:0] t_r0_c37_4;
  wire [7:0] t_r0_c37_5;
  wire [7:0] t_r0_c37_6;
  wire [7:0] t_r0_c37_7;
  wire [7:0] t_r0_c37_8;
  wire [7:0] t_r0_c37_9;
  wire [7:0] t_r0_c37_10;
  wire [7:0] t_r0_c37_11;
  wire [7:0] t_r0_c37_12;
  wire [7:0] t_r0_c38_0;
  wire [7:0] t_r0_c38_1;
  wire [7:0] t_r0_c38_2;
  wire [7:0] t_r0_c38_3;
  wire [7:0] t_r0_c38_4;
  wire [7:0] t_r0_c38_5;
  wire [7:0] t_r0_c38_6;
  wire [7:0] t_r0_c38_7;
  wire [7:0] t_r0_c38_8;
  wire [7:0] t_r0_c38_9;
  wire [7:0] t_r0_c38_10;
  wire [7:0] t_r0_c38_11;
  wire [7:0] t_r0_c38_12;
  wire [7:0] t_r0_c39_0;
  wire [7:0] t_r0_c39_1;
  wire [7:0] t_r0_c39_2;
  wire [7:0] t_r0_c39_3;
  wire [7:0] t_r0_c39_4;
  wire [7:0] t_r0_c39_5;
  wire [7:0] t_r0_c39_6;
  wire [7:0] t_r0_c39_7;
  wire [7:0] t_r0_c39_8;
  wire [7:0] t_r0_c39_9;
  wire [7:0] t_r0_c39_10;
  wire [7:0] t_r0_c39_11;
  wire [7:0] t_r0_c39_12;
  wire [7:0] t_r0_c40_0;
  wire [7:0] t_r0_c40_1;
  wire [7:0] t_r0_c40_2;
  wire [7:0] t_r0_c40_3;
  wire [7:0] t_r0_c40_4;
  wire [7:0] t_r0_c40_5;
  wire [7:0] t_r0_c40_6;
  wire [7:0] t_r0_c40_7;
  wire [7:0] t_r0_c40_8;
  wire [7:0] t_r0_c40_9;
  wire [7:0] t_r0_c40_10;
  wire [7:0] t_r0_c40_11;
  wire [7:0] t_r0_c40_12;
  wire [7:0] t_r0_c41_0;
  wire [7:0] t_r0_c41_1;
  wire [7:0] t_r0_c41_2;
  wire [7:0] t_r0_c41_3;
  wire [7:0] t_r0_c41_4;
  wire [7:0] t_r0_c41_5;
  wire [7:0] t_r0_c41_6;
  wire [7:0] t_r0_c41_7;
  wire [7:0] t_r0_c41_8;
  wire [7:0] t_r0_c41_9;
  wire [7:0] t_r0_c41_10;
  wire [7:0] t_r0_c41_11;
  wire [7:0] t_r0_c41_12;
  wire [7:0] t_r0_c42_0;
  wire [7:0] t_r0_c42_1;
  wire [7:0] t_r0_c42_2;
  wire [7:0] t_r0_c42_3;
  wire [7:0] t_r0_c42_4;
  wire [7:0] t_r0_c42_5;
  wire [7:0] t_r0_c42_6;
  wire [7:0] t_r0_c42_7;
  wire [7:0] t_r0_c42_8;
  wire [7:0] t_r0_c42_9;
  wire [7:0] t_r0_c42_10;
  wire [7:0] t_r0_c42_11;
  wire [7:0] t_r0_c42_12;
  wire [7:0] t_r0_c43_0;
  wire [7:0] t_r0_c43_1;
  wire [7:0] t_r0_c43_2;
  wire [7:0] t_r0_c43_3;
  wire [7:0] t_r0_c43_4;
  wire [7:0] t_r0_c43_5;
  wire [7:0] t_r0_c43_6;
  wire [7:0] t_r0_c43_7;
  wire [7:0] t_r0_c43_8;
  wire [7:0] t_r0_c43_9;
  wire [7:0] t_r0_c43_10;
  wire [7:0] t_r0_c43_11;
  wire [7:0] t_r0_c43_12;
  wire [7:0] t_r0_c44_0;
  wire [7:0] t_r0_c44_1;
  wire [7:0] t_r0_c44_2;
  wire [7:0] t_r0_c44_3;
  wire [7:0] t_r0_c44_4;
  wire [7:0] t_r0_c44_5;
  wire [7:0] t_r0_c44_6;
  wire [7:0] t_r0_c44_7;
  wire [7:0] t_r0_c44_8;
  wire [7:0] t_r0_c44_9;
  wire [7:0] t_r0_c44_10;
  wire [7:0] t_r0_c44_11;
  wire [7:0] t_r0_c44_12;
  wire [7:0] t_r0_c45_0;
  wire [7:0] t_r0_c45_1;
  wire [7:0] t_r0_c45_2;
  wire [7:0] t_r0_c45_3;
  wire [7:0] t_r0_c45_4;
  wire [7:0] t_r0_c45_5;
  wire [7:0] t_r0_c45_6;
  wire [7:0] t_r0_c45_7;
  wire [7:0] t_r0_c45_8;
  wire [7:0] t_r0_c45_9;
  wire [7:0] t_r0_c45_10;
  wire [7:0] t_r0_c45_11;
  wire [7:0] t_r0_c45_12;
  wire [7:0] t_r0_c46_0;
  wire [7:0] t_r0_c46_1;
  wire [7:0] t_r0_c46_2;
  wire [7:0] t_r0_c46_3;
  wire [7:0] t_r0_c46_4;
  wire [7:0] t_r0_c46_5;
  wire [7:0] t_r0_c46_6;
  wire [7:0] t_r0_c46_7;
  wire [7:0] t_r0_c46_8;
  wire [7:0] t_r0_c46_9;
  wire [7:0] t_r0_c46_10;
  wire [7:0] t_r0_c46_11;
  wire [7:0] t_r0_c46_12;
  wire [7:0] t_r0_c47_0;
  wire [7:0] t_r0_c47_1;
  wire [7:0] t_r0_c47_2;
  wire [7:0] t_r0_c47_3;
  wire [7:0] t_r0_c47_4;
  wire [7:0] t_r0_c47_5;
  wire [7:0] t_r0_c47_6;
  wire [7:0] t_r0_c47_7;
  wire [7:0] t_r0_c47_8;
  wire [7:0] t_r0_c47_9;
  wire [7:0] t_r0_c47_10;
  wire [7:0] t_r0_c47_11;
  wire [7:0] t_r0_c47_12;
  wire [7:0] t_r0_c48_0;
  wire [7:0] t_r0_c48_1;
  wire [7:0] t_r0_c48_2;
  wire [7:0] t_r0_c48_3;
  wire [7:0] t_r0_c48_4;
  wire [7:0] t_r0_c48_5;
  wire [7:0] t_r0_c48_6;
  wire [7:0] t_r0_c48_7;
  wire [7:0] t_r0_c48_8;
  wire [7:0] t_r0_c48_9;
  wire [7:0] t_r0_c48_10;
  wire [7:0] t_r0_c48_11;
  wire [7:0] t_r0_c48_12;
  wire [7:0] t_r0_c49_0;
  wire [7:0] t_r0_c49_1;
  wire [7:0] t_r0_c49_2;
  wire [7:0] t_r0_c49_3;
  wire [7:0] t_r0_c49_4;
  wire [7:0] t_r0_c49_5;
  wire [7:0] t_r0_c49_6;
  wire [7:0] t_r0_c49_7;
  wire [7:0] t_r0_c49_8;
  wire [7:0] t_r0_c49_9;
  wire [7:0] t_r0_c49_10;
  wire [7:0] t_r0_c49_11;
  wire [7:0] t_r0_c49_12;
  wire [7:0] t_r0_c50_0;
  wire [7:0] t_r0_c50_1;
  wire [7:0] t_r0_c50_2;
  wire [7:0] t_r0_c50_3;
  wire [7:0] t_r0_c50_4;
  wire [7:0] t_r0_c50_5;
  wire [7:0] t_r0_c50_6;
  wire [7:0] t_r0_c50_7;
  wire [7:0] t_r0_c50_8;
  wire [7:0] t_r0_c50_9;
  wire [7:0] t_r0_c50_10;
  wire [7:0] t_r0_c50_11;
  wire [7:0] t_r0_c50_12;
  wire [7:0] t_r0_c51_0;
  wire [7:0] t_r0_c51_1;
  wire [7:0] t_r0_c51_2;
  wire [7:0] t_r0_c51_3;
  wire [7:0] t_r0_c51_4;
  wire [7:0] t_r0_c51_5;
  wire [7:0] t_r0_c51_6;
  wire [7:0] t_r0_c51_7;
  wire [7:0] t_r0_c51_8;
  wire [7:0] t_r0_c51_9;
  wire [7:0] t_r0_c51_10;
  wire [7:0] t_r0_c51_11;
  wire [7:0] t_r0_c51_12;
  wire [7:0] t_r0_c52_0;
  wire [7:0] t_r0_c52_1;
  wire [7:0] t_r0_c52_2;
  wire [7:0] t_r0_c52_3;
  wire [7:0] t_r0_c52_4;
  wire [7:0] t_r0_c52_5;
  wire [7:0] t_r0_c52_6;
  wire [7:0] t_r0_c52_7;
  wire [7:0] t_r0_c52_8;
  wire [7:0] t_r0_c52_9;
  wire [7:0] t_r0_c52_10;
  wire [7:0] t_r0_c52_11;
  wire [7:0] t_r0_c52_12;
  wire [7:0] t_r0_c53_0;
  wire [7:0] t_r0_c53_1;
  wire [7:0] t_r0_c53_2;
  wire [7:0] t_r0_c53_3;
  wire [7:0] t_r0_c53_4;
  wire [7:0] t_r0_c53_5;
  wire [7:0] t_r0_c53_6;
  wire [7:0] t_r0_c53_7;
  wire [7:0] t_r0_c53_8;
  wire [7:0] t_r0_c53_9;
  wire [7:0] t_r0_c53_10;
  wire [7:0] t_r0_c53_11;
  wire [7:0] t_r0_c53_12;
  wire [7:0] t_r0_c54_0;
  wire [7:0] t_r0_c54_1;
  wire [7:0] t_r0_c54_2;
  wire [7:0] t_r0_c54_3;
  wire [7:0] t_r0_c54_4;
  wire [7:0] t_r0_c54_5;
  wire [7:0] t_r0_c54_6;
  wire [7:0] t_r0_c54_7;
  wire [7:0] t_r0_c54_8;
  wire [7:0] t_r0_c54_9;
  wire [7:0] t_r0_c54_10;
  wire [7:0] t_r0_c54_11;
  wire [7:0] t_r0_c54_12;
  wire [7:0] t_r0_c55_0;
  wire [7:0] t_r0_c55_1;
  wire [7:0] t_r0_c55_2;
  wire [7:0] t_r0_c55_3;
  wire [7:0] t_r0_c55_4;
  wire [7:0] t_r0_c55_5;
  wire [7:0] t_r0_c55_6;
  wire [7:0] t_r0_c55_7;
  wire [7:0] t_r0_c55_8;
  wire [7:0] t_r0_c55_9;
  wire [7:0] t_r0_c55_10;
  wire [7:0] t_r0_c55_11;
  wire [7:0] t_r0_c55_12;
  wire [7:0] t_r0_c56_0;
  wire [7:0] t_r0_c56_1;
  wire [7:0] t_r0_c56_2;
  wire [7:0] t_r0_c56_3;
  wire [7:0] t_r0_c56_4;
  wire [7:0] t_r0_c56_5;
  wire [7:0] t_r0_c56_6;
  wire [7:0] t_r0_c56_7;
  wire [7:0] t_r0_c56_8;
  wire [7:0] t_r0_c56_9;
  wire [7:0] t_r0_c56_10;
  wire [7:0] t_r0_c56_11;
  wire [7:0] t_r0_c56_12;
  wire [7:0] t_r0_c57_0;
  wire [7:0] t_r0_c57_1;
  wire [7:0] t_r0_c57_2;
  wire [7:0] t_r0_c57_3;
  wire [7:0] t_r0_c57_4;
  wire [7:0] t_r0_c57_5;
  wire [7:0] t_r0_c57_6;
  wire [7:0] t_r0_c57_7;
  wire [7:0] t_r0_c57_8;
  wire [7:0] t_r0_c57_9;
  wire [7:0] t_r0_c57_10;
  wire [7:0] t_r0_c57_11;
  wire [7:0] t_r0_c57_12;
  wire [7:0] t_r0_c58_0;
  wire [7:0] t_r0_c58_1;
  wire [7:0] t_r0_c58_2;
  wire [7:0] t_r0_c58_3;
  wire [7:0] t_r0_c58_4;
  wire [7:0] t_r0_c58_5;
  wire [7:0] t_r0_c58_6;
  wire [7:0] t_r0_c58_7;
  wire [7:0] t_r0_c58_8;
  wire [7:0] t_r0_c58_9;
  wire [7:0] t_r0_c58_10;
  wire [7:0] t_r0_c58_11;
  wire [7:0] t_r0_c58_12;
  wire [7:0] t_r0_c59_0;
  wire [7:0] t_r0_c59_1;
  wire [7:0] t_r0_c59_2;
  wire [7:0] t_r0_c59_3;
  wire [7:0] t_r0_c59_4;
  wire [7:0] t_r0_c59_5;
  wire [7:0] t_r0_c59_6;
  wire [7:0] t_r0_c59_7;
  wire [7:0] t_r0_c59_8;
  wire [7:0] t_r0_c59_9;
  wire [7:0] t_r0_c59_10;
  wire [7:0] t_r0_c59_11;
  wire [7:0] t_r0_c59_12;
  wire [7:0] t_r0_c60_0;
  wire [7:0] t_r0_c60_1;
  wire [7:0] t_r0_c60_2;
  wire [7:0] t_r0_c60_3;
  wire [7:0] t_r0_c60_4;
  wire [7:0] t_r0_c60_5;
  wire [7:0] t_r0_c60_6;
  wire [7:0] t_r0_c60_7;
  wire [7:0] t_r0_c60_8;
  wire [7:0] t_r0_c60_9;
  wire [7:0] t_r0_c60_10;
  wire [7:0] t_r0_c60_11;
  wire [7:0] t_r0_c60_12;
  wire [7:0] t_r0_c61_0;
  wire [7:0] t_r0_c61_1;
  wire [7:0] t_r0_c61_2;
  wire [7:0] t_r0_c61_3;
  wire [7:0] t_r0_c61_4;
  wire [7:0] t_r0_c61_5;
  wire [7:0] t_r0_c61_6;
  wire [7:0] t_r0_c61_7;
  wire [7:0] t_r0_c61_8;
  wire [7:0] t_r0_c61_9;
  wire [7:0] t_r0_c61_10;
  wire [7:0] t_r0_c61_11;
  wire [7:0] t_r0_c61_12;
  wire [7:0] t_r0_c62_0;
  wire [7:0] t_r0_c62_1;
  wire [7:0] t_r0_c62_2;
  wire [7:0] t_r0_c62_3;
  wire [7:0] t_r0_c62_4;
  wire [7:0] t_r0_c62_5;
  wire [7:0] t_r0_c62_6;
  wire [7:0] t_r0_c62_7;
  wire [7:0] t_r0_c62_8;
  wire [7:0] t_r0_c62_9;
  wire [7:0] t_r0_c62_10;
  wire [7:0] t_r0_c62_11;
  wire [7:0] t_r0_c62_12;
  wire [7:0] t_r0_c63_0;
  wire [7:0] t_r0_c63_1;
  wire [7:0] t_r0_c63_2;
  wire [7:0] t_r0_c63_3;
  wire [7:0] t_r0_c63_4;
  wire [7:0] t_r0_c63_5;
  wire [7:0] t_r0_c63_6;
  wire [7:0] t_r0_c63_7;
  wire [7:0] t_r0_c63_8;
  wire [7:0] t_r0_c63_9;
  wire [7:0] t_r0_c63_10;
  wire [7:0] t_r0_c63_11;
  wire [7:0] t_r0_c63_12;
  wire [7:0] t_r0_c64_0;
  wire [7:0] t_r0_c64_1;
  wire [7:0] t_r0_c64_2;
  wire [7:0] t_r0_c64_3;
  wire [7:0] t_r0_c64_4;
  wire [7:0] t_r0_c64_5;
  wire [7:0] t_r0_c64_6;
  wire [7:0] t_r0_c64_7;
  wire [7:0] t_r0_c64_8;
  wire [7:0] t_r0_c64_9;
  wire [7:0] t_r0_c64_10;
  wire [7:0] t_r0_c64_11;
  wire [7:0] t_r0_c64_12;
  wire [7:0] t_r0_c65_0;
  wire [7:0] t_r0_c65_1;
  wire [7:0] t_r0_c65_2;
  wire [7:0] t_r0_c65_3;
  wire [7:0] t_r0_c65_4;
  wire [7:0] t_r0_c65_5;
  wire [7:0] t_r0_c65_6;
  wire [7:0] t_r0_c65_7;
  wire [7:0] t_r0_c65_8;
  wire [7:0] t_r0_c65_9;
  wire [7:0] t_r0_c65_10;
  wire [7:0] t_r0_c65_11;
  wire [7:0] t_r0_c65_12;
  wire [7:0] t_r1_c0_0;
  wire [7:0] t_r1_c0_1;
  wire [7:0] t_r1_c0_2;
  wire [7:0] t_r1_c0_3;
  wire [7:0] t_r1_c0_4;
  wire [7:0] t_r1_c0_5;
  wire [7:0] t_r1_c0_6;
  wire [7:0] t_r1_c0_7;
  wire [7:0] t_r1_c0_8;
  wire [7:0] t_r1_c0_9;
  wire [7:0] t_r1_c0_10;
  wire [7:0] t_r1_c0_11;
  wire [7:0] t_r1_c0_12;
  wire [7:0] t_r1_c1_0;
  wire [7:0] t_r1_c1_1;
  wire [7:0] t_r1_c1_2;
  wire [7:0] t_r1_c1_3;
  wire [7:0] t_r1_c1_4;
  wire [7:0] t_r1_c1_5;
  wire [7:0] t_r1_c1_6;
  wire [7:0] t_r1_c1_7;
  wire [7:0] t_r1_c1_8;
  wire [7:0] t_r1_c1_9;
  wire [7:0] t_r1_c1_10;
  wire [7:0] t_r1_c1_11;
  wire [7:0] t_r1_c1_12;
  wire [7:0] t_r1_c2_0;
  wire [7:0] t_r1_c2_1;
  wire [7:0] t_r1_c2_2;
  wire [7:0] t_r1_c2_3;
  wire [7:0] t_r1_c2_4;
  wire [7:0] t_r1_c2_5;
  wire [7:0] t_r1_c2_6;
  wire [7:0] t_r1_c2_7;
  wire [7:0] t_r1_c2_8;
  wire [7:0] t_r1_c2_9;
  wire [7:0] t_r1_c2_10;
  wire [7:0] t_r1_c2_11;
  wire [7:0] t_r1_c2_12;
  wire [7:0] t_r1_c3_0;
  wire [7:0] t_r1_c3_1;
  wire [7:0] t_r1_c3_2;
  wire [7:0] t_r1_c3_3;
  wire [7:0] t_r1_c3_4;
  wire [7:0] t_r1_c3_5;
  wire [7:0] t_r1_c3_6;
  wire [7:0] t_r1_c3_7;
  wire [7:0] t_r1_c3_8;
  wire [7:0] t_r1_c3_9;
  wire [7:0] t_r1_c3_10;
  wire [7:0] t_r1_c3_11;
  wire [7:0] t_r1_c3_12;
  wire [7:0] t_r1_c4_0;
  wire [7:0] t_r1_c4_1;
  wire [7:0] t_r1_c4_2;
  wire [7:0] t_r1_c4_3;
  wire [7:0] t_r1_c4_4;
  wire [7:0] t_r1_c4_5;
  wire [7:0] t_r1_c4_6;
  wire [7:0] t_r1_c4_7;
  wire [7:0] t_r1_c4_8;
  wire [7:0] t_r1_c4_9;
  wire [7:0] t_r1_c4_10;
  wire [7:0] t_r1_c4_11;
  wire [7:0] t_r1_c4_12;
  wire [7:0] t_r1_c5_0;
  wire [7:0] t_r1_c5_1;
  wire [7:0] t_r1_c5_2;
  wire [7:0] t_r1_c5_3;
  wire [7:0] t_r1_c5_4;
  wire [7:0] t_r1_c5_5;
  wire [7:0] t_r1_c5_6;
  wire [7:0] t_r1_c5_7;
  wire [7:0] t_r1_c5_8;
  wire [7:0] t_r1_c5_9;
  wire [7:0] t_r1_c5_10;
  wire [7:0] t_r1_c5_11;
  wire [7:0] t_r1_c5_12;
  wire [7:0] t_r1_c6_0;
  wire [7:0] t_r1_c6_1;
  wire [7:0] t_r1_c6_2;
  wire [7:0] t_r1_c6_3;
  wire [7:0] t_r1_c6_4;
  wire [7:0] t_r1_c6_5;
  wire [7:0] t_r1_c6_6;
  wire [7:0] t_r1_c6_7;
  wire [7:0] t_r1_c6_8;
  wire [7:0] t_r1_c6_9;
  wire [7:0] t_r1_c6_10;
  wire [7:0] t_r1_c6_11;
  wire [7:0] t_r1_c6_12;
  wire [7:0] t_r1_c7_0;
  wire [7:0] t_r1_c7_1;
  wire [7:0] t_r1_c7_2;
  wire [7:0] t_r1_c7_3;
  wire [7:0] t_r1_c7_4;
  wire [7:0] t_r1_c7_5;
  wire [7:0] t_r1_c7_6;
  wire [7:0] t_r1_c7_7;
  wire [7:0] t_r1_c7_8;
  wire [7:0] t_r1_c7_9;
  wire [7:0] t_r1_c7_10;
  wire [7:0] t_r1_c7_11;
  wire [7:0] t_r1_c7_12;
  wire [7:0] t_r1_c8_0;
  wire [7:0] t_r1_c8_1;
  wire [7:0] t_r1_c8_2;
  wire [7:0] t_r1_c8_3;
  wire [7:0] t_r1_c8_4;
  wire [7:0] t_r1_c8_5;
  wire [7:0] t_r1_c8_6;
  wire [7:0] t_r1_c8_7;
  wire [7:0] t_r1_c8_8;
  wire [7:0] t_r1_c8_9;
  wire [7:0] t_r1_c8_10;
  wire [7:0] t_r1_c8_11;
  wire [7:0] t_r1_c8_12;
  wire [7:0] t_r1_c9_0;
  wire [7:0] t_r1_c9_1;
  wire [7:0] t_r1_c9_2;
  wire [7:0] t_r1_c9_3;
  wire [7:0] t_r1_c9_4;
  wire [7:0] t_r1_c9_5;
  wire [7:0] t_r1_c9_6;
  wire [7:0] t_r1_c9_7;
  wire [7:0] t_r1_c9_8;
  wire [7:0] t_r1_c9_9;
  wire [7:0] t_r1_c9_10;
  wire [7:0] t_r1_c9_11;
  wire [7:0] t_r1_c9_12;
  wire [7:0] t_r1_c10_0;
  wire [7:0] t_r1_c10_1;
  wire [7:0] t_r1_c10_2;
  wire [7:0] t_r1_c10_3;
  wire [7:0] t_r1_c10_4;
  wire [7:0] t_r1_c10_5;
  wire [7:0] t_r1_c10_6;
  wire [7:0] t_r1_c10_7;
  wire [7:0] t_r1_c10_8;
  wire [7:0] t_r1_c10_9;
  wire [7:0] t_r1_c10_10;
  wire [7:0] t_r1_c10_11;
  wire [7:0] t_r1_c10_12;
  wire [7:0] t_r1_c11_0;
  wire [7:0] t_r1_c11_1;
  wire [7:0] t_r1_c11_2;
  wire [7:0] t_r1_c11_3;
  wire [7:0] t_r1_c11_4;
  wire [7:0] t_r1_c11_5;
  wire [7:0] t_r1_c11_6;
  wire [7:0] t_r1_c11_7;
  wire [7:0] t_r1_c11_8;
  wire [7:0] t_r1_c11_9;
  wire [7:0] t_r1_c11_10;
  wire [7:0] t_r1_c11_11;
  wire [7:0] t_r1_c11_12;
  wire [7:0] t_r1_c12_0;
  wire [7:0] t_r1_c12_1;
  wire [7:0] t_r1_c12_2;
  wire [7:0] t_r1_c12_3;
  wire [7:0] t_r1_c12_4;
  wire [7:0] t_r1_c12_5;
  wire [7:0] t_r1_c12_6;
  wire [7:0] t_r1_c12_7;
  wire [7:0] t_r1_c12_8;
  wire [7:0] t_r1_c12_9;
  wire [7:0] t_r1_c12_10;
  wire [7:0] t_r1_c12_11;
  wire [7:0] t_r1_c12_12;
  wire [7:0] t_r1_c13_0;
  wire [7:0] t_r1_c13_1;
  wire [7:0] t_r1_c13_2;
  wire [7:0] t_r1_c13_3;
  wire [7:0] t_r1_c13_4;
  wire [7:0] t_r1_c13_5;
  wire [7:0] t_r1_c13_6;
  wire [7:0] t_r1_c13_7;
  wire [7:0] t_r1_c13_8;
  wire [7:0] t_r1_c13_9;
  wire [7:0] t_r1_c13_10;
  wire [7:0] t_r1_c13_11;
  wire [7:0] t_r1_c13_12;
  wire [7:0] t_r1_c14_0;
  wire [7:0] t_r1_c14_1;
  wire [7:0] t_r1_c14_2;
  wire [7:0] t_r1_c14_3;
  wire [7:0] t_r1_c14_4;
  wire [7:0] t_r1_c14_5;
  wire [7:0] t_r1_c14_6;
  wire [7:0] t_r1_c14_7;
  wire [7:0] t_r1_c14_8;
  wire [7:0] t_r1_c14_9;
  wire [7:0] t_r1_c14_10;
  wire [7:0] t_r1_c14_11;
  wire [7:0] t_r1_c14_12;
  wire [7:0] t_r1_c15_0;
  wire [7:0] t_r1_c15_1;
  wire [7:0] t_r1_c15_2;
  wire [7:0] t_r1_c15_3;
  wire [7:0] t_r1_c15_4;
  wire [7:0] t_r1_c15_5;
  wire [7:0] t_r1_c15_6;
  wire [7:0] t_r1_c15_7;
  wire [7:0] t_r1_c15_8;
  wire [7:0] t_r1_c15_9;
  wire [7:0] t_r1_c15_10;
  wire [7:0] t_r1_c15_11;
  wire [7:0] t_r1_c15_12;
  wire [7:0] t_r1_c16_0;
  wire [7:0] t_r1_c16_1;
  wire [7:0] t_r1_c16_2;
  wire [7:0] t_r1_c16_3;
  wire [7:0] t_r1_c16_4;
  wire [7:0] t_r1_c16_5;
  wire [7:0] t_r1_c16_6;
  wire [7:0] t_r1_c16_7;
  wire [7:0] t_r1_c16_8;
  wire [7:0] t_r1_c16_9;
  wire [7:0] t_r1_c16_10;
  wire [7:0] t_r1_c16_11;
  wire [7:0] t_r1_c16_12;
  wire [7:0] t_r1_c17_0;
  wire [7:0] t_r1_c17_1;
  wire [7:0] t_r1_c17_2;
  wire [7:0] t_r1_c17_3;
  wire [7:0] t_r1_c17_4;
  wire [7:0] t_r1_c17_5;
  wire [7:0] t_r1_c17_6;
  wire [7:0] t_r1_c17_7;
  wire [7:0] t_r1_c17_8;
  wire [7:0] t_r1_c17_9;
  wire [7:0] t_r1_c17_10;
  wire [7:0] t_r1_c17_11;
  wire [7:0] t_r1_c17_12;
  wire [7:0] t_r1_c18_0;
  wire [7:0] t_r1_c18_1;
  wire [7:0] t_r1_c18_2;
  wire [7:0] t_r1_c18_3;
  wire [7:0] t_r1_c18_4;
  wire [7:0] t_r1_c18_5;
  wire [7:0] t_r1_c18_6;
  wire [7:0] t_r1_c18_7;
  wire [7:0] t_r1_c18_8;
  wire [7:0] t_r1_c18_9;
  wire [7:0] t_r1_c18_10;
  wire [7:0] t_r1_c18_11;
  wire [7:0] t_r1_c18_12;
  wire [7:0] t_r1_c19_0;
  wire [7:0] t_r1_c19_1;
  wire [7:0] t_r1_c19_2;
  wire [7:0] t_r1_c19_3;
  wire [7:0] t_r1_c19_4;
  wire [7:0] t_r1_c19_5;
  wire [7:0] t_r1_c19_6;
  wire [7:0] t_r1_c19_7;
  wire [7:0] t_r1_c19_8;
  wire [7:0] t_r1_c19_9;
  wire [7:0] t_r1_c19_10;
  wire [7:0] t_r1_c19_11;
  wire [7:0] t_r1_c19_12;
  wire [7:0] t_r1_c20_0;
  wire [7:0] t_r1_c20_1;
  wire [7:0] t_r1_c20_2;
  wire [7:0] t_r1_c20_3;
  wire [7:0] t_r1_c20_4;
  wire [7:0] t_r1_c20_5;
  wire [7:0] t_r1_c20_6;
  wire [7:0] t_r1_c20_7;
  wire [7:0] t_r1_c20_8;
  wire [7:0] t_r1_c20_9;
  wire [7:0] t_r1_c20_10;
  wire [7:0] t_r1_c20_11;
  wire [7:0] t_r1_c20_12;
  wire [7:0] t_r1_c21_0;
  wire [7:0] t_r1_c21_1;
  wire [7:0] t_r1_c21_2;
  wire [7:0] t_r1_c21_3;
  wire [7:0] t_r1_c21_4;
  wire [7:0] t_r1_c21_5;
  wire [7:0] t_r1_c21_6;
  wire [7:0] t_r1_c21_7;
  wire [7:0] t_r1_c21_8;
  wire [7:0] t_r1_c21_9;
  wire [7:0] t_r1_c21_10;
  wire [7:0] t_r1_c21_11;
  wire [7:0] t_r1_c21_12;
  wire [7:0] t_r1_c22_0;
  wire [7:0] t_r1_c22_1;
  wire [7:0] t_r1_c22_2;
  wire [7:0] t_r1_c22_3;
  wire [7:0] t_r1_c22_4;
  wire [7:0] t_r1_c22_5;
  wire [7:0] t_r1_c22_6;
  wire [7:0] t_r1_c22_7;
  wire [7:0] t_r1_c22_8;
  wire [7:0] t_r1_c22_9;
  wire [7:0] t_r1_c22_10;
  wire [7:0] t_r1_c22_11;
  wire [7:0] t_r1_c22_12;
  wire [7:0] t_r1_c23_0;
  wire [7:0] t_r1_c23_1;
  wire [7:0] t_r1_c23_2;
  wire [7:0] t_r1_c23_3;
  wire [7:0] t_r1_c23_4;
  wire [7:0] t_r1_c23_5;
  wire [7:0] t_r1_c23_6;
  wire [7:0] t_r1_c23_7;
  wire [7:0] t_r1_c23_8;
  wire [7:0] t_r1_c23_9;
  wire [7:0] t_r1_c23_10;
  wire [7:0] t_r1_c23_11;
  wire [7:0] t_r1_c23_12;
  wire [7:0] t_r1_c24_0;
  wire [7:0] t_r1_c24_1;
  wire [7:0] t_r1_c24_2;
  wire [7:0] t_r1_c24_3;
  wire [7:0] t_r1_c24_4;
  wire [7:0] t_r1_c24_5;
  wire [7:0] t_r1_c24_6;
  wire [7:0] t_r1_c24_7;
  wire [7:0] t_r1_c24_8;
  wire [7:0] t_r1_c24_9;
  wire [7:0] t_r1_c24_10;
  wire [7:0] t_r1_c24_11;
  wire [7:0] t_r1_c24_12;
  wire [7:0] t_r1_c25_0;
  wire [7:0] t_r1_c25_1;
  wire [7:0] t_r1_c25_2;
  wire [7:0] t_r1_c25_3;
  wire [7:0] t_r1_c25_4;
  wire [7:0] t_r1_c25_5;
  wire [7:0] t_r1_c25_6;
  wire [7:0] t_r1_c25_7;
  wire [7:0] t_r1_c25_8;
  wire [7:0] t_r1_c25_9;
  wire [7:0] t_r1_c25_10;
  wire [7:0] t_r1_c25_11;
  wire [7:0] t_r1_c25_12;
  wire [7:0] t_r1_c26_0;
  wire [7:0] t_r1_c26_1;
  wire [7:0] t_r1_c26_2;
  wire [7:0] t_r1_c26_3;
  wire [7:0] t_r1_c26_4;
  wire [7:0] t_r1_c26_5;
  wire [7:0] t_r1_c26_6;
  wire [7:0] t_r1_c26_7;
  wire [7:0] t_r1_c26_8;
  wire [7:0] t_r1_c26_9;
  wire [7:0] t_r1_c26_10;
  wire [7:0] t_r1_c26_11;
  wire [7:0] t_r1_c26_12;
  wire [7:0] t_r1_c27_0;
  wire [7:0] t_r1_c27_1;
  wire [7:0] t_r1_c27_2;
  wire [7:0] t_r1_c27_3;
  wire [7:0] t_r1_c27_4;
  wire [7:0] t_r1_c27_5;
  wire [7:0] t_r1_c27_6;
  wire [7:0] t_r1_c27_7;
  wire [7:0] t_r1_c27_8;
  wire [7:0] t_r1_c27_9;
  wire [7:0] t_r1_c27_10;
  wire [7:0] t_r1_c27_11;
  wire [7:0] t_r1_c27_12;
  wire [7:0] t_r1_c28_0;
  wire [7:0] t_r1_c28_1;
  wire [7:0] t_r1_c28_2;
  wire [7:0] t_r1_c28_3;
  wire [7:0] t_r1_c28_4;
  wire [7:0] t_r1_c28_5;
  wire [7:0] t_r1_c28_6;
  wire [7:0] t_r1_c28_7;
  wire [7:0] t_r1_c28_8;
  wire [7:0] t_r1_c28_9;
  wire [7:0] t_r1_c28_10;
  wire [7:0] t_r1_c28_11;
  wire [7:0] t_r1_c28_12;
  wire [7:0] t_r1_c29_0;
  wire [7:0] t_r1_c29_1;
  wire [7:0] t_r1_c29_2;
  wire [7:0] t_r1_c29_3;
  wire [7:0] t_r1_c29_4;
  wire [7:0] t_r1_c29_5;
  wire [7:0] t_r1_c29_6;
  wire [7:0] t_r1_c29_7;
  wire [7:0] t_r1_c29_8;
  wire [7:0] t_r1_c29_9;
  wire [7:0] t_r1_c29_10;
  wire [7:0] t_r1_c29_11;
  wire [7:0] t_r1_c29_12;
  wire [7:0] t_r1_c30_0;
  wire [7:0] t_r1_c30_1;
  wire [7:0] t_r1_c30_2;
  wire [7:0] t_r1_c30_3;
  wire [7:0] t_r1_c30_4;
  wire [7:0] t_r1_c30_5;
  wire [7:0] t_r1_c30_6;
  wire [7:0] t_r1_c30_7;
  wire [7:0] t_r1_c30_8;
  wire [7:0] t_r1_c30_9;
  wire [7:0] t_r1_c30_10;
  wire [7:0] t_r1_c30_11;
  wire [7:0] t_r1_c30_12;
  wire [7:0] t_r1_c31_0;
  wire [7:0] t_r1_c31_1;
  wire [7:0] t_r1_c31_2;
  wire [7:0] t_r1_c31_3;
  wire [7:0] t_r1_c31_4;
  wire [7:0] t_r1_c31_5;
  wire [7:0] t_r1_c31_6;
  wire [7:0] t_r1_c31_7;
  wire [7:0] t_r1_c31_8;
  wire [7:0] t_r1_c31_9;
  wire [7:0] t_r1_c31_10;
  wire [7:0] t_r1_c31_11;
  wire [7:0] t_r1_c31_12;
  wire [7:0] t_r1_c32_0;
  wire [7:0] t_r1_c32_1;
  wire [7:0] t_r1_c32_2;
  wire [7:0] t_r1_c32_3;
  wire [7:0] t_r1_c32_4;
  wire [7:0] t_r1_c32_5;
  wire [7:0] t_r1_c32_6;
  wire [7:0] t_r1_c32_7;
  wire [7:0] t_r1_c32_8;
  wire [7:0] t_r1_c32_9;
  wire [7:0] t_r1_c32_10;
  wire [7:0] t_r1_c32_11;
  wire [7:0] t_r1_c32_12;
  wire [7:0] t_r1_c33_0;
  wire [7:0] t_r1_c33_1;
  wire [7:0] t_r1_c33_2;
  wire [7:0] t_r1_c33_3;
  wire [7:0] t_r1_c33_4;
  wire [7:0] t_r1_c33_5;
  wire [7:0] t_r1_c33_6;
  wire [7:0] t_r1_c33_7;
  wire [7:0] t_r1_c33_8;
  wire [7:0] t_r1_c33_9;
  wire [7:0] t_r1_c33_10;
  wire [7:0] t_r1_c33_11;
  wire [7:0] t_r1_c33_12;
  wire [7:0] t_r1_c34_0;
  wire [7:0] t_r1_c34_1;
  wire [7:0] t_r1_c34_2;
  wire [7:0] t_r1_c34_3;
  wire [7:0] t_r1_c34_4;
  wire [7:0] t_r1_c34_5;
  wire [7:0] t_r1_c34_6;
  wire [7:0] t_r1_c34_7;
  wire [7:0] t_r1_c34_8;
  wire [7:0] t_r1_c34_9;
  wire [7:0] t_r1_c34_10;
  wire [7:0] t_r1_c34_11;
  wire [7:0] t_r1_c34_12;
  wire [7:0] t_r1_c35_0;
  wire [7:0] t_r1_c35_1;
  wire [7:0] t_r1_c35_2;
  wire [7:0] t_r1_c35_3;
  wire [7:0] t_r1_c35_4;
  wire [7:0] t_r1_c35_5;
  wire [7:0] t_r1_c35_6;
  wire [7:0] t_r1_c35_7;
  wire [7:0] t_r1_c35_8;
  wire [7:0] t_r1_c35_9;
  wire [7:0] t_r1_c35_10;
  wire [7:0] t_r1_c35_11;
  wire [7:0] t_r1_c35_12;
  wire [7:0] t_r1_c36_0;
  wire [7:0] t_r1_c36_1;
  wire [7:0] t_r1_c36_2;
  wire [7:0] t_r1_c36_3;
  wire [7:0] t_r1_c36_4;
  wire [7:0] t_r1_c36_5;
  wire [7:0] t_r1_c36_6;
  wire [7:0] t_r1_c36_7;
  wire [7:0] t_r1_c36_8;
  wire [7:0] t_r1_c36_9;
  wire [7:0] t_r1_c36_10;
  wire [7:0] t_r1_c36_11;
  wire [7:0] t_r1_c36_12;
  wire [7:0] t_r1_c37_0;
  wire [7:0] t_r1_c37_1;
  wire [7:0] t_r1_c37_2;
  wire [7:0] t_r1_c37_3;
  wire [7:0] t_r1_c37_4;
  wire [7:0] t_r1_c37_5;
  wire [7:0] t_r1_c37_6;
  wire [7:0] t_r1_c37_7;
  wire [7:0] t_r1_c37_8;
  wire [7:0] t_r1_c37_9;
  wire [7:0] t_r1_c37_10;
  wire [7:0] t_r1_c37_11;
  wire [7:0] t_r1_c37_12;
  wire [7:0] t_r1_c38_0;
  wire [7:0] t_r1_c38_1;
  wire [7:0] t_r1_c38_2;
  wire [7:0] t_r1_c38_3;
  wire [7:0] t_r1_c38_4;
  wire [7:0] t_r1_c38_5;
  wire [7:0] t_r1_c38_6;
  wire [7:0] t_r1_c38_7;
  wire [7:0] t_r1_c38_8;
  wire [7:0] t_r1_c38_9;
  wire [7:0] t_r1_c38_10;
  wire [7:0] t_r1_c38_11;
  wire [7:0] t_r1_c38_12;
  wire [7:0] t_r1_c39_0;
  wire [7:0] t_r1_c39_1;
  wire [7:0] t_r1_c39_2;
  wire [7:0] t_r1_c39_3;
  wire [7:0] t_r1_c39_4;
  wire [7:0] t_r1_c39_5;
  wire [7:0] t_r1_c39_6;
  wire [7:0] t_r1_c39_7;
  wire [7:0] t_r1_c39_8;
  wire [7:0] t_r1_c39_9;
  wire [7:0] t_r1_c39_10;
  wire [7:0] t_r1_c39_11;
  wire [7:0] t_r1_c39_12;
  wire [7:0] t_r1_c40_0;
  wire [7:0] t_r1_c40_1;
  wire [7:0] t_r1_c40_2;
  wire [7:0] t_r1_c40_3;
  wire [7:0] t_r1_c40_4;
  wire [7:0] t_r1_c40_5;
  wire [7:0] t_r1_c40_6;
  wire [7:0] t_r1_c40_7;
  wire [7:0] t_r1_c40_8;
  wire [7:0] t_r1_c40_9;
  wire [7:0] t_r1_c40_10;
  wire [7:0] t_r1_c40_11;
  wire [7:0] t_r1_c40_12;
  wire [7:0] t_r1_c41_0;
  wire [7:0] t_r1_c41_1;
  wire [7:0] t_r1_c41_2;
  wire [7:0] t_r1_c41_3;
  wire [7:0] t_r1_c41_4;
  wire [7:0] t_r1_c41_5;
  wire [7:0] t_r1_c41_6;
  wire [7:0] t_r1_c41_7;
  wire [7:0] t_r1_c41_8;
  wire [7:0] t_r1_c41_9;
  wire [7:0] t_r1_c41_10;
  wire [7:0] t_r1_c41_11;
  wire [7:0] t_r1_c41_12;
  wire [7:0] t_r1_c42_0;
  wire [7:0] t_r1_c42_1;
  wire [7:0] t_r1_c42_2;
  wire [7:0] t_r1_c42_3;
  wire [7:0] t_r1_c42_4;
  wire [7:0] t_r1_c42_5;
  wire [7:0] t_r1_c42_6;
  wire [7:0] t_r1_c42_7;
  wire [7:0] t_r1_c42_8;
  wire [7:0] t_r1_c42_9;
  wire [7:0] t_r1_c42_10;
  wire [7:0] t_r1_c42_11;
  wire [7:0] t_r1_c42_12;
  wire [7:0] t_r1_c43_0;
  wire [7:0] t_r1_c43_1;
  wire [7:0] t_r1_c43_2;
  wire [7:0] t_r1_c43_3;
  wire [7:0] t_r1_c43_4;
  wire [7:0] t_r1_c43_5;
  wire [7:0] t_r1_c43_6;
  wire [7:0] t_r1_c43_7;
  wire [7:0] t_r1_c43_8;
  wire [7:0] t_r1_c43_9;
  wire [7:0] t_r1_c43_10;
  wire [7:0] t_r1_c43_11;
  wire [7:0] t_r1_c43_12;
  wire [7:0] t_r1_c44_0;
  wire [7:0] t_r1_c44_1;
  wire [7:0] t_r1_c44_2;
  wire [7:0] t_r1_c44_3;
  wire [7:0] t_r1_c44_4;
  wire [7:0] t_r1_c44_5;
  wire [7:0] t_r1_c44_6;
  wire [7:0] t_r1_c44_7;
  wire [7:0] t_r1_c44_8;
  wire [7:0] t_r1_c44_9;
  wire [7:0] t_r1_c44_10;
  wire [7:0] t_r1_c44_11;
  wire [7:0] t_r1_c44_12;
  wire [7:0] t_r1_c45_0;
  wire [7:0] t_r1_c45_1;
  wire [7:0] t_r1_c45_2;
  wire [7:0] t_r1_c45_3;
  wire [7:0] t_r1_c45_4;
  wire [7:0] t_r1_c45_5;
  wire [7:0] t_r1_c45_6;
  wire [7:0] t_r1_c45_7;
  wire [7:0] t_r1_c45_8;
  wire [7:0] t_r1_c45_9;
  wire [7:0] t_r1_c45_10;
  wire [7:0] t_r1_c45_11;
  wire [7:0] t_r1_c45_12;
  wire [7:0] t_r1_c46_0;
  wire [7:0] t_r1_c46_1;
  wire [7:0] t_r1_c46_2;
  wire [7:0] t_r1_c46_3;
  wire [7:0] t_r1_c46_4;
  wire [7:0] t_r1_c46_5;
  wire [7:0] t_r1_c46_6;
  wire [7:0] t_r1_c46_7;
  wire [7:0] t_r1_c46_8;
  wire [7:0] t_r1_c46_9;
  wire [7:0] t_r1_c46_10;
  wire [7:0] t_r1_c46_11;
  wire [7:0] t_r1_c46_12;
  wire [7:0] t_r1_c47_0;
  wire [7:0] t_r1_c47_1;
  wire [7:0] t_r1_c47_2;
  wire [7:0] t_r1_c47_3;
  wire [7:0] t_r1_c47_4;
  wire [7:0] t_r1_c47_5;
  wire [7:0] t_r1_c47_6;
  wire [7:0] t_r1_c47_7;
  wire [7:0] t_r1_c47_8;
  wire [7:0] t_r1_c47_9;
  wire [7:0] t_r1_c47_10;
  wire [7:0] t_r1_c47_11;
  wire [7:0] t_r1_c47_12;
  wire [7:0] t_r1_c48_0;
  wire [7:0] t_r1_c48_1;
  wire [7:0] t_r1_c48_2;
  wire [7:0] t_r1_c48_3;
  wire [7:0] t_r1_c48_4;
  wire [7:0] t_r1_c48_5;
  wire [7:0] t_r1_c48_6;
  wire [7:0] t_r1_c48_7;
  wire [7:0] t_r1_c48_8;
  wire [7:0] t_r1_c48_9;
  wire [7:0] t_r1_c48_10;
  wire [7:0] t_r1_c48_11;
  wire [7:0] t_r1_c48_12;
  wire [7:0] t_r1_c49_0;
  wire [7:0] t_r1_c49_1;
  wire [7:0] t_r1_c49_2;
  wire [7:0] t_r1_c49_3;
  wire [7:0] t_r1_c49_4;
  wire [7:0] t_r1_c49_5;
  wire [7:0] t_r1_c49_6;
  wire [7:0] t_r1_c49_7;
  wire [7:0] t_r1_c49_8;
  wire [7:0] t_r1_c49_9;
  wire [7:0] t_r1_c49_10;
  wire [7:0] t_r1_c49_11;
  wire [7:0] t_r1_c49_12;
  wire [7:0] t_r1_c50_0;
  wire [7:0] t_r1_c50_1;
  wire [7:0] t_r1_c50_2;
  wire [7:0] t_r1_c50_3;
  wire [7:0] t_r1_c50_4;
  wire [7:0] t_r1_c50_5;
  wire [7:0] t_r1_c50_6;
  wire [7:0] t_r1_c50_7;
  wire [7:0] t_r1_c50_8;
  wire [7:0] t_r1_c50_9;
  wire [7:0] t_r1_c50_10;
  wire [7:0] t_r1_c50_11;
  wire [7:0] t_r1_c50_12;
  wire [7:0] t_r1_c51_0;
  wire [7:0] t_r1_c51_1;
  wire [7:0] t_r1_c51_2;
  wire [7:0] t_r1_c51_3;
  wire [7:0] t_r1_c51_4;
  wire [7:0] t_r1_c51_5;
  wire [7:0] t_r1_c51_6;
  wire [7:0] t_r1_c51_7;
  wire [7:0] t_r1_c51_8;
  wire [7:0] t_r1_c51_9;
  wire [7:0] t_r1_c51_10;
  wire [7:0] t_r1_c51_11;
  wire [7:0] t_r1_c51_12;
  wire [7:0] t_r1_c52_0;
  wire [7:0] t_r1_c52_1;
  wire [7:0] t_r1_c52_2;
  wire [7:0] t_r1_c52_3;
  wire [7:0] t_r1_c52_4;
  wire [7:0] t_r1_c52_5;
  wire [7:0] t_r1_c52_6;
  wire [7:0] t_r1_c52_7;
  wire [7:0] t_r1_c52_8;
  wire [7:0] t_r1_c52_9;
  wire [7:0] t_r1_c52_10;
  wire [7:0] t_r1_c52_11;
  wire [7:0] t_r1_c52_12;
  wire [7:0] t_r1_c53_0;
  wire [7:0] t_r1_c53_1;
  wire [7:0] t_r1_c53_2;
  wire [7:0] t_r1_c53_3;
  wire [7:0] t_r1_c53_4;
  wire [7:0] t_r1_c53_5;
  wire [7:0] t_r1_c53_6;
  wire [7:0] t_r1_c53_7;
  wire [7:0] t_r1_c53_8;
  wire [7:0] t_r1_c53_9;
  wire [7:0] t_r1_c53_10;
  wire [7:0] t_r1_c53_11;
  wire [7:0] t_r1_c53_12;
  wire [7:0] t_r1_c54_0;
  wire [7:0] t_r1_c54_1;
  wire [7:0] t_r1_c54_2;
  wire [7:0] t_r1_c54_3;
  wire [7:0] t_r1_c54_4;
  wire [7:0] t_r1_c54_5;
  wire [7:0] t_r1_c54_6;
  wire [7:0] t_r1_c54_7;
  wire [7:0] t_r1_c54_8;
  wire [7:0] t_r1_c54_9;
  wire [7:0] t_r1_c54_10;
  wire [7:0] t_r1_c54_11;
  wire [7:0] t_r1_c54_12;
  wire [7:0] t_r1_c55_0;
  wire [7:0] t_r1_c55_1;
  wire [7:0] t_r1_c55_2;
  wire [7:0] t_r1_c55_3;
  wire [7:0] t_r1_c55_4;
  wire [7:0] t_r1_c55_5;
  wire [7:0] t_r1_c55_6;
  wire [7:0] t_r1_c55_7;
  wire [7:0] t_r1_c55_8;
  wire [7:0] t_r1_c55_9;
  wire [7:0] t_r1_c55_10;
  wire [7:0] t_r1_c55_11;
  wire [7:0] t_r1_c55_12;
  wire [7:0] t_r1_c56_0;
  wire [7:0] t_r1_c56_1;
  wire [7:0] t_r1_c56_2;
  wire [7:0] t_r1_c56_3;
  wire [7:0] t_r1_c56_4;
  wire [7:0] t_r1_c56_5;
  wire [7:0] t_r1_c56_6;
  wire [7:0] t_r1_c56_7;
  wire [7:0] t_r1_c56_8;
  wire [7:0] t_r1_c56_9;
  wire [7:0] t_r1_c56_10;
  wire [7:0] t_r1_c56_11;
  wire [7:0] t_r1_c56_12;
  wire [7:0] t_r1_c57_0;
  wire [7:0] t_r1_c57_1;
  wire [7:0] t_r1_c57_2;
  wire [7:0] t_r1_c57_3;
  wire [7:0] t_r1_c57_4;
  wire [7:0] t_r1_c57_5;
  wire [7:0] t_r1_c57_6;
  wire [7:0] t_r1_c57_7;
  wire [7:0] t_r1_c57_8;
  wire [7:0] t_r1_c57_9;
  wire [7:0] t_r1_c57_10;
  wire [7:0] t_r1_c57_11;
  wire [7:0] t_r1_c57_12;
  wire [7:0] t_r1_c58_0;
  wire [7:0] t_r1_c58_1;
  wire [7:0] t_r1_c58_2;
  wire [7:0] t_r1_c58_3;
  wire [7:0] t_r1_c58_4;
  wire [7:0] t_r1_c58_5;
  wire [7:0] t_r1_c58_6;
  wire [7:0] t_r1_c58_7;
  wire [7:0] t_r1_c58_8;
  wire [7:0] t_r1_c58_9;
  wire [7:0] t_r1_c58_10;
  wire [7:0] t_r1_c58_11;
  wire [7:0] t_r1_c58_12;
  wire [7:0] t_r1_c59_0;
  wire [7:0] t_r1_c59_1;
  wire [7:0] t_r1_c59_2;
  wire [7:0] t_r1_c59_3;
  wire [7:0] t_r1_c59_4;
  wire [7:0] t_r1_c59_5;
  wire [7:0] t_r1_c59_6;
  wire [7:0] t_r1_c59_7;
  wire [7:0] t_r1_c59_8;
  wire [7:0] t_r1_c59_9;
  wire [7:0] t_r1_c59_10;
  wire [7:0] t_r1_c59_11;
  wire [7:0] t_r1_c59_12;
  wire [7:0] t_r1_c60_0;
  wire [7:0] t_r1_c60_1;
  wire [7:0] t_r1_c60_2;
  wire [7:0] t_r1_c60_3;
  wire [7:0] t_r1_c60_4;
  wire [7:0] t_r1_c60_5;
  wire [7:0] t_r1_c60_6;
  wire [7:0] t_r1_c60_7;
  wire [7:0] t_r1_c60_8;
  wire [7:0] t_r1_c60_9;
  wire [7:0] t_r1_c60_10;
  wire [7:0] t_r1_c60_11;
  wire [7:0] t_r1_c60_12;
  wire [7:0] t_r1_c61_0;
  wire [7:0] t_r1_c61_1;
  wire [7:0] t_r1_c61_2;
  wire [7:0] t_r1_c61_3;
  wire [7:0] t_r1_c61_4;
  wire [7:0] t_r1_c61_5;
  wire [7:0] t_r1_c61_6;
  wire [7:0] t_r1_c61_7;
  wire [7:0] t_r1_c61_8;
  wire [7:0] t_r1_c61_9;
  wire [7:0] t_r1_c61_10;
  wire [7:0] t_r1_c61_11;
  wire [7:0] t_r1_c61_12;
  wire [7:0] t_r1_c62_0;
  wire [7:0] t_r1_c62_1;
  wire [7:0] t_r1_c62_2;
  wire [7:0] t_r1_c62_3;
  wire [7:0] t_r1_c62_4;
  wire [7:0] t_r1_c62_5;
  wire [7:0] t_r1_c62_6;
  wire [7:0] t_r1_c62_7;
  wire [7:0] t_r1_c62_8;
  wire [7:0] t_r1_c62_9;
  wire [7:0] t_r1_c62_10;
  wire [7:0] t_r1_c62_11;
  wire [7:0] t_r1_c62_12;
  wire [7:0] t_r1_c63_0;
  wire [7:0] t_r1_c63_1;
  wire [7:0] t_r1_c63_2;
  wire [7:0] t_r1_c63_3;
  wire [7:0] t_r1_c63_4;
  wire [7:0] t_r1_c63_5;
  wire [7:0] t_r1_c63_6;
  wire [7:0] t_r1_c63_7;
  wire [7:0] t_r1_c63_8;
  wire [7:0] t_r1_c63_9;
  wire [7:0] t_r1_c63_10;
  wire [7:0] t_r1_c63_11;
  wire [7:0] t_r1_c63_12;
  wire [7:0] t_r1_c64_0;
  wire [7:0] t_r1_c64_1;
  wire [7:0] t_r1_c64_2;
  wire [7:0] t_r1_c64_3;
  wire [7:0] t_r1_c64_4;
  wire [7:0] t_r1_c64_5;
  wire [7:0] t_r1_c64_6;
  wire [7:0] t_r1_c64_7;
  wire [7:0] t_r1_c64_8;
  wire [7:0] t_r1_c64_9;
  wire [7:0] t_r1_c64_10;
  wire [7:0] t_r1_c64_11;
  wire [7:0] t_r1_c64_12;
  wire [7:0] t_r1_c65_0;
  wire [7:0] t_r1_c65_1;
  wire [7:0] t_r1_c65_2;
  wire [7:0] t_r1_c65_3;
  wire [7:0] t_r1_c65_4;
  wire [7:0] t_r1_c65_5;
  wire [7:0] t_r1_c65_6;
  wire [7:0] t_r1_c65_7;
  wire [7:0] t_r1_c65_8;
  wire [7:0] t_r1_c65_9;
  wire [7:0] t_r1_c65_10;
  wire [7:0] t_r1_c65_11;
  wire [7:0] t_r1_c65_12;
  wire [7:0] t_r2_c0_0;
  wire [7:0] t_r2_c0_1;
  wire [7:0] t_r2_c0_2;
  wire [7:0] t_r2_c0_3;
  wire [7:0] t_r2_c0_4;
  wire [7:0] t_r2_c0_5;
  wire [7:0] t_r2_c0_6;
  wire [7:0] t_r2_c0_7;
  wire [7:0] t_r2_c0_8;
  wire [7:0] t_r2_c0_9;
  wire [7:0] t_r2_c0_10;
  wire [7:0] t_r2_c0_11;
  wire [7:0] t_r2_c0_12;
  wire [7:0] t_r2_c1_0;
  wire [7:0] t_r2_c1_1;
  wire [7:0] t_r2_c1_2;
  wire [7:0] t_r2_c1_3;
  wire [7:0] t_r2_c1_4;
  wire [7:0] t_r2_c1_5;
  wire [7:0] t_r2_c1_6;
  wire [7:0] t_r2_c1_7;
  wire [7:0] t_r2_c1_8;
  wire [7:0] t_r2_c1_9;
  wire [7:0] t_r2_c1_10;
  wire [7:0] t_r2_c1_11;
  wire [7:0] t_r2_c1_12;
  wire [7:0] t_r2_c2_0;
  wire [7:0] t_r2_c2_1;
  wire [7:0] t_r2_c2_2;
  wire [7:0] t_r2_c2_3;
  wire [7:0] t_r2_c2_4;
  wire [7:0] t_r2_c2_5;
  wire [7:0] t_r2_c2_6;
  wire [7:0] t_r2_c2_7;
  wire [7:0] t_r2_c2_8;
  wire [7:0] t_r2_c2_9;
  wire [7:0] t_r2_c2_10;
  wire [7:0] t_r2_c2_11;
  wire [7:0] t_r2_c2_12;
  wire [7:0] t_r2_c3_0;
  wire [7:0] t_r2_c3_1;
  wire [7:0] t_r2_c3_2;
  wire [7:0] t_r2_c3_3;
  wire [7:0] t_r2_c3_4;
  wire [7:0] t_r2_c3_5;
  wire [7:0] t_r2_c3_6;
  wire [7:0] t_r2_c3_7;
  wire [7:0] t_r2_c3_8;
  wire [7:0] t_r2_c3_9;
  wire [7:0] t_r2_c3_10;
  wire [7:0] t_r2_c3_11;
  wire [7:0] t_r2_c3_12;
  wire [7:0] t_r2_c4_0;
  wire [7:0] t_r2_c4_1;
  wire [7:0] t_r2_c4_2;
  wire [7:0] t_r2_c4_3;
  wire [7:0] t_r2_c4_4;
  wire [7:0] t_r2_c4_5;
  wire [7:0] t_r2_c4_6;
  wire [7:0] t_r2_c4_7;
  wire [7:0] t_r2_c4_8;
  wire [7:0] t_r2_c4_9;
  wire [7:0] t_r2_c4_10;
  wire [7:0] t_r2_c4_11;
  wire [7:0] t_r2_c4_12;
  wire [7:0] t_r2_c5_0;
  wire [7:0] t_r2_c5_1;
  wire [7:0] t_r2_c5_2;
  wire [7:0] t_r2_c5_3;
  wire [7:0] t_r2_c5_4;
  wire [7:0] t_r2_c5_5;
  wire [7:0] t_r2_c5_6;
  wire [7:0] t_r2_c5_7;
  wire [7:0] t_r2_c5_8;
  wire [7:0] t_r2_c5_9;
  wire [7:0] t_r2_c5_10;
  wire [7:0] t_r2_c5_11;
  wire [7:0] t_r2_c5_12;
  wire [7:0] t_r2_c6_0;
  wire [7:0] t_r2_c6_1;
  wire [7:0] t_r2_c6_2;
  wire [7:0] t_r2_c6_3;
  wire [7:0] t_r2_c6_4;
  wire [7:0] t_r2_c6_5;
  wire [7:0] t_r2_c6_6;
  wire [7:0] t_r2_c6_7;
  wire [7:0] t_r2_c6_8;
  wire [7:0] t_r2_c6_9;
  wire [7:0] t_r2_c6_10;
  wire [7:0] t_r2_c6_11;
  wire [7:0] t_r2_c6_12;
  wire [7:0] t_r2_c7_0;
  wire [7:0] t_r2_c7_1;
  wire [7:0] t_r2_c7_2;
  wire [7:0] t_r2_c7_3;
  wire [7:0] t_r2_c7_4;
  wire [7:0] t_r2_c7_5;
  wire [7:0] t_r2_c7_6;
  wire [7:0] t_r2_c7_7;
  wire [7:0] t_r2_c7_8;
  wire [7:0] t_r2_c7_9;
  wire [7:0] t_r2_c7_10;
  wire [7:0] t_r2_c7_11;
  wire [7:0] t_r2_c7_12;
  wire [7:0] t_r2_c8_0;
  wire [7:0] t_r2_c8_1;
  wire [7:0] t_r2_c8_2;
  wire [7:0] t_r2_c8_3;
  wire [7:0] t_r2_c8_4;
  wire [7:0] t_r2_c8_5;
  wire [7:0] t_r2_c8_6;
  wire [7:0] t_r2_c8_7;
  wire [7:0] t_r2_c8_8;
  wire [7:0] t_r2_c8_9;
  wire [7:0] t_r2_c8_10;
  wire [7:0] t_r2_c8_11;
  wire [7:0] t_r2_c8_12;
  wire [7:0] t_r2_c9_0;
  wire [7:0] t_r2_c9_1;
  wire [7:0] t_r2_c9_2;
  wire [7:0] t_r2_c9_3;
  wire [7:0] t_r2_c9_4;
  wire [7:0] t_r2_c9_5;
  wire [7:0] t_r2_c9_6;
  wire [7:0] t_r2_c9_7;
  wire [7:0] t_r2_c9_8;
  wire [7:0] t_r2_c9_9;
  wire [7:0] t_r2_c9_10;
  wire [7:0] t_r2_c9_11;
  wire [7:0] t_r2_c9_12;
  wire [7:0] t_r2_c10_0;
  wire [7:0] t_r2_c10_1;
  wire [7:0] t_r2_c10_2;
  wire [7:0] t_r2_c10_3;
  wire [7:0] t_r2_c10_4;
  wire [7:0] t_r2_c10_5;
  wire [7:0] t_r2_c10_6;
  wire [7:0] t_r2_c10_7;
  wire [7:0] t_r2_c10_8;
  wire [7:0] t_r2_c10_9;
  wire [7:0] t_r2_c10_10;
  wire [7:0] t_r2_c10_11;
  wire [7:0] t_r2_c10_12;
  wire [7:0] t_r2_c11_0;
  wire [7:0] t_r2_c11_1;
  wire [7:0] t_r2_c11_2;
  wire [7:0] t_r2_c11_3;
  wire [7:0] t_r2_c11_4;
  wire [7:0] t_r2_c11_5;
  wire [7:0] t_r2_c11_6;
  wire [7:0] t_r2_c11_7;
  wire [7:0] t_r2_c11_8;
  wire [7:0] t_r2_c11_9;
  wire [7:0] t_r2_c11_10;
  wire [7:0] t_r2_c11_11;
  wire [7:0] t_r2_c11_12;
  wire [7:0] t_r2_c12_0;
  wire [7:0] t_r2_c12_1;
  wire [7:0] t_r2_c12_2;
  wire [7:0] t_r2_c12_3;
  wire [7:0] t_r2_c12_4;
  wire [7:0] t_r2_c12_5;
  wire [7:0] t_r2_c12_6;
  wire [7:0] t_r2_c12_7;
  wire [7:0] t_r2_c12_8;
  wire [7:0] t_r2_c12_9;
  wire [7:0] t_r2_c12_10;
  wire [7:0] t_r2_c12_11;
  wire [7:0] t_r2_c12_12;
  wire [7:0] t_r2_c13_0;
  wire [7:0] t_r2_c13_1;
  wire [7:0] t_r2_c13_2;
  wire [7:0] t_r2_c13_3;
  wire [7:0] t_r2_c13_4;
  wire [7:0] t_r2_c13_5;
  wire [7:0] t_r2_c13_6;
  wire [7:0] t_r2_c13_7;
  wire [7:0] t_r2_c13_8;
  wire [7:0] t_r2_c13_9;
  wire [7:0] t_r2_c13_10;
  wire [7:0] t_r2_c13_11;
  wire [7:0] t_r2_c13_12;
  wire [7:0] t_r2_c14_0;
  wire [7:0] t_r2_c14_1;
  wire [7:0] t_r2_c14_2;
  wire [7:0] t_r2_c14_3;
  wire [7:0] t_r2_c14_4;
  wire [7:0] t_r2_c14_5;
  wire [7:0] t_r2_c14_6;
  wire [7:0] t_r2_c14_7;
  wire [7:0] t_r2_c14_8;
  wire [7:0] t_r2_c14_9;
  wire [7:0] t_r2_c14_10;
  wire [7:0] t_r2_c14_11;
  wire [7:0] t_r2_c14_12;
  wire [7:0] t_r2_c15_0;
  wire [7:0] t_r2_c15_1;
  wire [7:0] t_r2_c15_2;
  wire [7:0] t_r2_c15_3;
  wire [7:0] t_r2_c15_4;
  wire [7:0] t_r2_c15_5;
  wire [7:0] t_r2_c15_6;
  wire [7:0] t_r2_c15_7;
  wire [7:0] t_r2_c15_8;
  wire [7:0] t_r2_c15_9;
  wire [7:0] t_r2_c15_10;
  wire [7:0] t_r2_c15_11;
  wire [7:0] t_r2_c15_12;
  wire [7:0] t_r2_c16_0;
  wire [7:0] t_r2_c16_1;
  wire [7:0] t_r2_c16_2;
  wire [7:0] t_r2_c16_3;
  wire [7:0] t_r2_c16_4;
  wire [7:0] t_r2_c16_5;
  wire [7:0] t_r2_c16_6;
  wire [7:0] t_r2_c16_7;
  wire [7:0] t_r2_c16_8;
  wire [7:0] t_r2_c16_9;
  wire [7:0] t_r2_c16_10;
  wire [7:0] t_r2_c16_11;
  wire [7:0] t_r2_c16_12;
  wire [7:0] t_r2_c17_0;
  wire [7:0] t_r2_c17_1;
  wire [7:0] t_r2_c17_2;
  wire [7:0] t_r2_c17_3;
  wire [7:0] t_r2_c17_4;
  wire [7:0] t_r2_c17_5;
  wire [7:0] t_r2_c17_6;
  wire [7:0] t_r2_c17_7;
  wire [7:0] t_r2_c17_8;
  wire [7:0] t_r2_c17_9;
  wire [7:0] t_r2_c17_10;
  wire [7:0] t_r2_c17_11;
  wire [7:0] t_r2_c17_12;
  wire [7:0] t_r2_c18_0;
  wire [7:0] t_r2_c18_1;
  wire [7:0] t_r2_c18_2;
  wire [7:0] t_r2_c18_3;
  wire [7:0] t_r2_c18_4;
  wire [7:0] t_r2_c18_5;
  wire [7:0] t_r2_c18_6;
  wire [7:0] t_r2_c18_7;
  wire [7:0] t_r2_c18_8;
  wire [7:0] t_r2_c18_9;
  wire [7:0] t_r2_c18_10;
  wire [7:0] t_r2_c18_11;
  wire [7:0] t_r2_c18_12;
  wire [7:0] t_r2_c19_0;
  wire [7:0] t_r2_c19_1;
  wire [7:0] t_r2_c19_2;
  wire [7:0] t_r2_c19_3;
  wire [7:0] t_r2_c19_4;
  wire [7:0] t_r2_c19_5;
  wire [7:0] t_r2_c19_6;
  wire [7:0] t_r2_c19_7;
  wire [7:0] t_r2_c19_8;
  wire [7:0] t_r2_c19_9;
  wire [7:0] t_r2_c19_10;
  wire [7:0] t_r2_c19_11;
  wire [7:0] t_r2_c19_12;
  wire [7:0] t_r2_c20_0;
  wire [7:0] t_r2_c20_1;
  wire [7:0] t_r2_c20_2;
  wire [7:0] t_r2_c20_3;
  wire [7:0] t_r2_c20_4;
  wire [7:0] t_r2_c20_5;
  wire [7:0] t_r2_c20_6;
  wire [7:0] t_r2_c20_7;
  wire [7:0] t_r2_c20_8;
  wire [7:0] t_r2_c20_9;
  wire [7:0] t_r2_c20_10;
  wire [7:0] t_r2_c20_11;
  wire [7:0] t_r2_c20_12;
  wire [7:0] t_r2_c21_0;
  wire [7:0] t_r2_c21_1;
  wire [7:0] t_r2_c21_2;
  wire [7:0] t_r2_c21_3;
  wire [7:0] t_r2_c21_4;
  wire [7:0] t_r2_c21_5;
  wire [7:0] t_r2_c21_6;
  wire [7:0] t_r2_c21_7;
  wire [7:0] t_r2_c21_8;
  wire [7:0] t_r2_c21_9;
  wire [7:0] t_r2_c21_10;
  wire [7:0] t_r2_c21_11;
  wire [7:0] t_r2_c21_12;
  wire [7:0] t_r2_c22_0;
  wire [7:0] t_r2_c22_1;
  wire [7:0] t_r2_c22_2;
  wire [7:0] t_r2_c22_3;
  wire [7:0] t_r2_c22_4;
  wire [7:0] t_r2_c22_5;
  wire [7:0] t_r2_c22_6;
  wire [7:0] t_r2_c22_7;
  wire [7:0] t_r2_c22_8;
  wire [7:0] t_r2_c22_9;
  wire [7:0] t_r2_c22_10;
  wire [7:0] t_r2_c22_11;
  wire [7:0] t_r2_c22_12;
  wire [7:0] t_r2_c23_0;
  wire [7:0] t_r2_c23_1;
  wire [7:0] t_r2_c23_2;
  wire [7:0] t_r2_c23_3;
  wire [7:0] t_r2_c23_4;
  wire [7:0] t_r2_c23_5;
  wire [7:0] t_r2_c23_6;
  wire [7:0] t_r2_c23_7;
  wire [7:0] t_r2_c23_8;
  wire [7:0] t_r2_c23_9;
  wire [7:0] t_r2_c23_10;
  wire [7:0] t_r2_c23_11;
  wire [7:0] t_r2_c23_12;
  wire [7:0] t_r2_c24_0;
  wire [7:0] t_r2_c24_1;
  wire [7:0] t_r2_c24_2;
  wire [7:0] t_r2_c24_3;
  wire [7:0] t_r2_c24_4;
  wire [7:0] t_r2_c24_5;
  wire [7:0] t_r2_c24_6;
  wire [7:0] t_r2_c24_7;
  wire [7:0] t_r2_c24_8;
  wire [7:0] t_r2_c24_9;
  wire [7:0] t_r2_c24_10;
  wire [7:0] t_r2_c24_11;
  wire [7:0] t_r2_c24_12;
  wire [7:0] t_r2_c25_0;
  wire [7:0] t_r2_c25_1;
  wire [7:0] t_r2_c25_2;
  wire [7:0] t_r2_c25_3;
  wire [7:0] t_r2_c25_4;
  wire [7:0] t_r2_c25_5;
  wire [7:0] t_r2_c25_6;
  wire [7:0] t_r2_c25_7;
  wire [7:0] t_r2_c25_8;
  wire [7:0] t_r2_c25_9;
  wire [7:0] t_r2_c25_10;
  wire [7:0] t_r2_c25_11;
  wire [7:0] t_r2_c25_12;
  wire [7:0] t_r2_c26_0;
  wire [7:0] t_r2_c26_1;
  wire [7:0] t_r2_c26_2;
  wire [7:0] t_r2_c26_3;
  wire [7:0] t_r2_c26_4;
  wire [7:0] t_r2_c26_5;
  wire [7:0] t_r2_c26_6;
  wire [7:0] t_r2_c26_7;
  wire [7:0] t_r2_c26_8;
  wire [7:0] t_r2_c26_9;
  wire [7:0] t_r2_c26_10;
  wire [7:0] t_r2_c26_11;
  wire [7:0] t_r2_c26_12;
  wire [7:0] t_r2_c27_0;
  wire [7:0] t_r2_c27_1;
  wire [7:0] t_r2_c27_2;
  wire [7:0] t_r2_c27_3;
  wire [7:0] t_r2_c27_4;
  wire [7:0] t_r2_c27_5;
  wire [7:0] t_r2_c27_6;
  wire [7:0] t_r2_c27_7;
  wire [7:0] t_r2_c27_8;
  wire [7:0] t_r2_c27_9;
  wire [7:0] t_r2_c27_10;
  wire [7:0] t_r2_c27_11;
  wire [7:0] t_r2_c27_12;
  wire [7:0] t_r2_c28_0;
  wire [7:0] t_r2_c28_1;
  wire [7:0] t_r2_c28_2;
  wire [7:0] t_r2_c28_3;
  wire [7:0] t_r2_c28_4;
  wire [7:0] t_r2_c28_5;
  wire [7:0] t_r2_c28_6;
  wire [7:0] t_r2_c28_7;
  wire [7:0] t_r2_c28_8;
  wire [7:0] t_r2_c28_9;
  wire [7:0] t_r2_c28_10;
  wire [7:0] t_r2_c28_11;
  wire [7:0] t_r2_c28_12;
  wire [7:0] t_r2_c29_0;
  wire [7:0] t_r2_c29_1;
  wire [7:0] t_r2_c29_2;
  wire [7:0] t_r2_c29_3;
  wire [7:0] t_r2_c29_4;
  wire [7:0] t_r2_c29_5;
  wire [7:0] t_r2_c29_6;
  wire [7:0] t_r2_c29_7;
  wire [7:0] t_r2_c29_8;
  wire [7:0] t_r2_c29_9;
  wire [7:0] t_r2_c29_10;
  wire [7:0] t_r2_c29_11;
  wire [7:0] t_r2_c29_12;
  wire [7:0] t_r2_c30_0;
  wire [7:0] t_r2_c30_1;
  wire [7:0] t_r2_c30_2;
  wire [7:0] t_r2_c30_3;
  wire [7:0] t_r2_c30_4;
  wire [7:0] t_r2_c30_5;
  wire [7:0] t_r2_c30_6;
  wire [7:0] t_r2_c30_7;
  wire [7:0] t_r2_c30_8;
  wire [7:0] t_r2_c30_9;
  wire [7:0] t_r2_c30_10;
  wire [7:0] t_r2_c30_11;
  wire [7:0] t_r2_c30_12;
  wire [7:0] t_r2_c31_0;
  wire [7:0] t_r2_c31_1;
  wire [7:0] t_r2_c31_2;
  wire [7:0] t_r2_c31_3;
  wire [7:0] t_r2_c31_4;
  wire [7:0] t_r2_c31_5;
  wire [7:0] t_r2_c31_6;
  wire [7:0] t_r2_c31_7;
  wire [7:0] t_r2_c31_8;
  wire [7:0] t_r2_c31_9;
  wire [7:0] t_r2_c31_10;
  wire [7:0] t_r2_c31_11;
  wire [7:0] t_r2_c31_12;
  wire [7:0] t_r2_c32_0;
  wire [7:0] t_r2_c32_1;
  wire [7:0] t_r2_c32_2;
  wire [7:0] t_r2_c32_3;
  wire [7:0] t_r2_c32_4;
  wire [7:0] t_r2_c32_5;
  wire [7:0] t_r2_c32_6;
  wire [7:0] t_r2_c32_7;
  wire [7:0] t_r2_c32_8;
  wire [7:0] t_r2_c32_9;
  wire [7:0] t_r2_c32_10;
  wire [7:0] t_r2_c32_11;
  wire [7:0] t_r2_c32_12;
  wire [7:0] t_r2_c33_0;
  wire [7:0] t_r2_c33_1;
  wire [7:0] t_r2_c33_2;
  wire [7:0] t_r2_c33_3;
  wire [7:0] t_r2_c33_4;
  wire [7:0] t_r2_c33_5;
  wire [7:0] t_r2_c33_6;
  wire [7:0] t_r2_c33_7;
  wire [7:0] t_r2_c33_8;
  wire [7:0] t_r2_c33_9;
  wire [7:0] t_r2_c33_10;
  wire [7:0] t_r2_c33_11;
  wire [7:0] t_r2_c33_12;
  wire [7:0] t_r2_c34_0;
  wire [7:0] t_r2_c34_1;
  wire [7:0] t_r2_c34_2;
  wire [7:0] t_r2_c34_3;
  wire [7:0] t_r2_c34_4;
  wire [7:0] t_r2_c34_5;
  wire [7:0] t_r2_c34_6;
  wire [7:0] t_r2_c34_7;
  wire [7:0] t_r2_c34_8;
  wire [7:0] t_r2_c34_9;
  wire [7:0] t_r2_c34_10;
  wire [7:0] t_r2_c34_11;
  wire [7:0] t_r2_c34_12;
  wire [7:0] t_r2_c35_0;
  wire [7:0] t_r2_c35_1;
  wire [7:0] t_r2_c35_2;
  wire [7:0] t_r2_c35_3;
  wire [7:0] t_r2_c35_4;
  wire [7:0] t_r2_c35_5;
  wire [7:0] t_r2_c35_6;
  wire [7:0] t_r2_c35_7;
  wire [7:0] t_r2_c35_8;
  wire [7:0] t_r2_c35_9;
  wire [7:0] t_r2_c35_10;
  wire [7:0] t_r2_c35_11;
  wire [7:0] t_r2_c35_12;
  wire [7:0] t_r2_c36_0;
  wire [7:0] t_r2_c36_1;
  wire [7:0] t_r2_c36_2;
  wire [7:0] t_r2_c36_3;
  wire [7:0] t_r2_c36_4;
  wire [7:0] t_r2_c36_5;
  wire [7:0] t_r2_c36_6;
  wire [7:0] t_r2_c36_7;
  wire [7:0] t_r2_c36_8;
  wire [7:0] t_r2_c36_9;
  wire [7:0] t_r2_c36_10;
  wire [7:0] t_r2_c36_11;
  wire [7:0] t_r2_c36_12;
  wire [7:0] t_r2_c37_0;
  wire [7:0] t_r2_c37_1;
  wire [7:0] t_r2_c37_2;
  wire [7:0] t_r2_c37_3;
  wire [7:0] t_r2_c37_4;
  wire [7:0] t_r2_c37_5;
  wire [7:0] t_r2_c37_6;
  wire [7:0] t_r2_c37_7;
  wire [7:0] t_r2_c37_8;
  wire [7:0] t_r2_c37_9;
  wire [7:0] t_r2_c37_10;
  wire [7:0] t_r2_c37_11;
  wire [7:0] t_r2_c37_12;
  wire [7:0] t_r2_c38_0;
  wire [7:0] t_r2_c38_1;
  wire [7:0] t_r2_c38_2;
  wire [7:0] t_r2_c38_3;
  wire [7:0] t_r2_c38_4;
  wire [7:0] t_r2_c38_5;
  wire [7:0] t_r2_c38_6;
  wire [7:0] t_r2_c38_7;
  wire [7:0] t_r2_c38_8;
  wire [7:0] t_r2_c38_9;
  wire [7:0] t_r2_c38_10;
  wire [7:0] t_r2_c38_11;
  wire [7:0] t_r2_c38_12;
  wire [7:0] t_r2_c39_0;
  wire [7:0] t_r2_c39_1;
  wire [7:0] t_r2_c39_2;
  wire [7:0] t_r2_c39_3;
  wire [7:0] t_r2_c39_4;
  wire [7:0] t_r2_c39_5;
  wire [7:0] t_r2_c39_6;
  wire [7:0] t_r2_c39_7;
  wire [7:0] t_r2_c39_8;
  wire [7:0] t_r2_c39_9;
  wire [7:0] t_r2_c39_10;
  wire [7:0] t_r2_c39_11;
  wire [7:0] t_r2_c39_12;
  wire [7:0] t_r2_c40_0;
  wire [7:0] t_r2_c40_1;
  wire [7:0] t_r2_c40_2;
  wire [7:0] t_r2_c40_3;
  wire [7:0] t_r2_c40_4;
  wire [7:0] t_r2_c40_5;
  wire [7:0] t_r2_c40_6;
  wire [7:0] t_r2_c40_7;
  wire [7:0] t_r2_c40_8;
  wire [7:0] t_r2_c40_9;
  wire [7:0] t_r2_c40_10;
  wire [7:0] t_r2_c40_11;
  wire [7:0] t_r2_c40_12;
  wire [7:0] t_r2_c41_0;
  wire [7:0] t_r2_c41_1;
  wire [7:0] t_r2_c41_2;
  wire [7:0] t_r2_c41_3;
  wire [7:0] t_r2_c41_4;
  wire [7:0] t_r2_c41_5;
  wire [7:0] t_r2_c41_6;
  wire [7:0] t_r2_c41_7;
  wire [7:0] t_r2_c41_8;
  wire [7:0] t_r2_c41_9;
  wire [7:0] t_r2_c41_10;
  wire [7:0] t_r2_c41_11;
  wire [7:0] t_r2_c41_12;
  wire [7:0] t_r2_c42_0;
  wire [7:0] t_r2_c42_1;
  wire [7:0] t_r2_c42_2;
  wire [7:0] t_r2_c42_3;
  wire [7:0] t_r2_c42_4;
  wire [7:0] t_r2_c42_5;
  wire [7:0] t_r2_c42_6;
  wire [7:0] t_r2_c42_7;
  wire [7:0] t_r2_c42_8;
  wire [7:0] t_r2_c42_9;
  wire [7:0] t_r2_c42_10;
  wire [7:0] t_r2_c42_11;
  wire [7:0] t_r2_c42_12;
  wire [7:0] t_r2_c43_0;
  wire [7:0] t_r2_c43_1;
  wire [7:0] t_r2_c43_2;
  wire [7:0] t_r2_c43_3;
  wire [7:0] t_r2_c43_4;
  wire [7:0] t_r2_c43_5;
  wire [7:0] t_r2_c43_6;
  wire [7:0] t_r2_c43_7;
  wire [7:0] t_r2_c43_8;
  wire [7:0] t_r2_c43_9;
  wire [7:0] t_r2_c43_10;
  wire [7:0] t_r2_c43_11;
  wire [7:0] t_r2_c43_12;
  wire [7:0] t_r2_c44_0;
  wire [7:0] t_r2_c44_1;
  wire [7:0] t_r2_c44_2;
  wire [7:0] t_r2_c44_3;
  wire [7:0] t_r2_c44_4;
  wire [7:0] t_r2_c44_5;
  wire [7:0] t_r2_c44_6;
  wire [7:0] t_r2_c44_7;
  wire [7:0] t_r2_c44_8;
  wire [7:0] t_r2_c44_9;
  wire [7:0] t_r2_c44_10;
  wire [7:0] t_r2_c44_11;
  wire [7:0] t_r2_c44_12;
  wire [7:0] t_r2_c45_0;
  wire [7:0] t_r2_c45_1;
  wire [7:0] t_r2_c45_2;
  wire [7:0] t_r2_c45_3;
  wire [7:0] t_r2_c45_4;
  wire [7:0] t_r2_c45_5;
  wire [7:0] t_r2_c45_6;
  wire [7:0] t_r2_c45_7;
  wire [7:0] t_r2_c45_8;
  wire [7:0] t_r2_c45_9;
  wire [7:0] t_r2_c45_10;
  wire [7:0] t_r2_c45_11;
  wire [7:0] t_r2_c45_12;
  wire [7:0] t_r2_c46_0;
  wire [7:0] t_r2_c46_1;
  wire [7:0] t_r2_c46_2;
  wire [7:0] t_r2_c46_3;
  wire [7:0] t_r2_c46_4;
  wire [7:0] t_r2_c46_5;
  wire [7:0] t_r2_c46_6;
  wire [7:0] t_r2_c46_7;
  wire [7:0] t_r2_c46_8;
  wire [7:0] t_r2_c46_9;
  wire [7:0] t_r2_c46_10;
  wire [7:0] t_r2_c46_11;
  wire [7:0] t_r2_c46_12;
  wire [7:0] t_r2_c47_0;
  wire [7:0] t_r2_c47_1;
  wire [7:0] t_r2_c47_2;
  wire [7:0] t_r2_c47_3;
  wire [7:0] t_r2_c47_4;
  wire [7:0] t_r2_c47_5;
  wire [7:0] t_r2_c47_6;
  wire [7:0] t_r2_c47_7;
  wire [7:0] t_r2_c47_8;
  wire [7:0] t_r2_c47_9;
  wire [7:0] t_r2_c47_10;
  wire [7:0] t_r2_c47_11;
  wire [7:0] t_r2_c47_12;
  wire [7:0] t_r2_c48_0;
  wire [7:0] t_r2_c48_1;
  wire [7:0] t_r2_c48_2;
  wire [7:0] t_r2_c48_3;
  wire [7:0] t_r2_c48_4;
  wire [7:0] t_r2_c48_5;
  wire [7:0] t_r2_c48_6;
  wire [7:0] t_r2_c48_7;
  wire [7:0] t_r2_c48_8;
  wire [7:0] t_r2_c48_9;
  wire [7:0] t_r2_c48_10;
  wire [7:0] t_r2_c48_11;
  wire [7:0] t_r2_c48_12;
  wire [7:0] t_r2_c49_0;
  wire [7:0] t_r2_c49_1;
  wire [7:0] t_r2_c49_2;
  wire [7:0] t_r2_c49_3;
  wire [7:0] t_r2_c49_4;
  wire [7:0] t_r2_c49_5;
  wire [7:0] t_r2_c49_6;
  wire [7:0] t_r2_c49_7;
  wire [7:0] t_r2_c49_8;
  wire [7:0] t_r2_c49_9;
  wire [7:0] t_r2_c49_10;
  wire [7:0] t_r2_c49_11;
  wire [7:0] t_r2_c49_12;
  wire [7:0] t_r2_c50_0;
  wire [7:0] t_r2_c50_1;
  wire [7:0] t_r2_c50_2;
  wire [7:0] t_r2_c50_3;
  wire [7:0] t_r2_c50_4;
  wire [7:0] t_r2_c50_5;
  wire [7:0] t_r2_c50_6;
  wire [7:0] t_r2_c50_7;
  wire [7:0] t_r2_c50_8;
  wire [7:0] t_r2_c50_9;
  wire [7:0] t_r2_c50_10;
  wire [7:0] t_r2_c50_11;
  wire [7:0] t_r2_c50_12;
  wire [7:0] t_r2_c51_0;
  wire [7:0] t_r2_c51_1;
  wire [7:0] t_r2_c51_2;
  wire [7:0] t_r2_c51_3;
  wire [7:0] t_r2_c51_4;
  wire [7:0] t_r2_c51_5;
  wire [7:0] t_r2_c51_6;
  wire [7:0] t_r2_c51_7;
  wire [7:0] t_r2_c51_8;
  wire [7:0] t_r2_c51_9;
  wire [7:0] t_r2_c51_10;
  wire [7:0] t_r2_c51_11;
  wire [7:0] t_r2_c51_12;
  wire [7:0] t_r2_c52_0;
  wire [7:0] t_r2_c52_1;
  wire [7:0] t_r2_c52_2;
  wire [7:0] t_r2_c52_3;
  wire [7:0] t_r2_c52_4;
  wire [7:0] t_r2_c52_5;
  wire [7:0] t_r2_c52_6;
  wire [7:0] t_r2_c52_7;
  wire [7:0] t_r2_c52_8;
  wire [7:0] t_r2_c52_9;
  wire [7:0] t_r2_c52_10;
  wire [7:0] t_r2_c52_11;
  wire [7:0] t_r2_c52_12;
  wire [7:0] t_r2_c53_0;
  wire [7:0] t_r2_c53_1;
  wire [7:0] t_r2_c53_2;
  wire [7:0] t_r2_c53_3;
  wire [7:0] t_r2_c53_4;
  wire [7:0] t_r2_c53_5;
  wire [7:0] t_r2_c53_6;
  wire [7:0] t_r2_c53_7;
  wire [7:0] t_r2_c53_8;
  wire [7:0] t_r2_c53_9;
  wire [7:0] t_r2_c53_10;
  wire [7:0] t_r2_c53_11;
  wire [7:0] t_r2_c53_12;
  wire [7:0] t_r2_c54_0;
  wire [7:0] t_r2_c54_1;
  wire [7:0] t_r2_c54_2;
  wire [7:0] t_r2_c54_3;
  wire [7:0] t_r2_c54_4;
  wire [7:0] t_r2_c54_5;
  wire [7:0] t_r2_c54_6;
  wire [7:0] t_r2_c54_7;
  wire [7:0] t_r2_c54_8;
  wire [7:0] t_r2_c54_9;
  wire [7:0] t_r2_c54_10;
  wire [7:0] t_r2_c54_11;
  wire [7:0] t_r2_c54_12;
  wire [7:0] t_r2_c55_0;
  wire [7:0] t_r2_c55_1;
  wire [7:0] t_r2_c55_2;
  wire [7:0] t_r2_c55_3;
  wire [7:0] t_r2_c55_4;
  wire [7:0] t_r2_c55_5;
  wire [7:0] t_r2_c55_6;
  wire [7:0] t_r2_c55_7;
  wire [7:0] t_r2_c55_8;
  wire [7:0] t_r2_c55_9;
  wire [7:0] t_r2_c55_10;
  wire [7:0] t_r2_c55_11;
  wire [7:0] t_r2_c55_12;
  wire [7:0] t_r2_c56_0;
  wire [7:0] t_r2_c56_1;
  wire [7:0] t_r2_c56_2;
  wire [7:0] t_r2_c56_3;
  wire [7:0] t_r2_c56_4;
  wire [7:0] t_r2_c56_5;
  wire [7:0] t_r2_c56_6;
  wire [7:0] t_r2_c56_7;
  wire [7:0] t_r2_c56_8;
  wire [7:0] t_r2_c56_9;
  wire [7:0] t_r2_c56_10;
  wire [7:0] t_r2_c56_11;
  wire [7:0] t_r2_c56_12;
  wire [7:0] t_r2_c57_0;
  wire [7:0] t_r2_c57_1;
  wire [7:0] t_r2_c57_2;
  wire [7:0] t_r2_c57_3;
  wire [7:0] t_r2_c57_4;
  wire [7:0] t_r2_c57_5;
  wire [7:0] t_r2_c57_6;
  wire [7:0] t_r2_c57_7;
  wire [7:0] t_r2_c57_8;
  wire [7:0] t_r2_c57_9;
  wire [7:0] t_r2_c57_10;
  wire [7:0] t_r2_c57_11;
  wire [7:0] t_r2_c57_12;
  wire [7:0] t_r2_c58_0;
  wire [7:0] t_r2_c58_1;
  wire [7:0] t_r2_c58_2;
  wire [7:0] t_r2_c58_3;
  wire [7:0] t_r2_c58_4;
  wire [7:0] t_r2_c58_5;
  wire [7:0] t_r2_c58_6;
  wire [7:0] t_r2_c58_7;
  wire [7:0] t_r2_c58_8;
  wire [7:0] t_r2_c58_9;
  wire [7:0] t_r2_c58_10;
  wire [7:0] t_r2_c58_11;
  wire [7:0] t_r2_c58_12;
  wire [7:0] t_r2_c59_0;
  wire [7:0] t_r2_c59_1;
  wire [7:0] t_r2_c59_2;
  wire [7:0] t_r2_c59_3;
  wire [7:0] t_r2_c59_4;
  wire [7:0] t_r2_c59_5;
  wire [7:0] t_r2_c59_6;
  wire [7:0] t_r2_c59_7;
  wire [7:0] t_r2_c59_8;
  wire [7:0] t_r2_c59_9;
  wire [7:0] t_r2_c59_10;
  wire [7:0] t_r2_c59_11;
  wire [7:0] t_r2_c59_12;
  wire [7:0] t_r2_c60_0;
  wire [7:0] t_r2_c60_1;
  wire [7:0] t_r2_c60_2;
  wire [7:0] t_r2_c60_3;
  wire [7:0] t_r2_c60_4;
  wire [7:0] t_r2_c60_5;
  wire [7:0] t_r2_c60_6;
  wire [7:0] t_r2_c60_7;
  wire [7:0] t_r2_c60_8;
  wire [7:0] t_r2_c60_9;
  wire [7:0] t_r2_c60_10;
  wire [7:0] t_r2_c60_11;
  wire [7:0] t_r2_c60_12;
  wire [7:0] t_r2_c61_0;
  wire [7:0] t_r2_c61_1;
  wire [7:0] t_r2_c61_2;
  wire [7:0] t_r2_c61_3;
  wire [7:0] t_r2_c61_4;
  wire [7:0] t_r2_c61_5;
  wire [7:0] t_r2_c61_6;
  wire [7:0] t_r2_c61_7;
  wire [7:0] t_r2_c61_8;
  wire [7:0] t_r2_c61_9;
  wire [7:0] t_r2_c61_10;
  wire [7:0] t_r2_c61_11;
  wire [7:0] t_r2_c61_12;
  wire [7:0] t_r2_c62_0;
  wire [7:0] t_r2_c62_1;
  wire [7:0] t_r2_c62_2;
  wire [7:0] t_r2_c62_3;
  wire [7:0] t_r2_c62_4;
  wire [7:0] t_r2_c62_5;
  wire [7:0] t_r2_c62_6;
  wire [7:0] t_r2_c62_7;
  wire [7:0] t_r2_c62_8;
  wire [7:0] t_r2_c62_9;
  wire [7:0] t_r2_c62_10;
  wire [7:0] t_r2_c62_11;
  wire [7:0] t_r2_c62_12;
  wire [7:0] t_r2_c63_0;
  wire [7:0] t_r2_c63_1;
  wire [7:0] t_r2_c63_2;
  wire [7:0] t_r2_c63_3;
  wire [7:0] t_r2_c63_4;
  wire [7:0] t_r2_c63_5;
  wire [7:0] t_r2_c63_6;
  wire [7:0] t_r2_c63_7;
  wire [7:0] t_r2_c63_8;
  wire [7:0] t_r2_c63_9;
  wire [7:0] t_r2_c63_10;
  wire [7:0] t_r2_c63_11;
  wire [7:0] t_r2_c63_12;
  wire [7:0] t_r2_c64_0;
  wire [7:0] t_r2_c64_1;
  wire [7:0] t_r2_c64_2;
  wire [7:0] t_r2_c64_3;
  wire [7:0] t_r2_c64_4;
  wire [7:0] t_r2_c64_5;
  wire [7:0] t_r2_c64_6;
  wire [7:0] t_r2_c64_7;
  wire [7:0] t_r2_c64_8;
  wire [7:0] t_r2_c64_9;
  wire [7:0] t_r2_c64_10;
  wire [7:0] t_r2_c64_11;
  wire [7:0] t_r2_c64_12;
  wire [7:0] t_r2_c65_0;
  wire [7:0] t_r2_c65_1;
  wire [7:0] t_r2_c65_2;
  wire [7:0] t_r2_c65_3;
  wire [7:0] t_r2_c65_4;
  wire [7:0] t_r2_c65_5;
  wire [7:0] t_r2_c65_6;
  wire [7:0] t_r2_c65_7;
  wire [7:0] t_r2_c65_8;
  wire [7:0] t_r2_c65_9;
  wire [7:0] t_r2_c65_10;
  wire [7:0] t_r2_c65_11;
  wire [7:0] t_r2_c65_12;
  wire [7:0] t_r3_c0_0;
  wire [7:0] t_r3_c0_1;
  wire [7:0] t_r3_c0_2;
  wire [7:0] t_r3_c0_3;
  wire [7:0] t_r3_c0_4;
  wire [7:0] t_r3_c0_5;
  wire [7:0] t_r3_c0_6;
  wire [7:0] t_r3_c0_7;
  wire [7:0] t_r3_c0_8;
  wire [7:0] t_r3_c0_9;
  wire [7:0] t_r3_c0_10;
  wire [7:0] t_r3_c0_11;
  wire [7:0] t_r3_c0_12;
  wire [7:0] t_r3_c1_0;
  wire [7:0] t_r3_c1_1;
  wire [7:0] t_r3_c1_2;
  wire [7:0] t_r3_c1_3;
  wire [7:0] t_r3_c1_4;
  wire [7:0] t_r3_c1_5;
  wire [7:0] t_r3_c1_6;
  wire [7:0] t_r3_c1_7;
  wire [7:0] t_r3_c1_8;
  wire [7:0] t_r3_c1_9;
  wire [7:0] t_r3_c1_10;
  wire [7:0] t_r3_c1_11;
  wire [7:0] t_r3_c1_12;
  wire [7:0] t_r3_c2_0;
  wire [7:0] t_r3_c2_1;
  wire [7:0] t_r3_c2_2;
  wire [7:0] t_r3_c2_3;
  wire [7:0] t_r3_c2_4;
  wire [7:0] t_r3_c2_5;
  wire [7:0] t_r3_c2_6;
  wire [7:0] t_r3_c2_7;
  wire [7:0] t_r3_c2_8;
  wire [7:0] t_r3_c2_9;
  wire [7:0] t_r3_c2_10;
  wire [7:0] t_r3_c2_11;
  wire [7:0] t_r3_c2_12;
  wire [7:0] t_r3_c3_0;
  wire [7:0] t_r3_c3_1;
  wire [7:0] t_r3_c3_2;
  wire [7:0] t_r3_c3_3;
  wire [7:0] t_r3_c3_4;
  wire [7:0] t_r3_c3_5;
  wire [7:0] t_r3_c3_6;
  wire [7:0] t_r3_c3_7;
  wire [7:0] t_r3_c3_8;
  wire [7:0] t_r3_c3_9;
  wire [7:0] t_r3_c3_10;
  wire [7:0] t_r3_c3_11;
  wire [7:0] t_r3_c3_12;
  wire [7:0] t_r3_c4_0;
  wire [7:0] t_r3_c4_1;
  wire [7:0] t_r3_c4_2;
  wire [7:0] t_r3_c4_3;
  wire [7:0] t_r3_c4_4;
  wire [7:0] t_r3_c4_5;
  wire [7:0] t_r3_c4_6;
  wire [7:0] t_r3_c4_7;
  wire [7:0] t_r3_c4_8;
  wire [7:0] t_r3_c4_9;
  wire [7:0] t_r3_c4_10;
  wire [7:0] t_r3_c4_11;
  wire [7:0] t_r3_c4_12;
  wire [7:0] t_r3_c5_0;
  wire [7:0] t_r3_c5_1;
  wire [7:0] t_r3_c5_2;
  wire [7:0] t_r3_c5_3;
  wire [7:0] t_r3_c5_4;
  wire [7:0] t_r3_c5_5;
  wire [7:0] t_r3_c5_6;
  wire [7:0] t_r3_c5_7;
  wire [7:0] t_r3_c5_8;
  wire [7:0] t_r3_c5_9;
  wire [7:0] t_r3_c5_10;
  wire [7:0] t_r3_c5_11;
  wire [7:0] t_r3_c5_12;
  wire [7:0] t_r3_c6_0;
  wire [7:0] t_r3_c6_1;
  wire [7:0] t_r3_c6_2;
  wire [7:0] t_r3_c6_3;
  wire [7:0] t_r3_c6_4;
  wire [7:0] t_r3_c6_5;
  wire [7:0] t_r3_c6_6;
  wire [7:0] t_r3_c6_7;
  wire [7:0] t_r3_c6_8;
  wire [7:0] t_r3_c6_9;
  wire [7:0] t_r3_c6_10;
  wire [7:0] t_r3_c6_11;
  wire [7:0] t_r3_c6_12;
  wire [7:0] t_r3_c7_0;
  wire [7:0] t_r3_c7_1;
  wire [7:0] t_r3_c7_2;
  wire [7:0] t_r3_c7_3;
  wire [7:0] t_r3_c7_4;
  wire [7:0] t_r3_c7_5;
  wire [7:0] t_r3_c7_6;
  wire [7:0] t_r3_c7_7;
  wire [7:0] t_r3_c7_8;
  wire [7:0] t_r3_c7_9;
  wire [7:0] t_r3_c7_10;
  wire [7:0] t_r3_c7_11;
  wire [7:0] t_r3_c7_12;
  wire [7:0] t_r3_c8_0;
  wire [7:0] t_r3_c8_1;
  wire [7:0] t_r3_c8_2;
  wire [7:0] t_r3_c8_3;
  wire [7:0] t_r3_c8_4;
  wire [7:0] t_r3_c8_5;
  wire [7:0] t_r3_c8_6;
  wire [7:0] t_r3_c8_7;
  wire [7:0] t_r3_c8_8;
  wire [7:0] t_r3_c8_9;
  wire [7:0] t_r3_c8_10;
  wire [7:0] t_r3_c8_11;
  wire [7:0] t_r3_c8_12;
  wire [7:0] t_r3_c9_0;
  wire [7:0] t_r3_c9_1;
  wire [7:0] t_r3_c9_2;
  wire [7:0] t_r3_c9_3;
  wire [7:0] t_r3_c9_4;
  wire [7:0] t_r3_c9_5;
  wire [7:0] t_r3_c9_6;
  wire [7:0] t_r3_c9_7;
  wire [7:0] t_r3_c9_8;
  wire [7:0] t_r3_c9_9;
  wire [7:0] t_r3_c9_10;
  wire [7:0] t_r3_c9_11;
  wire [7:0] t_r3_c9_12;
  wire [7:0] t_r3_c10_0;
  wire [7:0] t_r3_c10_1;
  wire [7:0] t_r3_c10_2;
  wire [7:0] t_r3_c10_3;
  wire [7:0] t_r3_c10_4;
  wire [7:0] t_r3_c10_5;
  wire [7:0] t_r3_c10_6;
  wire [7:0] t_r3_c10_7;
  wire [7:0] t_r3_c10_8;
  wire [7:0] t_r3_c10_9;
  wire [7:0] t_r3_c10_10;
  wire [7:0] t_r3_c10_11;
  wire [7:0] t_r3_c10_12;
  wire [7:0] t_r3_c11_0;
  wire [7:0] t_r3_c11_1;
  wire [7:0] t_r3_c11_2;
  wire [7:0] t_r3_c11_3;
  wire [7:0] t_r3_c11_4;
  wire [7:0] t_r3_c11_5;
  wire [7:0] t_r3_c11_6;
  wire [7:0] t_r3_c11_7;
  wire [7:0] t_r3_c11_8;
  wire [7:0] t_r3_c11_9;
  wire [7:0] t_r3_c11_10;
  wire [7:0] t_r3_c11_11;
  wire [7:0] t_r3_c11_12;
  wire [7:0] t_r3_c12_0;
  wire [7:0] t_r3_c12_1;
  wire [7:0] t_r3_c12_2;
  wire [7:0] t_r3_c12_3;
  wire [7:0] t_r3_c12_4;
  wire [7:0] t_r3_c12_5;
  wire [7:0] t_r3_c12_6;
  wire [7:0] t_r3_c12_7;
  wire [7:0] t_r3_c12_8;
  wire [7:0] t_r3_c12_9;
  wire [7:0] t_r3_c12_10;
  wire [7:0] t_r3_c12_11;
  wire [7:0] t_r3_c12_12;
  wire [7:0] t_r3_c13_0;
  wire [7:0] t_r3_c13_1;
  wire [7:0] t_r3_c13_2;
  wire [7:0] t_r3_c13_3;
  wire [7:0] t_r3_c13_4;
  wire [7:0] t_r3_c13_5;
  wire [7:0] t_r3_c13_6;
  wire [7:0] t_r3_c13_7;
  wire [7:0] t_r3_c13_8;
  wire [7:0] t_r3_c13_9;
  wire [7:0] t_r3_c13_10;
  wire [7:0] t_r3_c13_11;
  wire [7:0] t_r3_c13_12;
  wire [7:0] t_r3_c14_0;
  wire [7:0] t_r3_c14_1;
  wire [7:0] t_r3_c14_2;
  wire [7:0] t_r3_c14_3;
  wire [7:0] t_r3_c14_4;
  wire [7:0] t_r3_c14_5;
  wire [7:0] t_r3_c14_6;
  wire [7:0] t_r3_c14_7;
  wire [7:0] t_r3_c14_8;
  wire [7:0] t_r3_c14_9;
  wire [7:0] t_r3_c14_10;
  wire [7:0] t_r3_c14_11;
  wire [7:0] t_r3_c14_12;
  wire [7:0] t_r3_c15_0;
  wire [7:0] t_r3_c15_1;
  wire [7:0] t_r3_c15_2;
  wire [7:0] t_r3_c15_3;
  wire [7:0] t_r3_c15_4;
  wire [7:0] t_r3_c15_5;
  wire [7:0] t_r3_c15_6;
  wire [7:0] t_r3_c15_7;
  wire [7:0] t_r3_c15_8;
  wire [7:0] t_r3_c15_9;
  wire [7:0] t_r3_c15_10;
  wire [7:0] t_r3_c15_11;
  wire [7:0] t_r3_c15_12;
  wire [7:0] t_r3_c16_0;
  wire [7:0] t_r3_c16_1;
  wire [7:0] t_r3_c16_2;
  wire [7:0] t_r3_c16_3;
  wire [7:0] t_r3_c16_4;
  wire [7:0] t_r3_c16_5;
  wire [7:0] t_r3_c16_6;
  wire [7:0] t_r3_c16_7;
  wire [7:0] t_r3_c16_8;
  wire [7:0] t_r3_c16_9;
  wire [7:0] t_r3_c16_10;
  wire [7:0] t_r3_c16_11;
  wire [7:0] t_r3_c16_12;
  wire [7:0] t_r3_c17_0;
  wire [7:0] t_r3_c17_1;
  wire [7:0] t_r3_c17_2;
  wire [7:0] t_r3_c17_3;
  wire [7:0] t_r3_c17_4;
  wire [7:0] t_r3_c17_5;
  wire [7:0] t_r3_c17_6;
  wire [7:0] t_r3_c17_7;
  wire [7:0] t_r3_c17_8;
  wire [7:0] t_r3_c17_9;
  wire [7:0] t_r3_c17_10;
  wire [7:0] t_r3_c17_11;
  wire [7:0] t_r3_c17_12;
  wire [7:0] t_r3_c18_0;
  wire [7:0] t_r3_c18_1;
  wire [7:0] t_r3_c18_2;
  wire [7:0] t_r3_c18_3;
  wire [7:0] t_r3_c18_4;
  wire [7:0] t_r3_c18_5;
  wire [7:0] t_r3_c18_6;
  wire [7:0] t_r3_c18_7;
  wire [7:0] t_r3_c18_8;
  wire [7:0] t_r3_c18_9;
  wire [7:0] t_r3_c18_10;
  wire [7:0] t_r3_c18_11;
  wire [7:0] t_r3_c18_12;
  wire [7:0] t_r3_c19_0;
  wire [7:0] t_r3_c19_1;
  wire [7:0] t_r3_c19_2;
  wire [7:0] t_r3_c19_3;
  wire [7:0] t_r3_c19_4;
  wire [7:0] t_r3_c19_5;
  wire [7:0] t_r3_c19_6;
  wire [7:0] t_r3_c19_7;
  wire [7:0] t_r3_c19_8;
  wire [7:0] t_r3_c19_9;
  wire [7:0] t_r3_c19_10;
  wire [7:0] t_r3_c19_11;
  wire [7:0] t_r3_c19_12;
  wire [7:0] t_r3_c20_0;
  wire [7:0] t_r3_c20_1;
  wire [7:0] t_r3_c20_2;
  wire [7:0] t_r3_c20_3;
  wire [7:0] t_r3_c20_4;
  wire [7:0] t_r3_c20_5;
  wire [7:0] t_r3_c20_6;
  wire [7:0] t_r3_c20_7;
  wire [7:0] t_r3_c20_8;
  wire [7:0] t_r3_c20_9;
  wire [7:0] t_r3_c20_10;
  wire [7:0] t_r3_c20_11;
  wire [7:0] t_r3_c20_12;
  wire [7:0] t_r3_c21_0;
  wire [7:0] t_r3_c21_1;
  wire [7:0] t_r3_c21_2;
  wire [7:0] t_r3_c21_3;
  wire [7:0] t_r3_c21_4;
  wire [7:0] t_r3_c21_5;
  wire [7:0] t_r3_c21_6;
  wire [7:0] t_r3_c21_7;
  wire [7:0] t_r3_c21_8;
  wire [7:0] t_r3_c21_9;
  wire [7:0] t_r3_c21_10;
  wire [7:0] t_r3_c21_11;
  wire [7:0] t_r3_c21_12;
  wire [7:0] t_r3_c22_0;
  wire [7:0] t_r3_c22_1;
  wire [7:0] t_r3_c22_2;
  wire [7:0] t_r3_c22_3;
  wire [7:0] t_r3_c22_4;
  wire [7:0] t_r3_c22_5;
  wire [7:0] t_r3_c22_6;
  wire [7:0] t_r3_c22_7;
  wire [7:0] t_r3_c22_8;
  wire [7:0] t_r3_c22_9;
  wire [7:0] t_r3_c22_10;
  wire [7:0] t_r3_c22_11;
  wire [7:0] t_r3_c22_12;
  wire [7:0] t_r3_c23_0;
  wire [7:0] t_r3_c23_1;
  wire [7:0] t_r3_c23_2;
  wire [7:0] t_r3_c23_3;
  wire [7:0] t_r3_c23_4;
  wire [7:0] t_r3_c23_5;
  wire [7:0] t_r3_c23_6;
  wire [7:0] t_r3_c23_7;
  wire [7:0] t_r3_c23_8;
  wire [7:0] t_r3_c23_9;
  wire [7:0] t_r3_c23_10;
  wire [7:0] t_r3_c23_11;
  wire [7:0] t_r3_c23_12;
  wire [7:0] t_r3_c24_0;
  wire [7:0] t_r3_c24_1;
  wire [7:0] t_r3_c24_2;
  wire [7:0] t_r3_c24_3;
  wire [7:0] t_r3_c24_4;
  wire [7:0] t_r3_c24_5;
  wire [7:0] t_r3_c24_6;
  wire [7:0] t_r3_c24_7;
  wire [7:0] t_r3_c24_8;
  wire [7:0] t_r3_c24_9;
  wire [7:0] t_r3_c24_10;
  wire [7:0] t_r3_c24_11;
  wire [7:0] t_r3_c24_12;
  wire [7:0] t_r3_c25_0;
  wire [7:0] t_r3_c25_1;
  wire [7:0] t_r3_c25_2;
  wire [7:0] t_r3_c25_3;
  wire [7:0] t_r3_c25_4;
  wire [7:0] t_r3_c25_5;
  wire [7:0] t_r3_c25_6;
  wire [7:0] t_r3_c25_7;
  wire [7:0] t_r3_c25_8;
  wire [7:0] t_r3_c25_9;
  wire [7:0] t_r3_c25_10;
  wire [7:0] t_r3_c25_11;
  wire [7:0] t_r3_c25_12;
  wire [7:0] t_r3_c26_0;
  wire [7:0] t_r3_c26_1;
  wire [7:0] t_r3_c26_2;
  wire [7:0] t_r3_c26_3;
  wire [7:0] t_r3_c26_4;
  wire [7:0] t_r3_c26_5;
  wire [7:0] t_r3_c26_6;
  wire [7:0] t_r3_c26_7;
  wire [7:0] t_r3_c26_8;
  wire [7:0] t_r3_c26_9;
  wire [7:0] t_r3_c26_10;
  wire [7:0] t_r3_c26_11;
  wire [7:0] t_r3_c26_12;
  wire [7:0] t_r3_c27_0;
  wire [7:0] t_r3_c27_1;
  wire [7:0] t_r3_c27_2;
  wire [7:0] t_r3_c27_3;
  wire [7:0] t_r3_c27_4;
  wire [7:0] t_r3_c27_5;
  wire [7:0] t_r3_c27_6;
  wire [7:0] t_r3_c27_7;
  wire [7:0] t_r3_c27_8;
  wire [7:0] t_r3_c27_9;
  wire [7:0] t_r3_c27_10;
  wire [7:0] t_r3_c27_11;
  wire [7:0] t_r3_c27_12;
  wire [7:0] t_r3_c28_0;
  wire [7:0] t_r3_c28_1;
  wire [7:0] t_r3_c28_2;
  wire [7:0] t_r3_c28_3;
  wire [7:0] t_r3_c28_4;
  wire [7:0] t_r3_c28_5;
  wire [7:0] t_r3_c28_6;
  wire [7:0] t_r3_c28_7;
  wire [7:0] t_r3_c28_8;
  wire [7:0] t_r3_c28_9;
  wire [7:0] t_r3_c28_10;
  wire [7:0] t_r3_c28_11;
  wire [7:0] t_r3_c28_12;
  wire [7:0] t_r3_c29_0;
  wire [7:0] t_r3_c29_1;
  wire [7:0] t_r3_c29_2;
  wire [7:0] t_r3_c29_3;
  wire [7:0] t_r3_c29_4;
  wire [7:0] t_r3_c29_5;
  wire [7:0] t_r3_c29_6;
  wire [7:0] t_r3_c29_7;
  wire [7:0] t_r3_c29_8;
  wire [7:0] t_r3_c29_9;
  wire [7:0] t_r3_c29_10;
  wire [7:0] t_r3_c29_11;
  wire [7:0] t_r3_c29_12;
  wire [7:0] t_r3_c30_0;
  wire [7:0] t_r3_c30_1;
  wire [7:0] t_r3_c30_2;
  wire [7:0] t_r3_c30_3;
  wire [7:0] t_r3_c30_4;
  wire [7:0] t_r3_c30_5;
  wire [7:0] t_r3_c30_6;
  wire [7:0] t_r3_c30_7;
  wire [7:0] t_r3_c30_8;
  wire [7:0] t_r3_c30_9;
  wire [7:0] t_r3_c30_10;
  wire [7:0] t_r3_c30_11;
  wire [7:0] t_r3_c30_12;
  wire [7:0] t_r3_c31_0;
  wire [7:0] t_r3_c31_1;
  wire [7:0] t_r3_c31_2;
  wire [7:0] t_r3_c31_3;
  wire [7:0] t_r3_c31_4;
  wire [7:0] t_r3_c31_5;
  wire [7:0] t_r3_c31_6;
  wire [7:0] t_r3_c31_7;
  wire [7:0] t_r3_c31_8;
  wire [7:0] t_r3_c31_9;
  wire [7:0] t_r3_c31_10;
  wire [7:0] t_r3_c31_11;
  wire [7:0] t_r3_c31_12;
  wire [7:0] t_r3_c32_0;
  wire [7:0] t_r3_c32_1;
  wire [7:0] t_r3_c32_2;
  wire [7:0] t_r3_c32_3;
  wire [7:0] t_r3_c32_4;
  wire [7:0] t_r3_c32_5;
  wire [7:0] t_r3_c32_6;
  wire [7:0] t_r3_c32_7;
  wire [7:0] t_r3_c32_8;
  wire [7:0] t_r3_c32_9;
  wire [7:0] t_r3_c32_10;
  wire [7:0] t_r3_c32_11;
  wire [7:0] t_r3_c32_12;
  wire [7:0] t_r3_c33_0;
  wire [7:0] t_r3_c33_1;
  wire [7:0] t_r3_c33_2;
  wire [7:0] t_r3_c33_3;
  wire [7:0] t_r3_c33_4;
  wire [7:0] t_r3_c33_5;
  wire [7:0] t_r3_c33_6;
  wire [7:0] t_r3_c33_7;
  wire [7:0] t_r3_c33_8;
  wire [7:0] t_r3_c33_9;
  wire [7:0] t_r3_c33_10;
  wire [7:0] t_r3_c33_11;
  wire [7:0] t_r3_c33_12;
  wire [7:0] t_r3_c34_0;
  wire [7:0] t_r3_c34_1;
  wire [7:0] t_r3_c34_2;
  wire [7:0] t_r3_c34_3;
  wire [7:0] t_r3_c34_4;
  wire [7:0] t_r3_c34_5;
  wire [7:0] t_r3_c34_6;
  wire [7:0] t_r3_c34_7;
  wire [7:0] t_r3_c34_8;
  wire [7:0] t_r3_c34_9;
  wire [7:0] t_r3_c34_10;
  wire [7:0] t_r3_c34_11;
  wire [7:0] t_r3_c34_12;
  wire [7:0] t_r3_c35_0;
  wire [7:0] t_r3_c35_1;
  wire [7:0] t_r3_c35_2;
  wire [7:0] t_r3_c35_3;
  wire [7:0] t_r3_c35_4;
  wire [7:0] t_r3_c35_5;
  wire [7:0] t_r3_c35_6;
  wire [7:0] t_r3_c35_7;
  wire [7:0] t_r3_c35_8;
  wire [7:0] t_r3_c35_9;
  wire [7:0] t_r3_c35_10;
  wire [7:0] t_r3_c35_11;
  wire [7:0] t_r3_c35_12;
  wire [7:0] t_r3_c36_0;
  wire [7:0] t_r3_c36_1;
  wire [7:0] t_r3_c36_2;
  wire [7:0] t_r3_c36_3;
  wire [7:0] t_r3_c36_4;
  wire [7:0] t_r3_c36_5;
  wire [7:0] t_r3_c36_6;
  wire [7:0] t_r3_c36_7;
  wire [7:0] t_r3_c36_8;
  wire [7:0] t_r3_c36_9;
  wire [7:0] t_r3_c36_10;
  wire [7:0] t_r3_c36_11;
  wire [7:0] t_r3_c36_12;
  wire [7:0] t_r3_c37_0;
  wire [7:0] t_r3_c37_1;
  wire [7:0] t_r3_c37_2;
  wire [7:0] t_r3_c37_3;
  wire [7:0] t_r3_c37_4;
  wire [7:0] t_r3_c37_5;
  wire [7:0] t_r3_c37_6;
  wire [7:0] t_r3_c37_7;
  wire [7:0] t_r3_c37_8;
  wire [7:0] t_r3_c37_9;
  wire [7:0] t_r3_c37_10;
  wire [7:0] t_r3_c37_11;
  wire [7:0] t_r3_c37_12;
  wire [7:0] t_r3_c38_0;
  wire [7:0] t_r3_c38_1;
  wire [7:0] t_r3_c38_2;
  wire [7:0] t_r3_c38_3;
  wire [7:0] t_r3_c38_4;
  wire [7:0] t_r3_c38_5;
  wire [7:0] t_r3_c38_6;
  wire [7:0] t_r3_c38_7;
  wire [7:0] t_r3_c38_8;
  wire [7:0] t_r3_c38_9;
  wire [7:0] t_r3_c38_10;
  wire [7:0] t_r3_c38_11;
  wire [7:0] t_r3_c38_12;
  wire [7:0] t_r3_c39_0;
  wire [7:0] t_r3_c39_1;
  wire [7:0] t_r3_c39_2;
  wire [7:0] t_r3_c39_3;
  wire [7:0] t_r3_c39_4;
  wire [7:0] t_r3_c39_5;
  wire [7:0] t_r3_c39_6;
  wire [7:0] t_r3_c39_7;
  wire [7:0] t_r3_c39_8;
  wire [7:0] t_r3_c39_9;
  wire [7:0] t_r3_c39_10;
  wire [7:0] t_r3_c39_11;
  wire [7:0] t_r3_c39_12;
  wire [7:0] t_r3_c40_0;
  wire [7:0] t_r3_c40_1;
  wire [7:0] t_r3_c40_2;
  wire [7:0] t_r3_c40_3;
  wire [7:0] t_r3_c40_4;
  wire [7:0] t_r3_c40_5;
  wire [7:0] t_r3_c40_6;
  wire [7:0] t_r3_c40_7;
  wire [7:0] t_r3_c40_8;
  wire [7:0] t_r3_c40_9;
  wire [7:0] t_r3_c40_10;
  wire [7:0] t_r3_c40_11;
  wire [7:0] t_r3_c40_12;
  wire [7:0] t_r3_c41_0;
  wire [7:0] t_r3_c41_1;
  wire [7:0] t_r3_c41_2;
  wire [7:0] t_r3_c41_3;
  wire [7:0] t_r3_c41_4;
  wire [7:0] t_r3_c41_5;
  wire [7:0] t_r3_c41_6;
  wire [7:0] t_r3_c41_7;
  wire [7:0] t_r3_c41_8;
  wire [7:0] t_r3_c41_9;
  wire [7:0] t_r3_c41_10;
  wire [7:0] t_r3_c41_11;
  wire [7:0] t_r3_c41_12;
  wire [7:0] t_r3_c42_0;
  wire [7:0] t_r3_c42_1;
  wire [7:0] t_r3_c42_2;
  wire [7:0] t_r3_c42_3;
  wire [7:0] t_r3_c42_4;
  wire [7:0] t_r3_c42_5;
  wire [7:0] t_r3_c42_6;
  wire [7:0] t_r3_c42_7;
  wire [7:0] t_r3_c42_8;
  wire [7:0] t_r3_c42_9;
  wire [7:0] t_r3_c42_10;
  wire [7:0] t_r3_c42_11;
  wire [7:0] t_r3_c42_12;
  wire [7:0] t_r3_c43_0;
  wire [7:0] t_r3_c43_1;
  wire [7:0] t_r3_c43_2;
  wire [7:0] t_r3_c43_3;
  wire [7:0] t_r3_c43_4;
  wire [7:0] t_r3_c43_5;
  wire [7:0] t_r3_c43_6;
  wire [7:0] t_r3_c43_7;
  wire [7:0] t_r3_c43_8;
  wire [7:0] t_r3_c43_9;
  wire [7:0] t_r3_c43_10;
  wire [7:0] t_r3_c43_11;
  wire [7:0] t_r3_c43_12;
  wire [7:0] t_r3_c44_0;
  wire [7:0] t_r3_c44_1;
  wire [7:0] t_r3_c44_2;
  wire [7:0] t_r3_c44_3;
  wire [7:0] t_r3_c44_4;
  wire [7:0] t_r3_c44_5;
  wire [7:0] t_r3_c44_6;
  wire [7:0] t_r3_c44_7;
  wire [7:0] t_r3_c44_8;
  wire [7:0] t_r3_c44_9;
  wire [7:0] t_r3_c44_10;
  wire [7:0] t_r3_c44_11;
  wire [7:0] t_r3_c44_12;
  wire [7:0] t_r3_c45_0;
  wire [7:0] t_r3_c45_1;
  wire [7:0] t_r3_c45_2;
  wire [7:0] t_r3_c45_3;
  wire [7:0] t_r3_c45_4;
  wire [7:0] t_r3_c45_5;
  wire [7:0] t_r3_c45_6;
  wire [7:0] t_r3_c45_7;
  wire [7:0] t_r3_c45_8;
  wire [7:0] t_r3_c45_9;
  wire [7:0] t_r3_c45_10;
  wire [7:0] t_r3_c45_11;
  wire [7:0] t_r3_c45_12;
  wire [7:0] t_r3_c46_0;
  wire [7:0] t_r3_c46_1;
  wire [7:0] t_r3_c46_2;
  wire [7:0] t_r3_c46_3;
  wire [7:0] t_r3_c46_4;
  wire [7:0] t_r3_c46_5;
  wire [7:0] t_r3_c46_6;
  wire [7:0] t_r3_c46_7;
  wire [7:0] t_r3_c46_8;
  wire [7:0] t_r3_c46_9;
  wire [7:0] t_r3_c46_10;
  wire [7:0] t_r3_c46_11;
  wire [7:0] t_r3_c46_12;
  wire [7:0] t_r3_c47_0;
  wire [7:0] t_r3_c47_1;
  wire [7:0] t_r3_c47_2;
  wire [7:0] t_r3_c47_3;
  wire [7:0] t_r3_c47_4;
  wire [7:0] t_r3_c47_5;
  wire [7:0] t_r3_c47_6;
  wire [7:0] t_r3_c47_7;
  wire [7:0] t_r3_c47_8;
  wire [7:0] t_r3_c47_9;
  wire [7:0] t_r3_c47_10;
  wire [7:0] t_r3_c47_11;
  wire [7:0] t_r3_c47_12;
  wire [7:0] t_r3_c48_0;
  wire [7:0] t_r3_c48_1;
  wire [7:0] t_r3_c48_2;
  wire [7:0] t_r3_c48_3;
  wire [7:0] t_r3_c48_4;
  wire [7:0] t_r3_c48_5;
  wire [7:0] t_r3_c48_6;
  wire [7:0] t_r3_c48_7;
  wire [7:0] t_r3_c48_8;
  wire [7:0] t_r3_c48_9;
  wire [7:0] t_r3_c48_10;
  wire [7:0] t_r3_c48_11;
  wire [7:0] t_r3_c48_12;
  wire [7:0] t_r3_c49_0;
  wire [7:0] t_r3_c49_1;
  wire [7:0] t_r3_c49_2;
  wire [7:0] t_r3_c49_3;
  wire [7:0] t_r3_c49_4;
  wire [7:0] t_r3_c49_5;
  wire [7:0] t_r3_c49_6;
  wire [7:0] t_r3_c49_7;
  wire [7:0] t_r3_c49_8;
  wire [7:0] t_r3_c49_9;
  wire [7:0] t_r3_c49_10;
  wire [7:0] t_r3_c49_11;
  wire [7:0] t_r3_c49_12;
  wire [7:0] t_r3_c50_0;
  wire [7:0] t_r3_c50_1;
  wire [7:0] t_r3_c50_2;
  wire [7:0] t_r3_c50_3;
  wire [7:0] t_r3_c50_4;
  wire [7:0] t_r3_c50_5;
  wire [7:0] t_r3_c50_6;
  wire [7:0] t_r3_c50_7;
  wire [7:0] t_r3_c50_8;
  wire [7:0] t_r3_c50_9;
  wire [7:0] t_r3_c50_10;
  wire [7:0] t_r3_c50_11;
  wire [7:0] t_r3_c50_12;
  wire [7:0] t_r3_c51_0;
  wire [7:0] t_r3_c51_1;
  wire [7:0] t_r3_c51_2;
  wire [7:0] t_r3_c51_3;
  wire [7:0] t_r3_c51_4;
  wire [7:0] t_r3_c51_5;
  wire [7:0] t_r3_c51_6;
  wire [7:0] t_r3_c51_7;
  wire [7:0] t_r3_c51_8;
  wire [7:0] t_r3_c51_9;
  wire [7:0] t_r3_c51_10;
  wire [7:0] t_r3_c51_11;
  wire [7:0] t_r3_c51_12;
  wire [7:0] t_r3_c52_0;
  wire [7:0] t_r3_c52_1;
  wire [7:0] t_r3_c52_2;
  wire [7:0] t_r3_c52_3;
  wire [7:0] t_r3_c52_4;
  wire [7:0] t_r3_c52_5;
  wire [7:0] t_r3_c52_6;
  wire [7:0] t_r3_c52_7;
  wire [7:0] t_r3_c52_8;
  wire [7:0] t_r3_c52_9;
  wire [7:0] t_r3_c52_10;
  wire [7:0] t_r3_c52_11;
  wire [7:0] t_r3_c52_12;
  wire [7:0] t_r3_c53_0;
  wire [7:0] t_r3_c53_1;
  wire [7:0] t_r3_c53_2;
  wire [7:0] t_r3_c53_3;
  wire [7:0] t_r3_c53_4;
  wire [7:0] t_r3_c53_5;
  wire [7:0] t_r3_c53_6;
  wire [7:0] t_r3_c53_7;
  wire [7:0] t_r3_c53_8;
  wire [7:0] t_r3_c53_9;
  wire [7:0] t_r3_c53_10;
  wire [7:0] t_r3_c53_11;
  wire [7:0] t_r3_c53_12;
  wire [7:0] t_r3_c54_0;
  wire [7:0] t_r3_c54_1;
  wire [7:0] t_r3_c54_2;
  wire [7:0] t_r3_c54_3;
  wire [7:0] t_r3_c54_4;
  wire [7:0] t_r3_c54_5;
  wire [7:0] t_r3_c54_6;
  wire [7:0] t_r3_c54_7;
  wire [7:0] t_r3_c54_8;
  wire [7:0] t_r3_c54_9;
  wire [7:0] t_r3_c54_10;
  wire [7:0] t_r3_c54_11;
  wire [7:0] t_r3_c54_12;
  wire [7:0] t_r3_c55_0;
  wire [7:0] t_r3_c55_1;
  wire [7:0] t_r3_c55_2;
  wire [7:0] t_r3_c55_3;
  wire [7:0] t_r3_c55_4;
  wire [7:0] t_r3_c55_5;
  wire [7:0] t_r3_c55_6;
  wire [7:0] t_r3_c55_7;
  wire [7:0] t_r3_c55_8;
  wire [7:0] t_r3_c55_9;
  wire [7:0] t_r3_c55_10;
  wire [7:0] t_r3_c55_11;
  wire [7:0] t_r3_c55_12;
  wire [7:0] t_r3_c56_0;
  wire [7:0] t_r3_c56_1;
  wire [7:0] t_r3_c56_2;
  wire [7:0] t_r3_c56_3;
  wire [7:0] t_r3_c56_4;
  wire [7:0] t_r3_c56_5;
  wire [7:0] t_r3_c56_6;
  wire [7:0] t_r3_c56_7;
  wire [7:0] t_r3_c56_8;
  wire [7:0] t_r3_c56_9;
  wire [7:0] t_r3_c56_10;
  wire [7:0] t_r3_c56_11;
  wire [7:0] t_r3_c56_12;
  wire [7:0] t_r3_c57_0;
  wire [7:0] t_r3_c57_1;
  wire [7:0] t_r3_c57_2;
  wire [7:0] t_r3_c57_3;
  wire [7:0] t_r3_c57_4;
  wire [7:0] t_r3_c57_5;
  wire [7:0] t_r3_c57_6;
  wire [7:0] t_r3_c57_7;
  wire [7:0] t_r3_c57_8;
  wire [7:0] t_r3_c57_9;
  wire [7:0] t_r3_c57_10;
  wire [7:0] t_r3_c57_11;
  wire [7:0] t_r3_c57_12;
  wire [7:0] t_r3_c58_0;
  wire [7:0] t_r3_c58_1;
  wire [7:0] t_r3_c58_2;
  wire [7:0] t_r3_c58_3;
  wire [7:0] t_r3_c58_4;
  wire [7:0] t_r3_c58_5;
  wire [7:0] t_r3_c58_6;
  wire [7:0] t_r3_c58_7;
  wire [7:0] t_r3_c58_8;
  wire [7:0] t_r3_c58_9;
  wire [7:0] t_r3_c58_10;
  wire [7:0] t_r3_c58_11;
  wire [7:0] t_r3_c58_12;
  wire [7:0] t_r3_c59_0;
  wire [7:0] t_r3_c59_1;
  wire [7:0] t_r3_c59_2;
  wire [7:0] t_r3_c59_3;
  wire [7:0] t_r3_c59_4;
  wire [7:0] t_r3_c59_5;
  wire [7:0] t_r3_c59_6;
  wire [7:0] t_r3_c59_7;
  wire [7:0] t_r3_c59_8;
  wire [7:0] t_r3_c59_9;
  wire [7:0] t_r3_c59_10;
  wire [7:0] t_r3_c59_11;
  wire [7:0] t_r3_c59_12;
  wire [7:0] t_r3_c60_0;
  wire [7:0] t_r3_c60_1;
  wire [7:0] t_r3_c60_2;
  wire [7:0] t_r3_c60_3;
  wire [7:0] t_r3_c60_4;
  wire [7:0] t_r3_c60_5;
  wire [7:0] t_r3_c60_6;
  wire [7:0] t_r3_c60_7;
  wire [7:0] t_r3_c60_8;
  wire [7:0] t_r3_c60_9;
  wire [7:0] t_r3_c60_10;
  wire [7:0] t_r3_c60_11;
  wire [7:0] t_r3_c60_12;
  wire [7:0] t_r3_c61_0;
  wire [7:0] t_r3_c61_1;
  wire [7:0] t_r3_c61_2;
  wire [7:0] t_r3_c61_3;
  wire [7:0] t_r3_c61_4;
  wire [7:0] t_r3_c61_5;
  wire [7:0] t_r3_c61_6;
  wire [7:0] t_r3_c61_7;
  wire [7:0] t_r3_c61_8;
  wire [7:0] t_r3_c61_9;
  wire [7:0] t_r3_c61_10;
  wire [7:0] t_r3_c61_11;
  wire [7:0] t_r3_c61_12;
  wire [7:0] t_r3_c62_0;
  wire [7:0] t_r3_c62_1;
  wire [7:0] t_r3_c62_2;
  wire [7:0] t_r3_c62_3;
  wire [7:0] t_r3_c62_4;
  wire [7:0] t_r3_c62_5;
  wire [7:0] t_r3_c62_6;
  wire [7:0] t_r3_c62_7;
  wire [7:0] t_r3_c62_8;
  wire [7:0] t_r3_c62_9;
  wire [7:0] t_r3_c62_10;
  wire [7:0] t_r3_c62_11;
  wire [7:0] t_r3_c62_12;
  wire [7:0] t_r3_c63_0;
  wire [7:0] t_r3_c63_1;
  wire [7:0] t_r3_c63_2;
  wire [7:0] t_r3_c63_3;
  wire [7:0] t_r3_c63_4;
  wire [7:0] t_r3_c63_5;
  wire [7:0] t_r3_c63_6;
  wire [7:0] t_r3_c63_7;
  wire [7:0] t_r3_c63_8;
  wire [7:0] t_r3_c63_9;
  wire [7:0] t_r3_c63_10;
  wire [7:0] t_r3_c63_11;
  wire [7:0] t_r3_c63_12;
  wire [7:0] t_r3_c64_0;
  wire [7:0] t_r3_c64_1;
  wire [7:0] t_r3_c64_2;
  wire [7:0] t_r3_c64_3;
  wire [7:0] t_r3_c64_4;
  wire [7:0] t_r3_c64_5;
  wire [7:0] t_r3_c64_6;
  wire [7:0] t_r3_c64_7;
  wire [7:0] t_r3_c64_8;
  wire [7:0] t_r3_c64_9;
  wire [7:0] t_r3_c64_10;
  wire [7:0] t_r3_c64_11;
  wire [7:0] t_r3_c64_12;
  wire [7:0] t_r3_c65_0;
  wire [7:0] t_r3_c65_1;
  wire [7:0] t_r3_c65_2;
  wire [7:0] t_r3_c65_3;
  wire [7:0] t_r3_c65_4;
  wire [7:0] t_r3_c65_5;
  wire [7:0] t_r3_c65_6;
  wire [7:0] t_r3_c65_7;
  wire [7:0] t_r3_c65_8;
  wire [7:0] t_r3_c65_9;
  wire [7:0] t_r3_c65_10;
  wire [7:0] t_r3_c65_11;
  wire [7:0] t_r3_c65_12;
  wire [7:0] t_r4_c0_0;
  wire [7:0] t_r4_c0_1;
  wire [7:0] t_r4_c0_2;
  wire [7:0] t_r4_c0_3;
  wire [7:0] t_r4_c0_4;
  wire [7:0] t_r4_c0_5;
  wire [7:0] t_r4_c0_6;
  wire [7:0] t_r4_c0_7;
  wire [7:0] t_r4_c0_8;
  wire [7:0] t_r4_c0_9;
  wire [7:0] t_r4_c0_10;
  wire [7:0] t_r4_c0_11;
  wire [7:0] t_r4_c0_12;
  wire [7:0] t_r4_c1_0;
  wire [7:0] t_r4_c1_1;
  wire [7:0] t_r4_c1_2;
  wire [7:0] t_r4_c1_3;
  wire [7:0] t_r4_c1_4;
  wire [7:0] t_r4_c1_5;
  wire [7:0] t_r4_c1_6;
  wire [7:0] t_r4_c1_7;
  wire [7:0] t_r4_c1_8;
  wire [7:0] t_r4_c1_9;
  wire [7:0] t_r4_c1_10;
  wire [7:0] t_r4_c1_11;
  wire [7:0] t_r4_c1_12;
  wire [7:0] t_r4_c2_0;
  wire [7:0] t_r4_c2_1;
  wire [7:0] t_r4_c2_2;
  wire [7:0] t_r4_c2_3;
  wire [7:0] t_r4_c2_4;
  wire [7:0] t_r4_c2_5;
  wire [7:0] t_r4_c2_6;
  wire [7:0] t_r4_c2_7;
  wire [7:0] t_r4_c2_8;
  wire [7:0] t_r4_c2_9;
  wire [7:0] t_r4_c2_10;
  wire [7:0] t_r4_c2_11;
  wire [7:0] t_r4_c2_12;
  wire [7:0] t_r4_c3_0;
  wire [7:0] t_r4_c3_1;
  wire [7:0] t_r4_c3_2;
  wire [7:0] t_r4_c3_3;
  wire [7:0] t_r4_c3_4;
  wire [7:0] t_r4_c3_5;
  wire [7:0] t_r4_c3_6;
  wire [7:0] t_r4_c3_7;
  wire [7:0] t_r4_c3_8;
  wire [7:0] t_r4_c3_9;
  wire [7:0] t_r4_c3_10;
  wire [7:0] t_r4_c3_11;
  wire [7:0] t_r4_c3_12;
  wire [7:0] t_r4_c4_0;
  wire [7:0] t_r4_c4_1;
  wire [7:0] t_r4_c4_2;
  wire [7:0] t_r4_c4_3;
  wire [7:0] t_r4_c4_4;
  wire [7:0] t_r4_c4_5;
  wire [7:0] t_r4_c4_6;
  wire [7:0] t_r4_c4_7;
  wire [7:0] t_r4_c4_8;
  wire [7:0] t_r4_c4_9;
  wire [7:0] t_r4_c4_10;
  wire [7:0] t_r4_c4_11;
  wire [7:0] t_r4_c4_12;
  wire [7:0] t_r4_c5_0;
  wire [7:0] t_r4_c5_1;
  wire [7:0] t_r4_c5_2;
  wire [7:0] t_r4_c5_3;
  wire [7:0] t_r4_c5_4;
  wire [7:0] t_r4_c5_5;
  wire [7:0] t_r4_c5_6;
  wire [7:0] t_r4_c5_7;
  wire [7:0] t_r4_c5_8;
  wire [7:0] t_r4_c5_9;
  wire [7:0] t_r4_c5_10;
  wire [7:0] t_r4_c5_11;
  wire [7:0] t_r4_c5_12;
  wire [7:0] t_r4_c6_0;
  wire [7:0] t_r4_c6_1;
  wire [7:0] t_r4_c6_2;
  wire [7:0] t_r4_c6_3;
  wire [7:0] t_r4_c6_4;
  wire [7:0] t_r4_c6_5;
  wire [7:0] t_r4_c6_6;
  wire [7:0] t_r4_c6_7;
  wire [7:0] t_r4_c6_8;
  wire [7:0] t_r4_c6_9;
  wire [7:0] t_r4_c6_10;
  wire [7:0] t_r4_c6_11;
  wire [7:0] t_r4_c6_12;
  wire [7:0] t_r4_c7_0;
  wire [7:0] t_r4_c7_1;
  wire [7:0] t_r4_c7_2;
  wire [7:0] t_r4_c7_3;
  wire [7:0] t_r4_c7_4;
  wire [7:0] t_r4_c7_5;
  wire [7:0] t_r4_c7_6;
  wire [7:0] t_r4_c7_7;
  wire [7:0] t_r4_c7_8;
  wire [7:0] t_r4_c7_9;
  wire [7:0] t_r4_c7_10;
  wire [7:0] t_r4_c7_11;
  wire [7:0] t_r4_c7_12;
  wire [7:0] t_r4_c8_0;
  wire [7:0] t_r4_c8_1;
  wire [7:0] t_r4_c8_2;
  wire [7:0] t_r4_c8_3;
  wire [7:0] t_r4_c8_4;
  wire [7:0] t_r4_c8_5;
  wire [7:0] t_r4_c8_6;
  wire [7:0] t_r4_c8_7;
  wire [7:0] t_r4_c8_8;
  wire [7:0] t_r4_c8_9;
  wire [7:0] t_r4_c8_10;
  wire [7:0] t_r4_c8_11;
  wire [7:0] t_r4_c8_12;
  wire [7:0] t_r4_c9_0;
  wire [7:0] t_r4_c9_1;
  wire [7:0] t_r4_c9_2;
  wire [7:0] t_r4_c9_3;
  wire [7:0] t_r4_c9_4;
  wire [7:0] t_r4_c9_5;
  wire [7:0] t_r4_c9_6;
  wire [7:0] t_r4_c9_7;
  wire [7:0] t_r4_c9_8;
  wire [7:0] t_r4_c9_9;
  wire [7:0] t_r4_c9_10;
  wire [7:0] t_r4_c9_11;
  wire [7:0] t_r4_c9_12;
  wire [7:0] t_r4_c10_0;
  wire [7:0] t_r4_c10_1;
  wire [7:0] t_r4_c10_2;
  wire [7:0] t_r4_c10_3;
  wire [7:0] t_r4_c10_4;
  wire [7:0] t_r4_c10_5;
  wire [7:0] t_r4_c10_6;
  wire [7:0] t_r4_c10_7;
  wire [7:0] t_r4_c10_8;
  wire [7:0] t_r4_c10_9;
  wire [7:0] t_r4_c10_10;
  wire [7:0] t_r4_c10_11;
  wire [7:0] t_r4_c10_12;
  wire [7:0] t_r4_c11_0;
  wire [7:0] t_r4_c11_1;
  wire [7:0] t_r4_c11_2;
  wire [7:0] t_r4_c11_3;
  wire [7:0] t_r4_c11_4;
  wire [7:0] t_r4_c11_5;
  wire [7:0] t_r4_c11_6;
  wire [7:0] t_r4_c11_7;
  wire [7:0] t_r4_c11_8;
  wire [7:0] t_r4_c11_9;
  wire [7:0] t_r4_c11_10;
  wire [7:0] t_r4_c11_11;
  wire [7:0] t_r4_c11_12;
  wire [7:0] t_r4_c12_0;
  wire [7:0] t_r4_c12_1;
  wire [7:0] t_r4_c12_2;
  wire [7:0] t_r4_c12_3;
  wire [7:0] t_r4_c12_4;
  wire [7:0] t_r4_c12_5;
  wire [7:0] t_r4_c12_6;
  wire [7:0] t_r4_c12_7;
  wire [7:0] t_r4_c12_8;
  wire [7:0] t_r4_c12_9;
  wire [7:0] t_r4_c12_10;
  wire [7:0] t_r4_c12_11;
  wire [7:0] t_r4_c12_12;
  wire [7:0] t_r4_c13_0;
  wire [7:0] t_r4_c13_1;
  wire [7:0] t_r4_c13_2;
  wire [7:0] t_r4_c13_3;
  wire [7:0] t_r4_c13_4;
  wire [7:0] t_r4_c13_5;
  wire [7:0] t_r4_c13_6;
  wire [7:0] t_r4_c13_7;
  wire [7:0] t_r4_c13_8;
  wire [7:0] t_r4_c13_9;
  wire [7:0] t_r4_c13_10;
  wire [7:0] t_r4_c13_11;
  wire [7:0] t_r4_c13_12;
  wire [7:0] t_r4_c14_0;
  wire [7:0] t_r4_c14_1;
  wire [7:0] t_r4_c14_2;
  wire [7:0] t_r4_c14_3;
  wire [7:0] t_r4_c14_4;
  wire [7:0] t_r4_c14_5;
  wire [7:0] t_r4_c14_6;
  wire [7:0] t_r4_c14_7;
  wire [7:0] t_r4_c14_8;
  wire [7:0] t_r4_c14_9;
  wire [7:0] t_r4_c14_10;
  wire [7:0] t_r4_c14_11;
  wire [7:0] t_r4_c14_12;
  wire [7:0] t_r4_c15_0;
  wire [7:0] t_r4_c15_1;
  wire [7:0] t_r4_c15_2;
  wire [7:0] t_r4_c15_3;
  wire [7:0] t_r4_c15_4;
  wire [7:0] t_r4_c15_5;
  wire [7:0] t_r4_c15_6;
  wire [7:0] t_r4_c15_7;
  wire [7:0] t_r4_c15_8;
  wire [7:0] t_r4_c15_9;
  wire [7:0] t_r4_c15_10;
  wire [7:0] t_r4_c15_11;
  wire [7:0] t_r4_c15_12;
  wire [7:0] t_r4_c16_0;
  wire [7:0] t_r4_c16_1;
  wire [7:0] t_r4_c16_2;
  wire [7:0] t_r4_c16_3;
  wire [7:0] t_r4_c16_4;
  wire [7:0] t_r4_c16_5;
  wire [7:0] t_r4_c16_6;
  wire [7:0] t_r4_c16_7;
  wire [7:0] t_r4_c16_8;
  wire [7:0] t_r4_c16_9;
  wire [7:0] t_r4_c16_10;
  wire [7:0] t_r4_c16_11;
  wire [7:0] t_r4_c16_12;
  wire [7:0] t_r4_c17_0;
  wire [7:0] t_r4_c17_1;
  wire [7:0] t_r4_c17_2;
  wire [7:0] t_r4_c17_3;
  wire [7:0] t_r4_c17_4;
  wire [7:0] t_r4_c17_5;
  wire [7:0] t_r4_c17_6;
  wire [7:0] t_r4_c17_7;
  wire [7:0] t_r4_c17_8;
  wire [7:0] t_r4_c17_9;
  wire [7:0] t_r4_c17_10;
  wire [7:0] t_r4_c17_11;
  wire [7:0] t_r4_c17_12;
  wire [7:0] t_r4_c18_0;
  wire [7:0] t_r4_c18_1;
  wire [7:0] t_r4_c18_2;
  wire [7:0] t_r4_c18_3;
  wire [7:0] t_r4_c18_4;
  wire [7:0] t_r4_c18_5;
  wire [7:0] t_r4_c18_6;
  wire [7:0] t_r4_c18_7;
  wire [7:0] t_r4_c18_8;
  wire [7:0] t_r4_c18_9;
  wire [7:0] t_r4_c18_10;
  wire [7:0] t_r4_c18_11;
  wire [7:0] t_r4_c18_12;
  wire [7:0] t_r4_c19_0;
  wire [7:0] t_r4_c19_1;
  wire [7:0] t_r4_c19_2;
  wire [7:0] t_r4_c19_3;
  wire [7:0] t_r4_c19_4;
  wire [7:0] t_r4_c19_5;
  wire [7:0] t_r4_c19_6;
  wire [7:0] t_r4_c19_7;
  wire [7:0] t_r4_c19_8;
  wire [7:0] t_r4_c19_9;
  wire [7:0] t_r4_c19_10;
  wire [7:0] t_r4_c19_11;
  wire [7:0] t_r4_c19_12;
  wire [7:0] t_r4_c20_0;
  wire [7:0] t_r4_c20_1;
  wire [7:0] t_r4_c20_2;
  wire [7:0] t_r4_c20_3;
  wire [7:0] t_r4_c20_4;
  wire [7:0] t_r4_c20_5;
  wire [7:0] t_r4_c20_6;
  wire [7:0] t_r4_c20_7;
  wire [7:0] t_r4_c20_8;
  wire [7:0] t_r4_c20_9;
  wire [7:0] t_r4_c20_10;
  wire [7:0] t_r4_c20_11;
  wire [7:0] t_r4_c20_12;
  wire [7:0] t_r4_c21_0;
  wire [7:0] t_r4_c21_1;
  wire [7:0] t_r4_c21_2;
  wire [7:0] t_r4_c21_3;
  wire [7:0] t_r4_c21_4;
  wire [7:0] t_r4_c21_5;
  wire [7:0] t_r4_c21_6;
  wire [7:0] t_r4_c21_7;
  wire [7:0] t_r4_c21_8;
  wire [7:0] t_r4_c21_9;
  wire [7:0] t_r4_c21_10;
  wire [7:0] t_r4_c21_11;
  wire [7:0] t_r4_c21_12;
  wire [7:0] t_r4_c22_0;
  wire [7:0] t_r4_c22_1;
  wire [7:0] t_r4_c22_2;
  wire [7:0] t_r4_c22_3;
  wire [7:0] t_r4_c22_4;
  wire [7:0] t_r4_c22_5;
  wire [7:0] t_r4_c22_6;
  wire [7:0] t_r4_c22_7;
  wire [7:0] t_r4_c22_8;
  wire [7:0] t_r4_c22_9;
  wire [7:0] t_r4_c22_10;
  wire [7:0] t_r4_c22_11;
  wire [7:0] t_r4_c22_12;
  wire [7:0] t_r4_c23_0;
  wire [7:0] t_r4_c23_1;
  wire [7:0] t_r4_c23_2;
  wire [7:0] t_r4_c23_3;
  wire [7:0] t_r4_c23_4;
  wire [7:0] t_r4_c23_5;
  wire [7:0] t_r4_c23_6;
  wire [7:0] t_r4_c23_7;
  wire [7:0] t_r4_c23_8;
  wire [7:0] t_r4_c23_9;
  wire [7:0] t_r4_c23_10;
  wire [7:0] t_r4_c23_11;
  wire [7:0] t_r4_c23_12;
  wire [7:0] t_r4_c24_0;
  wire [7:0] t_r4_c24_1;
  wire [7:0] t_r4_c24_2;
  wire [7:0] t_r4_c24_3;
  wire [7:0] t_r4_c24_4;
  wire [7:0] t_r4_c24_5;
  wire [7:0] t_r4_c24_6;
  wire [7:0] t_r4_c24_7;
  wire [7:0] t_r4_c24_8;
  wire [7:0] t_r4_c24_9;
  wire [7:0] t_r4_c24_10;
  wire [7:0] t_r4_c24_11;
  wire [7:0] t_r4_c24_12;
  wire [7:0] t_r4_c25_0;
  wire [7:0] t_r4_c25_1;
  wire [7:0] t_r4_c25_2;
  wire [7:0] t_r4_c25_3;
  wire [7:0] t_r4_c25_4;
  wire [7:0] t_r4_c25_5;
  wire [7:0] t_r4_c25_6;
  wire [7:0] t_r4_c25_7;
  wire [7:0] t_r4_c25_8;
  wire [7:0] t_r4_c25_9;
  wire [7:0] t_r4_c25_10;
  wire [7:0] t_r4_c25_11;
  wire [7:0] t_r4_c25_12;
  wire [7:0] t_r4_c26_0;
  wire [7:0] t_r4_c26_1;
  wire [7:0] t_r4_c26_2;
  wire [7:0] t_r4_c26_3;
  wire [7:0] t_r4_c26_4;
  wire [7:0] t_r4_c26_5;
  wire [7:0] t_r4_c26_6;
  wire [7:0] t_r4_c26_7;
  wire [7:0] t_r4_c26_8;
  wire [7:0] t_r4_c26_9;
  wire [7:0] t_r4_c26_10;
  wire [7:0] t_r4_c26_11;
  wire [7:0] t_r4_c26_12;
  wire [7:0] t_r4_c27_0;
  wire [7:0] t_r4_c27_1;
  wire [7:0] t_r4_c27_2;
  wire [7:0] t_r4_c27_3;
  wire [7:0] t_r4_c27_4;
  wire [7:0] t_r4_c27_5;
  wire [7:0] t_r4_c27_6;
  wire [7:0] t_r4_c27_7;
  wire [7:0] t_r4_c27_8;
  wire [7:0] t_r4_c27_9;
  wire [7:0] t_r4_c27_10;
  wire [7:0] t_r4_c27_11;
  wire [7:0] t_r4_c27_12;
  wire [7:0] t_r4_c28_0;
  wire [7:0] t_r4_c28_1;
  wire [7:0] t_r4_c28_2;
  wire [7:0] t_r4_c28_3;
  wire [7:0] t_r4_c28_4;
  wire [7:0] t_r4_c28_5;
  wire [7:0] t_r4_c28_6;
  wire [7:0] t_r4_c28_7;
  wire [7:0] t_r4_c28_8;
  wire [7:0] t_r4_c28_9;
  wire [7:0] t_r4_c28_10;
  wire [7:0] t_r4_c28_11;
  wire [7:0] t_r4_c28_12;
  wire [7:0] t_r4_c29_0;
  wire [7:0] t_r4_c29_1;
  wire [7:0] t_r4_c29_2;
  wire [7:0] t_r4_c29_3;
  wire [7:0] t_r4_c29_4;
  wire [7:0] t_r4_c29_5;
  wire [7:0] t_r4_c29_6;
  wire [7:0] t_r4_c29_7;
  wire [7:0] t_r4_c29_8;
  wire [7:0] t_r4_c29_9;
  wire [7:0] t_r4_c29_10;
  wire [7:0] t_r4_c29_11;
  wire [7:0] t_r4_c29_12;
  wire [7:0] t_r4_c30_0;
  wire [7:0] t_r4_c30_1;
  wire [7:0] t_r4_c30_2;
  wire [7:0] t_r4_c30_3;
  wire [7:0] t_r4_c30_4;
  wire [7:0] t_r4_c30_5;
  wire [7:0] t_r4_c30_6;
  wire [7:0] t_r4_c30_7;
  wire [7:0] t_r4_c30_8;
  wire [7:0] t_r4_c30_9;
  wire [7:0] t_r4_c30_10;
  wire [7:0] t_r4_c30_11;
  wire [7:0] t_r4_c30_12;
  wire [7:0] t_r4_c31_0;
  wire [7:0] t_r4_c31_1;
  wire [7:0] t_r4_c31_2;
  wire [7:0] t_r4_c31_3;
  wire [7:0] t_r4_c31_4;
  wire [7:0] t_r4_c31_5;
  wire [7:0] t_r4_c31_6;
  wire [7:0] t_r4_c31_7;
  wire [7:0] t_r4_c31_8;
  wire [7:0] t_r4_c31_9;
  wire [7:0] t_r4_c31_10;
  wire [7:0] t_r4_c31_11;
  wire [7:0] t_r4_c31_12;
  wire [7:0] t_r4_c32_0;
  wire [7:0] t_r4_c32_1;
  wire [7:0] t_r4_c32_2;
  wire [7:0] t_r4_c32_3;
  wire [7:0] t_r4_c32_4;
  wire [7:0] t_r4_c32_5;
  wire [7:0] t_r4_c32_6;
  wire [7:0] t_r4_c32_7;
  wire [7:0] t_r4_c32_8;
  wire [7:0] t_r4_c32_9;
  wire [7:0] t_r4_c32_10;
  wire [7:0] t_r4_c32_11;
  wire [7:0] t_r4_c32_12;
  wire [7:0] t_r4_c33_0;
  wire [7:0] t_r4_c33_1;
  wire [7:0] t_r4_c33_2;
  wire [7:0] t_r4_c33_3;
  wire [7:0] t_r4_c33_4;
  wire [7:0] t_r4_c33_5;
  wire [7:0] t_r4_c33_6;
  wire [7:0] t_r4_c33_7;
  wire [7:0] t_r4_c33_8;
  wire [7:0] t_r4_c33_9;
  wire [7:0] t_r4_c33_10;
  wire [7:0] t_r4_c33_11;
  wire [7:0] t_r4_c33_12;
  wire [7:0] t_r4_c34_0;
  wire [7:0] t_r4_c34_1;
  wire [7:0] t_r4_c34_2;
  wire [7:0] t_r4_c34_3;
  wire [7:0] t_r4_c34_4;
  wire [7:0] t_r4_c34_5;
  wire [7:0] t_r4_c34_6;
  wire [7:0] t_r4_c34_7;
  wire [7:0] t_r4_c34_8;
  wire [7:0] t_r4_c34_9;
  wire [7:0] t_r4_c34_10;
  wire [7:0] t_r4_c34_11;
  wire [7:0] t_r4_c34_12;
  wire [7:0] t_r4_c35_0;
  wire [7:0] t_r4_c35_1;
  wire [7:0] t_r4_c35_2;
  wire [7:0] t_r4_c35_3;
  wire [7:0] t_r4_c35_4;
  wire [7:0] t_r4_c35_5;
  wire [7:0] t_r4_c35_6;
  wire [7:0] t_r4_c35_7;
  wire [7:0] t_r4_c35_8;
  wire [7:0] t_r4_c35_9;
  wire [7:0] t_r4_c35_10;
  wire [7:0] t_r4_c35_11;
  wire [7:0] t_r4_c35_12;
  wire [7:0] t_r4_c36_0;
  wire [7:0] t_r4_c36_1;
  wire [7:0] t_r4_c36_2;
  wire [7:0] t_r4_c36_3;
  wire [7:0] t_r4_c36_4;
  wire [7:0] t_r4_c36_5;
  wire [7:0] t_r4_c36_6;
  wire [7:0] t_r4_c36_7;
  wire [7:0] t_r4_c36_8;
  wire [7:0] t_r4_c36_9;
  wire [7:0] t_r4_c36_10;
  wire [7:0] t_r4_c36_11;
  wire [7:0] t_r4_c36_12;
  wire [7:0] t_r4_c37_0;
  wire [7:0] t_r4_c37_1;
  wire [7:0] t_r4_c37_2;
  wire [7:0] t_r4_c37_3;
  wire [7:0] t_r4_c37_4;
  wire [7:0] t_r4_c37_5;
  wire [7:0] t_r4_c37_6;
  wire [7:0] t_r4_c37_7;
  wire [7:0] t_r4_c37_8;
  wire [7:0] t_r4_c37_9;
  wire [7:0] t_r4_c37_10;
  wire [7:0] t_r4_c37_11;
  wire [7:0] t_r4_c37_12;
  wire [7:0] t_r4_c38_0;
  wire [7:0] t_r4_c38_1;
  wire [7:0] t_r4_c38_2;
  wire [7:0] t_r4_c38_3;
  wire [7:0] t_r4_c38_4;
  wire [7:0] t_r4_c38_5;
  wire [7:0] t_r4_c38_6;
  wire [7:0] t_r4_c38_7;
  wire [7:0] t_r4_c38_8;
  wire [7:0] t_r4_c38_9;
  wire [7:0] t_r4_c38_10;
  wire [7:0] t_r4_c38_11;
  wire [7:0] t_r4_c38_12;
  wire [7:0] t_r4_c39_0;
  wire [7:0] t_r4_c39_1;
  wire [7:0] t_r4_c39_2;
  wire [7:0] t_r4_c39_3;
  wire [7:0] t_r4_c39_4;
  wire [7:0] t_r4_c39_5;
  wire [7:0] t_r4_c39_6;
  wire [7:0] t_r4_c39_7;
  wire [7:0] t_r4_c39_8;
  wire [7:0] t_r4_c39_9;
  wire [7:0] t_r4_c39_10;
  wire [7:0] t_r4_c39_11;
  wire [7:0] t_r4_c39_12;
  wire [7:0] t_r4_c40_0;
  wire [7:0] t_r4_c40_1;
  wire [7:0] t_r4_c40_2;
  wire [7:0] t_r4_c40_3;
  wire [7:0] t_r4_c40_4;
  wire [7:0] t_r4_c40_5;
  wire [7:0] t_r4_c40_6;
  wire [7:0] t_r4_c40_7;
  wire [7:0] t_r4_c40_8;
  wire [7:0] t_r4_c40_9;
  wire [7:0] t_r4_c40_10;
  wire [7:0] t_r4_c40_11;
  wire [7:0] t_r4_c40_12;
  wire [7:0] t_r4_c41_0;
  wire [7:0] t_r4_c41_1;
  wire [7:0] t_r4_c41_2;
  wire [7:0] t_r4_c41_3;
  wire [7:0] t_r4_c41_4;
  wire [7:0] t_r4_c41_5;
  wire [7:0] t_r4_c41_6;
  wire [7:0] t_r4_c41_7;
  wire [7:0] t_r4_c41_8;
  wire [7:0] t_r4_c41_9;
  wire [7:0] t_r4_c41_10;
  wire [7:0] t_r4_c41_11;
  wire [7:0] t_r4_c41_12;
  wire [7:0] t_r4_c42_0;
  wire [7:0] t_r4_c42_1;
  wire [7:0] t_r4_c42_2;
  wire [7:0] t_r4_c42_3;
  wire [7:0] t_r4_c42_4;
  wire [7:0] t_r4_c42_5;
  wire [7:0] t_r4_c42_6;
  wire [7:0] t_r4_c42_7;
  wire [7:0] t_r4_c42_8;
  wire [7:0] t_r4_c42_9;
  wire [7:0] t_r4_c42_10;
  wire [7:0] t_r4_c42_11;
  wire [7:0] t_r4_c42_12;
  wire [7:0] t_r4_c43_0;
  wire [7:0] t_r4_c43_1;
  wire [7:0] t_r4_c43_2;
  wire [7:0] t_r4_c43_3;
  wire [7:0] t_r4_c43_4;
  wire [7:0] t_r4_c43_5;
  wire [7:0] t_r4_c43_6;
  wire [7:0] t_r4_c43_7;
  wire [7:0] t_r4_c43_8;
  wire [7:0] t_r4_c43_9;
  wire [7:0] t_r4_c43_10;
  wire [7:0] t_r4_c43_11;
  wire [7:0] t_r4_c43_12;
  wire [7:0] t_r4_c44_0;
  wire [7:0] t_r4_c44_1;
  wire [7:0] t_r4_c44_2;
  wire [7:0] t_r4_c44_3;
  wire [7:0] t_r4_c44_4;
  wire [7:0] t_r4_c44_5;
  wire [7:0] t_r4_c44_6;
  wire [7:0] t_r4_c44_7;
  wire [7:0] t_r4_c44_8;
  wire [7:0] t_r4_c44_9;
  wire [7:0] t_r4_c44_10;
  wire [7:0] t_r4_c44_11;
  wire [7:0] t_r4_c44_12;
  wire [7:0] t_r4_c45_0;
  wire [7:0] t_r4_c45_1;
  wire [7:0] t_r4_c45_2;
  wire [7:0] t_r4_c45_3;
  wire [7:0] t_r4_c45_4;
  wire [7:0] t_r4_c45_5;
  wire [7:0] t_r4_c45_6;
  wire [7:0] t_r4_c45_7;
  wire [7:0] t_r4_c45_8;
  wire [7:0] t_r4_c45_9;
  wire [7:0] t_r4_c45_10;
  wire [7:0] t_r4_c45_11;
  wire [7:0] t_r4_c45_12;
  wire [7:0] t_r4_c46_0;
  wire [7:0] t_r4_c46_1;
  wire [7:0] t_r4_c46_2;
  wire [7:0] t_r4_c46_3;
  wire [7:0] t_r4_c46_4;
  wire [7:0] t_r4_c46_5;
  wire [7:0] t_r4_c46_6;
  wire [7:0] t_r4_c46_7;
  wire [7:0] t_r4_c46_8;
  wire [7:0] t_r4_c46_9;
  wire [7:0] t_r4_c46_10;
  wire [7:0] t_r4_c46_11;
  wire [7:0] t_r4_c46_12;
  wire [7:0] t_r4_c47_0;
  wire [7:0] t_r4_c47_1;
  wire [7:0] t_r4_c47_2;
  wire [7:0] t_r4_c47_3;
  wire [7:0] t_r4_c47_4;
  wire [7:0] t_r4_c47_5;
  wire [7:0] t_r4_c47_6;
  wire [7:0] t_r4_c47_7;
  wire [7:0] t_r4_c47_8;
  wire [7:0] t_r4_c47_9;
  wire [7:0] t_r4_c47_10;
  wire [7:0] t_r4_c47_11;
  wire [7:0] t_r4_c47_12;
  wire [7:0] t_r4_c48_0;
  wire [7:0] t_r4_c48_1;
  wire [7:0] t_r4_c48_2;
  wire [7:0] t_r4_c48_3;
  wire [7:0] t_r4_c48_4;
  wire [7:0] t_r4_c48_5;
  wire [7:0] t_r4_c48_6;
  wire [7:0] t_r4_c48_7;
  wire [7:0] t_r4_c48_8;
  wire [7:0] t_r4_c48_9;
  wire [7:0] t_r4_c48_10;
  wire [7:0] t_r4_c48_11;
  wire [7:0] t_r4_c48_12;
  wire [7:0] t_r4_c49_0;
  wire [7:0] t_r4_c49_1;
  wire [7:0] t_r4_c49_2;
  wire [7:0] t_r4_c49_3;
  wire [7:0] t_r4_c49_4;
  wire [7:0] t_r4_c49_5;
  wire [7:0] t_r4_c49_6;
  wire [7:0] t_r4_c49_7;
  wire [7:0] t_r4_c49_8;
  wire [7:0] t_r4_c49_9;
  wire [7:0] t_r4_c49_10;
  wire [7:0] t_r4_c49_11;
  wire [7:0] t_r4_c49_12;
  wire [7:0] t_r4_c50_0;
  wire [7:0] t_r4_c50_1;
  wire [7:0] t_r4_c50_2;
  wire [7:0] t_r4_c50_3;
  wire [7:0] t_r4_c50_4;
  wire [7:0] t_r4_c50_5;
  wire [7:0] t_r4_c50_6;
  wire [7:0] t_r4_c50_7;
  wire [7:0] t_r4_c50_8;
  wire [7:0] t_r4_c50_9;
  wire [7:0] t_r4_c50_10;
  wire [7:0] t_r4_c50_11;
  wire [7:0] t_r4_c50_12;
  wire [7:0] t_r4_c51_0;
  wire [7:0] t_r4_c51_1;
  wire [7:0] t_r4_c51_2;
  wire [7:0] t_r4_c51_3;
  wire [7:0] t_r4_c51_4;
  wire [7:0] t_r4_c51_5;
  wire [7:0] t_r4_c51_6;
  wire [7:0] t_r4_c51_7;
  wire [7:0] t_r4_c51_8;
  wire [7:0] t_r4_c51_9;
  wire [7:0] t_r4_c51_10;
  wire [7:0] t_r4_c51_11;
  wire [7:0] t_r4_c51_12;
  wire [7:0] t_r4_c52_0;
  wire [7:0] t_r4_c52_1;
  wire [7:0] t_r4_c52_2;
  wire [7:0] t_r4_c52_3;
  wire [7:0] t_r4_c52_4;
  wire [7:0] t_r4_c52_5;
  wire [7:0] t_r4_c52_6;
  wire [7:0] t_r4_c52_7;
  wire [7:0] t_r4_c52_8;
  wire [7:0] t_r4_c52_9;
  wire [7:0] t_r4_c52_10;
  wire [7:0] t_r4_c52_11;
  wire [7:0] t_r4_c52_12;
  wire [7:0] t_r4_c53_0;
  wire [7:0] t_r4_c53_1;
  wire [7:0] t_r4_c53_2;
  wire [7:0] t_r4_c53_3;
  wire [7:0] t_r4_c53_4;
  wire [7:0] t_r4_c53_5;
  wire [7:0] t_r4_c53_6;
  wire [7:0] t_r4_c53_7;
  wire [7:0] t_r4_c53_8;
  wire [7:0] t_r4_c53_9;
  wire [7:0] t_r4_c53_10;
  wire [7:0] t_r4_c53_11;
  wire [7:0] t_r4_c53_12;
  wire [7:0] t_r4_c54_0;
  wire [7:0] t_r4_c54_1;
  wire [7:0] t_r4_c54_2;
  wire [7:0] t_r4_c54_3;
  wire [7:0] t_r4_c54_4;
  wire [7:0] t_r4_c54_5;
  wire [7:0] t_r4_c54_6;
  wire [7:0] t_r4_c54_7;
  wire [7:0] t_r4_c54_8;
  wire [7:0] t_r4_c54_9;
  wire [7:0] t_r4_c54_10;
  wire [7:0] t_r4_c54_11;
  wire [7:0] t_r4_c54_12;
  wire [7:0] t_r4_c55_0;
  wire [7:0] t_r4_c55_1;
  wire [7:0] t_r4_c55_2;
  wire [7:0] t_r4_c55_3;
  wire [7:0] t_r4_c55_4;
  wire [7:0] t_r4_c55_5;
  wire [7:0] t_r4_c55_6;
  wire [7:0] t_r4_c55_7;
  wire [7:0] t_r4_c55_8;
  wire [7:0] t_r4_c55_9;
  wire [7:0] t_r4_c55_10;
  wire [7:0] t_r4_c55_11;
  wire [7:0] t_r4_c55_12;
  wire [7:0] t_r4_c56_0;
  wire [7:0] t_r4_c56_1;
  wire [7:0] t_r4_c56_2;
  wire [7:0] t_r4_c56_3;
  wire [7:0] t_r4_c56_4;
  wire [7:0] t_r4_c56_5;
  wire [7:0] t_r4_c56_6;
  wire [7:0] t_r4_c56_7;
  wire [7:0] t_r4_c56_8;
  wire [7:0] t_r4_c56_9;
  wire [7:0] t_r4_c56_10;
  wire [7:0] t_r4_c56_11;
  wire [7:0] t_r4_c56_12;
  wire [7:0] t_r4_c57_0;
  wire [7:0] t_r4_c57_1;
  wire [7:0] t_r4_c57_2;
  wire [7:0] t_r4_c57_3;
  wire [7:0] t_r4_c57_4;
  wire [7:0] t_r4_c57_5;
  wire [7:0] t_r4_c57_6;
  wire [7:0] t_r4_c57_7;
  wire [7:0] t_r4_c57_8;
  wire [7:0] t_r4_c57_9;
  wire [7:0] t_r4_c57_10;
  wire [7:0] t_r4_c57_11;
  wire [7:0] t_r4_c57_12;
  wire [7:0] t_r4_c58_0;
  wire [7:0] t_r4_c58_1;
  wire [7:0] t_r4_c58_2;
  wire [7:0] t_r4_c58_3;
  wire [7:0] t_r4_c58_4;
  wire [7:0] t_r4_c58_5;
  wire [7:0] t_r4_c58_6;
  wire [7:0] t_r4_c58_7;
  wire [7:0] t_r4_c58_8;
  wire [7:0] t_r4_c58_9;
  wire [7:0] t_r4_c58_10;
  wire [7:0] t_r4_c58_11;
  wire [7:0] t_r4_c58_12;
  wire [7:0] t_r4_c59_0;
  wire [7:0] t_r4_c59_1;
  wire [7:0] t_r4_c59_2;
  wire [7:0] t_r4_c59_3;
  wire [7:0] t_r4_c59_4;
  wire [7:0] t_r4_c59_5;
  wire [7:0] t_r4_c59_6;
  wire [7:0] t_r4_c59_7;
  wire [7:0] t_r4_c59_8;
  wire [7:0] t_r4_c59_9;
  wire [7:0] t_r4_c59_10;
  wire [7:0] t_r4_c59_11;
  wire [7:0] t_r4_c59_12;
  wire [7:0] t_r4_c60_0;
  wire [7:0] t_r4_c60_1;
  wire [7:0] t_r4_c60_2;
  wire [7:0] t_r4_c60_3;
  wire [7:0] t_r4_c60_4;
  wire [7:0] t_r4_c60_5;
  wire [7:0] t_r4_c60_6;
  wire [7:0] t_r4_c60_7;
  wire [7:0] t_r4_c60_8;
  wire [7:0] t_r4_c60_9;
  wire [7:0] t_r4_c60_10;
  wire [7:0] t_r4_c60_11;
  wire [7:0] t_r4_c60_12;
  wire [7:0] t_r4_c61_0;
  wire [7:0] t_r4_c61_1;
  wire [7:0] t_r4_c61_2;
  wire [7:0] t_r4_c61_3;
  wire [7:0] t_r4_c61_4;
  wire [7:0] t_r4_c61_5;
  wire [7:0] t_r4_c61_6;
  wire [7:0] t_r4_c61_7;
  wire [7:0] t_r4_c61_8;
  wire [7:0] t_r4_c61_9;
  wire [7:0] t_r4_c61_10;
  wire [7:0] t_r4_c61_11;
  wire [7:0] t_r4_c61_12;
  wire [7:0] t_r4_c62_0;
  wire [7:0] t_r4_c62_1;
  wire [7:0] t_r4_c62_2;
  wire [7:0] t_r4_c62_3;
  wire [7:0] t_r4_c62_4;
  wire [7:0] t_r4_c62_5;
  wire [7:0] t_r4_c62_6;
  wire [7:0] t_r4_c62_7;
  wire [7:0] t_r4_c62_8;
  wire [7:0] t_r4_c62_9;
  wire [7:0] t_r4_c62_10;
  wire [7:0] t_r4_c62_11;
  wire [7:0] t_r4_c62_12;
  wire [7:0] t_r4_c63_0;
  wire [7:0] t_r4_c63_1;
  wire [7:0] t_r4_c63_2;
  wire [7:0] t_r4_c63_3;
  wire [7:0] t_r4_c63_4;
  wire [7:0] t_r4_c63_5;
  wire [7:0] t_r4_c63_6;
  wire [7:0] t_r4_c63_7;
  wire [7:0] t_r4_c63_8;
  wire [7:0] t_r4_c63_9;
  wire [7:0] t_r4_c63_10;
  wire [7:0] t_r4_c63_11;
  wire [7:0] t_r4_c63_12;
  wire [7:0] t_r4_c64_0;
  wire [7:0] t_r4_c64_1;
  wire [7:0] t_r4_c64_2;
  wire [7:0] t_r4_c64_3;
  wire [7:0] t_r4_c64_4;
  wire [7:0] t_r4_c64_5;
  wire [7:0] t_r4_c64_6;
  wire [7:0] t_r4_c64_7;
  wire [7:0] t_r4_c64_8;
  wire [7:0] t_r4_c64_9;
  wire [7:0] t_r4_c64_10;
  wire [7:0] t_r4_c64_11;
  wire [7:0] t_r4_c64_12;
  wire [7:0] t_r4_c65_0;
  wire [7:0] t_r4_c65_1;
  wire [7:0] t_r4_c65_2;
  wire [7:0] t_r4_c65_3;
  wire [7:0] t_r4_c65_4;
  wire [7:0] t_r4_c65_5;
  wire [7:0] t_r4_c65_6;
  wire [7:0] t_r4_c65_7;
  wire [7:0] t_r4_c65_8;
  wire [7:0] t_r4_c65_9;
  wire [7:0] t_r4_c65_10;
  wire [7:0] t_r4_c65_11;
  wire [7:0] t_r4_c65_12;
  wire [7:0] t_r5_c0_0;
  wire [7:0] t_r5_c0_1;
  wire [7:0] t_r5_c0_2;
  wire [7:0] t_r5_c0_3;
  wire [7:0] t_r5_c0_4;
  wire [7:0] t_r5_c0_5;
  wire [7:0] t_r5_c0_6;
  wire [7:0] t_r5_c0_7;
  wire [7:0] t_r5_c0_8;
  wire [7:0] t_r5_c0_9;
  wire [7:0] t_r5_c0_10;
  wire [7:0] t_r5_c0_11;
  wire [7:0] t_r5_c0_12;
  wire [7:0] t_r5_c1_0;
  wire [7:0] t_r5_c1_1;
  wire [7:0] t_r5_c1_2;
  wire [7:0] t_r5_c1_3;
  wire [7:0] t_r5_c1_4;
  wire [7:0] t_r5_c1_5;
  wire [7:0] t_r5_c1_6;
  wire [7:0] t_r5_c1_7;
  wire [7:0] t_r5_c1_8;
  wire [7:0] t_r5_c1_9;
  wire [7:0] t_r5_c1_10;
  wire [7:0] t_r5_c1_11;
  wire [7:0] t_r5_c1_12;
  wire [7:0] t_r5_c2_0;
  wire [7:0] t_r5_c2_1;
  wire [7:0] t_r5_c2_2;
  wire [7:0] t_r5_c2_3;
  wire [7:0] t_r5_c2_4;
  wire [7:0] t_r5_c2_5;
  wire [7:0] t_r5_c2_6;
  wire [7:0] t_r5_c2_7;
  wire [7:0] t_r5_c2_8;
  wire [7:0] t_r5_c2_9;
  wire [7:0] t_r5_c2_10;
  wire [7:0] t_r5_c2_11;
  wire [7:0] t_r5_c2_12;
  wire [7:0] t_r5_c3_0;
  wire [7:0] t_r5_c3_1;
  wire [7:0] t_r5_c3_2;
  wire [7:0] t_r5_c3_3;
  wire [7:0] t_r5_c3_4;
  wire [7:0] t_r5_c3_5;
  wire [7:0] t_r5_c3_6;
  wire [7:0] t_r5_c3_7;
  wire [7:0] t_r5_c3_8;
  wire [7:0] t_r5_c3_9;
  wire [7:0] t_r5_c3_10;
  wire [7:0] t_r5_c3_11;
  wire [7:0] t_r5_c3_12;
  wire [7:0] t_r5_c4_0;
  wire [7:0] t_r5_c4_1;
  wire [7:0] t_r5_c4_2;
  wire [7:0] t_r5_c4_3;
  wire [7:0] t_r5_c4_4;
  wire [7:0] t_r5_c4_5;
  wire [7:0] t_r5_c4_6;
  wire [7:0] t_r5_c4_7;
  wire [7:0] t_r5_c4_8;
  wire [7:0] t_r5_c4_9;
  wire [7:0] t_r5_c4_10;
  wire [7:0] t_r5_c4_11;
  wire [7:0] t_r5_c4_12;
  wire [7:0] t_r5_c5_0;
  wire [7:0] t_r5_c5_1;
  wire [7:0] t_r5_c5_2;
  wire [7:0] t_r5_c5_3;
  wire [7:0] t_r5_c5_4;
  wire [7:0] t_r5_c5_5;
  wire [7:0] t_r5_c5_6;
  wire [7:0] t_r5_c5_7;
  wire [7:0] t_r5_c5_8;
  wire [7:0] t_r5_c5_9;
  wire [7:0] t_r5_c5_10;
  wire [7:0] t_r5_c5_11;
  wire [7:0] t_r5_c5_12;
  wire [7:0] t_r5_c6_0;
  wire [7:0] t_r5_c6_1;
  wire [7:0] t_r5_c6_2;
  wire [7:0] t_r5_c6_3;
  wire [7:0] t_r5_c6_4;
  wire [7:0] t_r5_c6_5;
  wire [7:0] t_r5_c6_6;
  wire [7:0] t_r5_c6_7;
  wire [7:0] t_r5_c6_8;
  wire [7:0] t_r5_c6_9;
  wire [7:0] t_r5_c6_10;
  wire [7:0] t_r5_c6_11;
  wire [7:0] t_r5_c6_12;
  wire [7:0] t_r5_c7_0;
  wire [7:0] t_r5_c7_1;
  wire [7:0] t_r5_c7_2;
  wire [7:0] t_r5_c7_3;
  wire [7:0] t_r5_c7_4;
  wire [7:0] t_r5_c7_5;
  wire [7:0] t_r5_c7_6;
  wire [7:0] t_r5_c7_7;
  wire [7:0] t_r5_c7_8;
  wire [7:0] t_r5_c7_9;
  wire [7:0] t_r5_c7_10;
  wire [7:0] t_r5_c7_11;
  wire [7:0] t_r5_c7_12;
  wire [7:0] t_r5_c8_0;
  wire [7:0] t_r5_c8_1;
  wire [7:0] t_r5_c8_2;
  wire [7:0] t_r5_c8_3;
  wire [7:0] t_r5_c8_4;
  wire [7:0] t_r5_c8_5;
  wire [7:0] t_r5_c8_6;
  wire [7:0] t_r5_c8_7;
  wire [7:0] t_r5_c8_8;
  wire [7:0] t_r5_c8_9;
  wire [7:0] t_r5_c8_10;
  wire [7:0] t_r5_c8_11;
  wire [7:0] t_r5_c8_12;
  wire [7:0] t_r5_c9_0;
  wire [7:0] t_r5_c9_1;
  wire [7:0] t_r5_c9_2;
  wire [7:0] t_r5_c9_3;
  wire [7:0] t_r5_c9_4;
  wire [7:0] t_r5_c9_5;
  wire [7:0] t_r5_c9_6;
  wire [7:0] t_r5_c9_7;
  wire [7:0] t_r5_c9_8;
  wire [7:0] t_r5_c9_9;
  wire [7:0] t_r5_c9_10;
  wire [7:0] t_r5_c9_11;
  wire [7:0] t_r5_c9_12;
  wire [7:0] t_r5_c10_0;
  wire [7:0] t_r5_c10_1;
  wire [7:0] t_r5_c10_2;
  wire [7:0] t_r5_c10_3;
  wire [7:0] t_r5_c10_4;
  wire [7:0] t_r5_c10_5;
  wire [7:0] t_r5_c10_6;
  wire [7:0] t_r5_c10_7;
  wire [7:0] t_r5_c10_8;
  wire [7:0] t_r5_c10_9;
  wire [7:0] t_r5_c10_10;
  wire [7:0] t_r5_c10_11;
  wire [7:0] t_r5_c10_12;
  wire [7:0] t_r5_c11_0;
  wire [7:0] t_r5_c11_1;
  wire [7:0] t_r5_c11_2;
  wire [7:0] t_r5_c11_3;
  wire [7:0] t_r5_c11_4;
  wire [7:0] t_r5_c11_5;
  wire [7:0] t_r5_c11_6;
  wire [7:0] t_r5_c11_7;
  wire [7:0] t_r5_c11_8;
  wire [7:0] t_r5_c11_9;
  wire [7:0] t_r5_c11_10;
  wire [7:0] t_r5_c11_11;
  wire [7:0] t_r5_c11_12;
  wire [7:0] t_r5_c12_0;
  wire [7:0] t_r5_c12_1;
  wire [7:0] t_r5_c12_2;
  wire [7:0] t_r5_c12_3;
  wire [7:0] t_r5_c12_4;
  wire [7:0] t_r5_c12_5;
  wire [7:0] t_r5_c12_6;
  wire [7:0] t_r5_c12_7;
  wire [7:0] t_r5_c12_8;
  wire [7:0] t_r5_c12_9;
  wire [7:0] t_r5_c12_10;
  wire [7:0] t_r5_c12_11;
  wire [7:0] t_r5_c12_12;
  wire [7:0] t_r5_c13_0;
  wire [7:0] t_r5_c13_1;
  wire [7:0] t_r5_c13_2;
  wire [7:0] t_r5_c13_3;
  wire [7:0] t_r5_c13_4;
  wire [7:0] t_r5_c13_5;
  wire [7:0] t_r5_c13_6;
  wire [7:0] t_r5_c13_7;
  wire [7:0] t_r5_c13_8;
  wire [7:0] t_r5_c13_9;
  wire [7:0] t_r5_c13_10;
  wire [7:0] t_r5_c13_11;
  wire [7:0] t_r5_c13_12;
  wire [7:0] t_r5_c14_0;
  wire [7:0] t_r5_c14_1;
  wire [7:0] t_r5_c14_2;
  wire [7:0] t_r5_c14_3;
  wire [7:0] t_r5_c14_4;
  wire [7:0] t_r5_c14_5;
  wire [7:0] t_r5_c14_6;
  wire [7:0] t_r5_c14_7;
  wire [7:0] t_r5_c14_8;
  wire [7:0] t_r5_c14_9;
  wire [7:0] t_r5_c14_10;
  wire [7:0] t_r5_c14_11;
  wire [7:0] t_r5_c14_12;
  wire [7:0] t_r5_c15_0;
  wire [7:0] t_r5_c15_1;
  wire [7:0] t_r5_c15_2;
  wire [7:0] t_r5_c15_3;
  wire [7:0] t_r5_c15_4;
  wire [7:0] t_r5_c15_5;
  wire [7:0] t_r5_c15_6;
  wire [7:0] t_r5_c15_7;
  wire [7:0] t_r5_c15_8;
  wire [7:0] t_r5_c15_9;
  wire [7:0] t_r5_c15_10;
  wire [7:0] t_r5_c15_11;
  wire [7:0] t_r5_c15_12;
  wire [7:0] t_r5_c16_0;
  wire [7:0] t_r5_c16_1;
  wire [7:0] t_r5_c16_2;
  wire [7:0] t_r5_c16_3;
  wire [7:0] t_r5_c16_4;
  wire [7:0] t_r5_c16_5;
  wire [7:0] t_r5_c16_6;
  wire [7:0] t_r5_c16_7;
  wire [7:0] t_r5_c16_8;
  wire [7:0] t_r5_c16_9;
  wire [7:0] t_r5_c16_10;
  wire [7:0] t_r5_c16_11;
  wire [7:0] t_r5_c16_12;
  wire [7:0] t_r5_c17_0;
  wire [7:0] t_r5_c17_1;
  wire [7:0] t_r5_c17_2;
  wire [7:0] t_r5_c17_3;
  wire [7:0] t_r5_c17_4;
  wire [7:0] t_r5_c17_5;
  wire [7:0] t_r5_c17_6;
  wire [7:0] t_r5_c17_7;
  wire [7:0] t_r5_c17_8;
  wire [7:0] t_r5_c17_9;
  wire [7:0] t_r5_c17_10;
  wire [7:0] t_r5_c17_11;
  wire [7:0] t_r5_c17_12;
  wire [7:0] t_r5_c18_0;
  wire [7:0] t_r5_c18_1;
  wire [7:0] t_r5_c18_2;
  wire [7:0] t_r5_c18_3;
  wire [7:0] t_r5_c18_4;
  wire [7:0] t_r5_c18_5;
  wire [7:0] t_r5_c18_6;
  wire [7:0] t_r5_c18_7;
  wire [7:0] t_r5_c18_8;
  wire [7:0] t_r5_c18_9;
  wire [7:0] t_r5_c18_10;
  wire [7:0] t_r5_c18_11;
  wire [7:0] t_r5_c18_12;
  wire [7:0] t_r5_c19_0;
  wire [7:0] t_r5_c19_1;
  wire [7:0] t_r5_c19_2;
  wire [7:0] t_r5_c19_3;
  wire [7:0] t_r5_c19_4;
  wire [7:0] t_r5_c19_5;
  wire [7:0] t_r5_c19_6;
  wire [7:0] t_r5_c19_7;
  wire [7:0] t_r5_c19_8;
  wire [7:0] t_r5_c19_9;
  wire [7:0] t_r5_c19_10;
  wire [7:0] t_r5_c19_11;
  wire [7:0] t_r5_c19_12;
  wire [7:0] t_r5_c20_0;
  wire [7:0] t_r5_c20_1;
  wire [7:0] t_r5_c20_2;
  wire [7:0] t_r5_c20_3;
  wire [7:0] t_r5_c20_4;
  wire [7:0] t_r5_c20_5;
  wire [7:0] t_r5_c20_6;
  wire [7:0] t_r5_c20_7;
  wire [7:0] t_r5_c20_8;
  wire [7:0] t_r5_c20_9;
  wire [7:0] t_r5_c20_10;
  wire [7:0] t_r5_c20_11;
  wire [7:0] t_r5_c20_12;
  wire [7:0] t_r5_c21_0;
  wire [7:0] t_r5_c21_1;
  wire [7:0] t_r5_c21_2;
  wire [7:0] t_r5_c21_3;
  wire [7:0] t_r5_c21_4;
  wire [7:0] t_r5_c21_5;
  wire [7:0] t_r5_c21_6;
  wire [7:0] t_r5_c21_7;
  wire [7:0] t_r5_c21_8;
  wire [7:0] t_r5_c21_9;
  wire [7:0] t_r5_c21_10;
  wire [7:0] t_r5_c21_11;
  wire [7:0] t_r5_c21_12;
  wire [7:0] t_r5_c22_0;
  wire [7:0] t_r5_c22_1;
  wire [7:0] t_r5_c22_2;
  wire [7:0] t_r5_c22_3;
  wire [7:0] t_r5_c22_4;
  wire [7:0] t_r5_c22_5;
  wire [7:0] t_r5_c22_6;
  wire [7:0] t_r5_c22_7;
  wire [7:0] t_r5_c22_8;
  wire [7:0] t_r5_c22_9;
  wire [7:0] t_r5_c22_10;
  wire [7:0] t_r5_c22_11;
  wire [7:0] t_r5_c22_12;
  wire [7:0] t_r5_c23_0;
  wire [7:0] t_r5_c23_1;
  wire [7:0] t_r5_c23_2;
  wire [7:0] t_r5_c23_3;
  wire [7:0] t_r5_c23_4;
  wire [7:0] t_r5_c23_5;
  wire [7:0] t_r5_c23_6;
  wire [7:0] t_r5_c23_7;
  wire [7:0] t_r5_c23_8;
  wire [7:0] t_r5_c23_9;
  wire [7:0] t_r5_c23_10;
  wire [7:0] t_r5_c23_11;
  wire [7:0] t_r5_c23_12;
  wire [7:0] t_r5_c24_0;
  wire [7:0] t_r5_c24_1;
  wire [7:0] t_r5_c24_2;
  wire [7:0] t_r5_c24_3;
  wire [7:0] t_r5_c24_4;
  wire [7:0] t_r5_c24_5;
  wire [7:0] t_r5_c24_6;
  wire [7:0] t_r5_c24_7;
  wire [7:0] t_r5_c24_8;
  wire [7:0] t_r5_c24_9;
  wire [7:0] t_r5_c24_10;
  wire [7:0] t_r5_c24_11;
  wire [7:0] t_r5_c24_12;
  wire [7:0] t_r5_c25_0;
  wire [7:0] t_r5_c25_1;
  wire [7:0] t_r5_c25_2;
  wire [7:0] t_r5_c25_3;
  wire [7:0] t_r5_c25_4;
  wire [7:0] t_r5_c25_5;
  wire [7:0] t_r5_c25_6;
  wire [7:0] t_r5_c25_7;
  wire [7:0] t_r5_c25_8;
  wire [7:0] t_r5_c25_9;
  wire [7:0] t_r5_c25_10;
  wire [7:0] t_r5_c25_11;
  wire [7:0] t_r5_c25_12;
  wire [7:0] t_r5_c26_0;
  wire [7:0] t_r5_c26_1;
  wire [7:0] t_r5_c26_2;
  wire [7:0] t_r5_c26_3;
  wire [7:0] t_r5_c26_4;
  wire [7:0] t_r5_c26_5;
  wire [7:0] t_r5_c26_6;
  wire [7:0] t_r5_c26_7;
  wire [7:0] t_r5_c26_8;
  wire [7:0] t_r5_c26_9;
  wire [7:0] t_r5_c26_10;
  wire [7:0] t_r5_c26_11;
  wire [7:0] t_r5_c26_12;
  wire [7:0] t_r5_c27_0;
  wire [7:0] t_r5_c27_1;
  wire [7:0] t_r5_c27_2;
  wire [7:0] t_r5_c27_3;
  wire [7:0] t_r5_c27_4;
  wire [7:0] t_r5_c27_5;
  wire [7:0] t_r5_c27_6;
  wire [7:0] t_r5_c27_7;
  wire [7:0] t_r5_c27_8;
  wire [7:0] t_r5_c27_9;
  wire [7:0] t_r5_c27_10;
  wire [7:0] t_r5_c27_11;
  wire [7:0] t_r5_c27_12;
  wire [7:0] t_r5_c28_0;
  wire [7:0] t_r5_c28_1;
  wire [7:0] t_r5_c28_2;
  wire [7:0] t_r5_c28_3;
  wire [7:0] t_r5_c28_4;
  wire [7:0] t_r5_c28_5;
  wire [7:0] t_r5_c28_6;
  wire [7:0] t_r5_c28_7;
  wire [7:0] t_r5_c28_8;
  wire [7:0] t_r5_c28_9;
  wire [7:0] t_r5_c28_10;
  wire [7:0] t_r5_c28_11;
  wire [7:0] t_r5_c28_12;
  wire [7:0] t_r5_c29_0;
  wire [7:0] t_r5_c29_1;
  wire [7:0] t_r5_c29_2;
  wire [7:0] t_r5_c29_3;
  wire [7:0] t_r5_c29_4;
  wire [7:0] t_r5_c29_5;
  wire [7:0] t_r5_c29_6;
  wire [7:0] t_r5_c29_7;
  wire [7:0] t_r5_c29_8;
  wire [7:0] t_r5_c29_9;
  wire [7:0] t_r5_c29_10;
  wire [7:0] t_r5_c29_11;
  wire [7:0] t_r5_c29_12;
  wire [7:0] t_r5_c30_0;
  wire [7:0] t_r5_c30_1;
  wire [7:0] t_r5_c30_2;
  wire [7:0] t_r5_c30_3;
  wire [7:0] t_r5_c30_4;
  wire [7:0] t_r5_c30_5;
  wire [7:0] t_r5_c30_6;
  wire [7:0] t_r5_c30_7;
  wire [7:0] t_r5_c30_8;
  wire [7:0] t_r5_c30_9;
  wire [7:0] t_r5_c30_10;
  wire [7:0] t_r5_c30_11;
  wire [7:0] t_r5_c30_12;
  wire [7:0] t_r5_c31_0;
  wire [7:0] t_r5_c31_1;
  wire [7:0] t_r5_c31_2;
  wire [7:0] t_r5_c31_3;
  wire [7:0] t_r5_c31_4;
  wire [7:0] t_r5_c31_5;
  wire [7:0] t_r5_c31_6;
  wire [7:0] t_r5_c31_7;
  wire [7:0] t_r5_c31_8;
  wire [7:0] t_r5_c31_9;
  wire [7:0] t_r5_c31_10;
  wire [7:0] t_r5_c31_11;
  wire [7:0] t_r5_c31_12;
  wire [7:0] t_r5_c32_0;
  wire [7:0] t_r5_c32_1;
  wire [7:0] t_r5_c32_2;
  wire [7:0] t_r5_c32_3;
  wire [7:0] t_r5_c32_4;
  wire [7:0] t_r5_c32_5;
  wire [7:0] t_r5_c32_6;
  wire [7:0] t_r5_c32_7;
  wire [7:0] t_r5_c32_8;
  wire [7:0] t_r5_c32_9;
  wire [7:0] t_r5_c32_10;
  wire [7:0] t_r5_c32_11;
  wire [7:0] t_r5_c32_12;
  wire [7:0] t_r5_c33_0;
  wire [7:0] t_r5_c33_1;
  wire [7:0] t_r5_c33_2;
  wire [7:0] t_r5_c33_3;
  wire [7:0] t_r5_c33_4;
  wire [7:0] t_r5_c33_5;
  wire [7:0] t_r5_c33_6;
  wire [7:0] t_r5_c33_7;
  wire [7:0] t_r5_c33_8;
  wire [7:0] t_r5_c33_9;
  wire [7:0] t_r5_c33_10;
  wire [7:0] t_r5_c33_11;
  wire [7:0] t_r5_c33_12;
  wire [7:0] t_r5_c34_0;
  wire [7:0] t_r5_c34_1;
  wire [7:0] t_r5_c34_2;
  wire [7:0] t_r5_c34_3;
  wire [7:0] t_r5_c34_4;
  wire [7:0] t_r5_c34_5;
  wire [7:0] t_r5_c34_6;
  wire [7:0] t_r5_c34_7;
  wire [7:0] t_r5_c34_8;
  wire [7:0] t_r5_c34_9;
  wire [7:0] t_r5_c34_10;
  wire [7:0] t_r5_c34_11;
  wire [7:0] t_r5_c34_12;
  wire [7:0] t_r5_c35_0;
  wire [7:0] t_r5_c35_1;
  wire [7:0] t_r5_c35_2;
  wire [7:0] t_r5_c35_3;
  wire [7:0] t_r5_c35_4;
  wire [7:0] t_r5_c35_5;
  wire [7:0] t_r5_c35_6;
  wire [7:0] t_r5_c35_7;
  wire [7:0] t_r5_c35_8;
  wire [7:0] t_r5_c35_9;
  wire [7:0] t_r5_c35_10;
  wire [7:0] t_r5_c35_11;
  wire [7:0] t_r5_c35_12;
  wire [7:0] t_r5_c36_0;
  wire [7:0] t_r5_c36_1;
  wire [7:0] t_r5_c36_2;
  wire [7:0] t_r5_c36_3;
  wire [7:0] t_r5_c36_4;
  wire [7:0] t_r5_c36_5;
  wire [7:0] t_r5_c36_6;
  wire [7:0] t_r5_c36_7;
  wire [7:0] t_r5_c36_8;
  wire [7:0] t_r5_c36_9;
  wire [7:0] t_r5_c36_10;
  wire [7:0] t_r5_c36_11;
  wire [7:0] t_r5_c36_12;
  wire [7:0] t_r5_c37_0;
  wire [7:0] t_r5_c37_1;
  wire [7:0] t_r5_c37_2;
  wire [7:0] t_r5_c37_3;
  wire [7:0] t_r5_c37_4;
  wire [7:0] t_r5_c37_5;
  wire [7:0] t_r5_c37_6;
  wire [7:0] t_r5_c37_7;
  wire [7:0] t_r5_c37_8;
  wire [7:0] t_r5_c37_9;
  wire [7:0] t_r5_c37_10;
  wire [7:0] t_r5_c37_11;
  wire [7:0] t_r5_c37_12;
  wire [7:0] t_r5_c38_0;
  wire [7:0] t_r5_c38_1;
  wire [7:0] t_r5_c38_2;
  wire [7:0] t_r5_c38_3;
  wire [7:0] t_r5_c38_4;
  wire [7:0] t_r5_c38_5;
  wire [7:0] t_r5_c38_6;
  wire [7:0] t_r5_c38_7;
  wire [7:0] t_r5_c38_8;
  wire [7:0] t_r5_c38_9;
  wire [7:0] t_r5_c38_10;
  wire [7:0] t_r5_c38_11;
  wire [7:0] t_r5_c38_12;
  wire [7:0] t_r5_c39_0;
  wire [7:0] t_r5_c39_1;
  wire [7:0] t_r5_c39_2;
  wire [7:0] t_r5_c39_3;
  wire [7:0] t_r5_c39_4;
  wire [7:0] t_r5_c39_5;
  wire [7:0] t_r5_c39_6;
  wire [7:0] t_r5_c39_7;
  wire [7:0] t_r5_c39_8;
  wire [7:0] t_r5_c39_9;
  wire [7:0] t_r5_c39_10;
  wire [7:0] t_r5_c39_11;
  wire [7:0] t_r5_c39_12;
  wire [7:0] t_r5_c40_0;
  wire [7:0] t_r5_c40_1;
  wire [7:0] t_r5_c40_2;
  wire [7:0] t_r5_c40_3;
  wire [7:0] t_r5_c40_4;
  wire [7:0] t_r5_c40_5;
  wire [7:0] t_r5_c40_6;
  wire [7:0] t_r5_c40_7;
  wire [7:0] t_r5_c40_8;
  wire [7:0] t_r5_c40_9;
  wire [7:0] t_r5_c40_10;
  wire [7:0] t_r5_c40_11;
  wire [7:0] t_r5_c40_12;
  wire [7:0] t_r5_c41_0;
  wire [7:0] t_r5_c41_1;
  wire [7:0] t_r5_c41_2;
  wire [7:0] t_r5_c41_3;
  wire [7:0] t_r5_c41_4;
  wire [7:0] t_r5_c41_5;
  wire [7:0] t_r5_c41_6;
  wire [7:0] t_r5_c41_7;
  wire [7:0] t_r5_c41_8;
  wire [7:0] t_r5_c41_9;
  wire [7:0] t_r5_c41_10;
  wire [7:0] t_r5_c41_11;
  wire [7:0] t_r5_c41_12;
  wire [7:0] t_r5_c42_0;
  wire [7:0] t_r5_c42_1;
  wire [7:0] t_r5_c42_2;
  wire [7:0] t_r5_c42_3;
  wire [7:0] t_r5_c42_4;
  wire [7:0] t_r5_c42_5;
  wire [7:0] t_r5_c42_6;
  wire [7:0] t_r5_c42_7;
  wire [7:0] t_r5_c42_8;
  wire [7:0] t_r5_c42_9;
  wire [7:0] t_r5_c42_10;
  wire [7:0] t_r5_c42_11;
  wire [7:0] t_r5_c42_12;
  wire [7:0] t_r5_c43_0;
  wire [7:0] t_r5_c43_1;
  wire [7:0] t_r5_c43_2;
  wire [7:0] t_r5_c43_3;
  wire [7:0] t_r5_c43_4;
  wire [7:0] t_r5_c43_5;
  wire [7:0] t_r5_c43_6;
  wire [7:0] t_r5_c43_7;
  wire [7:0] t_r5_c43_8;
  wire [7:0] t_r5_c43_9;
  wire [7:0] t_r5_c43_10;
  wire [7:0] t_r5_c43_11;
  wire [7:0] t_r5_c43_12;
  wire [7:0] t_r5_c44_0;
  wire [7:0] t_r5_c44_1;
  wire [7:0] t_r5_c44_2;
  wire [7:0] t_r5_c44_3;
  wire [7:0] t_r5_c44_4;
  wire [7:0] t_r5_c44_5;
  wire [7:0] t_r5_c44_6;
  wire [7:0] t_r5_c44_7;
  wire [7:0] t_r5_c44_8;
  wire [7:0] t_r5_c44_9;
  wire [7:0] t_r5_c44_10;
  wire [7:0] t_r5_c44_11;
  wire [7:0] t_r5_c44_12;
  wire [7:0] t_r5_c45_0;
  wire [7:0] t_r5_c45_1;
  wire [7:0] t_r5_c45_2;
  wire [7:0] t_r5_c45_3;
  wire [7:0] t_r5_c45_4;
  wire [7:0] t_r5_c45_5;
  wire [7:0] t_r5_c45_6;
  wire [7:0] t_r5_c45_7;
  wire [7:0] t_r5_c45_8;
  wire [7:0] t_r5_c45_9;
  wire [7:0] t_r5_c45_10;
  wire [7:0] t_r5_c45_11;
  wire [7:0] t_r5_c45_12;
  wire [7:0] t_r5_c46_0;
  wire [7:0] t_r5_c46_1;
  wire [7:0] t_r5_c46_2;
  wire [7:0] t_r5_c46_3;
  wire [7:0] t_r5_c46_4;
  wire [7:0] t_r5_c46_5;
  wire [7:0] t_r5_c46_6;
  wire [7:0] t_r5_c46_7;
  wire [7:0] t_r5_c46_8;
  wire [7:0] t_r5_c46_9;
  wire [7:0] t_r5_c46_10;
  wire [7:0] t_r5_c46_11;
  wire [7:0] t_r5_c46_12;
  wire [7:0] t_r5_c47_0;
  wire [7:0] t_r5_c47_1;
  wire [7:0] t_r5_c47_2;
  wire [7:0] t_r5_c47_3;
  wire [7:0] t_r5_c47_4;
  wire [7:0] t_r5_c47_5;
  wire [7:0] t_r5_c47_6;
  wire [7:0] t_r5_c47_7;
  wire [7:0] t_r5_c47_8;
  wire [7:0] t_r5_c47_9;
  wire [7:0] t_r5_c47_10;
  wire [7:0] t_r5_c47_11;
  wire [7:0] t_r5_c47_12;
  wire [7:0] t_r5_c48_0;
  wire [7:0] t_r5_c48_1;
  wire [7:0] t_r5_c48_2;
  wire [7:0] t_r5_c48_3;
  wire [7:0] t_r5_c48_4;
  wire [7:0] t_r5_c48_5;
  wire [7:0] t_r5_c48_6;
  wire [7:0] t_r5_c48_7;
  wire [7:0] t_r5_c48_8;
  wire [7:0] t_r5_c48_9;
  wire [7:0] t_r5_c48_10;
  wire [7:0] t_r5_c48_11;
  wire [7:0] t_r5_c48_12;
  wire [7:0] t_r5_c49_0;
  wire [7:0] t_r5_c49_1;
  wire [7:0] t_r5_c49_2;
  wire [7:0] t_r5_c49_3;
  wire [7:0] t_r5_c49_4;
  wire [7:0] t_r5_c49_5;
  wire [7:0] t_r5_c49_6;
  wire [7:0] t_r5_c49_7;
  wire [7:0] t_r5_c49_8;
  wire [7:0] t_r5_c49_9;
  wire [7:0] t_r5_c49_10;
  wire [7:0] t_r5_c49_11;
  wire [7:0] t_r5_c49_12;
  wire [7:0] t_r5_c50_0;
  wire [7:0] t_r5_c50_1;
  wire [7:0] t_r5_c50_2;
  wire [7:0] t_r5_c50_3;
  wire [7:0] t_r5_c50_4;
  wire [7:0] t_r5_c50_5;
  wire [7:0] t_r5_c50_6;
  wire [7:0] t_r5_c50_7;
  wire [7:0] t_r5_c50_8;
  wire [7:0] t_r5_c50_9;
  wire [7:0] t_r5_c50_10;
  wire [7:0] t_r5_c50_11;
  wire [7:0] t_r5_c50_12;
  wire [7:0] t_r5_c51_0;
  wire [7:0] t_r5_c51_1;
  wire [7:0] t_r5_c51_2;
  wire [7:0] t_r5_c51_3;
  wire [7:0] t_r5_c51_4;
  wire [7:0] t_r5_c51_5;
  wire [7:0] t_r5_c51_6;
  wire [7:0] t_r5_c51_7;
  wire [7:0] t_r5_c51_8;
  wire [7:0] t_r5_c51_9;
  wire [7:0] t_r5_c51_10;
  wire [7:0] t_r5_c51_11;
  wire [7:0] t_r5_c51_12;
  wire [7:0] t_r5_c52_0;
  wire [7:0] t_r5_c52_1;
  wire [7:0] t_r5_c52_2;
  wire [7:0] t_r5_c52_3;
  wire [7:0] t_r5_c52_4;
  wire [7:0] t_r5_c52_5;
  wire [7:0] t_r5_c52_6;
  wire [7:0] t_r5_c52_7;
  wire [7:0] t_r5_c52_8;
  wire [7:0] t_r5_c52_9;
  wire [7:0] t_r5_c52_10;
  wire [7:0] t_r5_c52_11;
  wire [7:0] t_r5_c52_12;
  wire [7:0] t_r5_c53_0;
  wire [7:0] t_r5_c53_1;
  wire [7:0] t_r5_c53_2;
  wire [7:0] t_r5_c53_3;
  wire [7:0] t_r5_c53_4;
  wire [7:0] t_r5_c53_5;
  wire [7:0] t_r5_c53_6;
  wire [7:0] t_r5_c53_7;
  wire [7:0] t_r5_c53_8;
  wire [7:0] t_r5_c53_9;
  wire [7:0] t_r5_c53_10;
  wire [7:0] t_r5_c53_11;
  wire [7:0] t_r5_c53_12;
  wire [7:0] t_r5_c54_0;
  wire [7:0] t_r5_c54_1;
  wire [7:0] t_r5_c54_2;
  wire [7:0] t_r5_c54_3;
  wire [7:0] t_r5_c54_4;
  wire [7:0] t_r5_c54_5;
  wire [7:0] t_r5_c54_6;
  wire [7:0] t_r5_c54_7;
  wire [7:0] t_r5_c54_8;
  wire [7:0] t_r5_c54_9;
  wire [7:0] t_r5_c54_10;
  wire [7:0] t_r5_c54_11;
  wire [7:0] t_r5_c54_12;
  wire [7:0] t_r5_c55_0;
  wire [7:0] t_r5_c55_1;
  wire [7:0] t_r5_c55_2;
  wire [7:0] t_r5_c55_3;
  wire [7:0] t_r5_c55_4;
  wire [7:0] t_r5_c55_5;
  wire [7:0] t_r5_c55_6;
  wire [7:0] t_r5_c55_7;
  wire [7:0] t_r5_c55_8;
  wire [7:0] t_r5_c55_9;
  wire [7:0] t_r5_c55_10;
  wire [7:0] t_r5_c55_11;
  wire [7:0] t_r5_c55_12;
  wire [7:0] t_r5_c56_0;
  wire [7:0] t_r5_c56_1;
  wire [7:0] t_r5_c56_2;
  wire [7:0] t_r5_c56_3;
  wire [7:0] t_r5_c56_4;
  wire [7:0] t_r5_c56_5;
  wire [7:0] t_r5_c56_6;
  wire [7:0] t_r5_c56_7;
  wire [7:0] t_r5_c56_8;
  wire [7:0] t_r5_c56_9;
  wire [7:0] t_r5_c56_10;
  wire [7:0] t_r5_c56_11;
  wire [7:0] t_r5_c56_12;
  wire [7:0] t_r5_c57_0;
  wire [7:0] t_r5_c57_1;
  wire [7:0] t_r5_c57_2;
  wire [7:0] t_r5_c57_3;
  wire [7:0] t_r5_c57_4;
  wire [7:0] t_r5_c57_5;
  wire [7:0] t_r5_c57_6;
  wire [7:0] t_r5_c57_7;
  wire [7:0] t_r5_c57_8;
  wire [7:0] t_r5_c57_9;
  wire [7:0] t_r5_c57_10;
  wire [7:0] t_r5_c57_11;
  wire [7:0] t_r5_c57_12;
  wire [7:0] t_r5_c58_0;
  wire [7:0] t_r5_c58_1;
  wire [7:0] t_r5_c58_2;
  wire [7:0] t_r5_c58_3;
  wire [7:0] t_r5_c58_4;
  wire [7:0] t_r5_c58_5;
  wire [7:0] t_r5_c58_6;
  wire [7:0] t_r5_c58_7;
  wire [7:0] t_r5_c58_8;
  wire [7:0] t_r5_c58_9;
  wire [7:0] t_r5_c58_10;
  wire [7:0] t_r5_c58_11;
  wire [7:0] t_r5_c58_12;
  wire [7:0] t_r5_c59_0;
  wire [7:0] t_r5_c59_1;
  wire [7:0] t_r5_c59_2;
  wire [7:0] t_r5_c59_3;
  wire [7:0] t_r5_c59_4;
  wire [7:0] t_r5_c59_5;
  wire [7:0] t_r5_c59_6;
  wire [7:0] t_r5_c59_7;
  wire [7:0] t_r5_c59_8;
  wire [7:0] t_r5_c59_9;
  wire [7:0] t_r5_c59_10;
  wire [7:0] t_r5_c59_11;
  wire [7:0] t_r5_c59_12;
  wire [7:0] t_r5_c60_0;
  wire [7:0] t_r5_c60_1;
  wire [7:0] t_r5_c60_2;
  wire [7:0] t_r5_c60_3;
  wire [7:0] t_r5_c60_4;
  wire [7:0] t_r5_c60_5;
  wire [7:0] t_r5_c60_6;
  wire [7:0] t_r5_c60_7;
  wire [7:0] t_r5_c60_8;
  wire [7:0] t_r5_c60_9;
  wire [7:0] t_r5_c60_10;
  wire [7:0] t_r5_c60_11;
  wire [7:0] t_r5_c60_12;
  wire [7:0] t_r5_c61_0;
  wire [7:0] t_r5_c61_1;
  wire [7:0] t_r5_c61_2;
  wire [7:0] t_r5_c61_3;
  wire [7:0] t_r5_c61_4;
  wire [7:0] t_r5_c61_5;
  wire [7:0] t_r5_c61_6;
  wire [7:0] t_r5_c61_7;
  wire [7:0] t_r5_c61_8;
  wire [7:0] t_r5_c61_9;
  wire [7:0] t_r5_c61_10;
  wire [7:0] t_r5_c61_11;
  wire [7:0] t_r5_c61_12;
  wire [7:0] t_r5_c62_0;
  wire [7:0] t_r5_c62_1;
  wire [7:0] t_r5_c62_2;
  wire [7:0] t_r5_c62_3;
  wire [7:0] t_r5_c62_4;
  wire [7:0] t_r5_c62_5;
  wire [7:0] t_r5_c62_6;
  wire [7:0] t_r5_c62_7;
  wire [7:0] t_r5_c62_8;
  wire [7:0] t_r5_c62_9;
  wire [7:0] t_r5_c62_10;
  wire [7:0] t_r5_c62_11;
  wire [7:0] t_r5_c62_12;
  wire [7:0] t_r5_c63_0;
  wire [7:0] t_r5_c63_1;
  wire [7:0] t_r5_c63_2;
  wire [7:0] t_r5_c63_3;
  wire [7:0] t_r5_c63_4;
  wire [7:0] t_r5_c63_5;
  wire [7:0] t_r5_c63_6;
  wire [7:0] t_r5_c63_7;
  wire [7:0] t_r5_c63_8;
  wire [7:0] t_r5_c63_9;
  wire [7:0] t_r5_c63_10;
  wire [7:0] t_r5_c63_11;
  wire [7:0] t_r5_c63_12;
  wire [7:0] t_r5_c64_0;
  wire [7:0] t_r5_c64_1;
  wire [7:0] t_r5_c64_2;
  wire [7:0] t_r5_c64_3;
  wire [7:0] t_r5_c64_4;
  wire [7:0] t_r5_c64_5;
  wire [7:0] t_r5_c64_6;
  wire [7:0] t_r5_c64_7;
  wire [7:0] t_r5_c64_8;
  wire [7:0] t_r5_c64_9;
  wire [7:0] t_r5_c64_10;
  wire [7:0] t_r5_c64_11;
  wire [7:0] t_r5_c64_12;
  wire [7:0] t_r5_c65_0;
  wire [7:0] t_r5_c65_1;
  wire [7:0] t_r5_c65_2;
  wire [7:0] t_r5_c65_3;
  wire [7:0] t_r5_c65_4;
  wire [7:0] t_r5_c65_5;
  wire [7:0] t_r5_c65_6;
  wire [7:0] t_r5_c65_7;
  wire [7:0] t_r5_c65_8;
  wire [7:0] t_r5_c65_9;
  wire [7:0] t_r5_c65_10;
  wire [7:0] t_r5_c65_11;
  wire [7:0] t_r5_c65_12;
  wire [7:0] t_r6_c0_0;
  wire [7:0] t_r6_c0_1;
  wire [7:0] t_r6_c0_2;
  wire [7:0] t_r6_c0_3;
  wire [7:0] t_r6_c0_4;
  wire [7:0] t_r6_c0_5;
  wire [7:0] t_r6_c0_6;
  wire [7:0] t_r6_c0_7;
  wire [7:0] t_r6_c0_8;
  wire [7:0] t_r6_c0_9;
  wire [7:0] t_r6_c0_10;
  wire [7:0] t_r6_c0_11;
  wire [7:0] t_r6_c0_12;
  wire [7:0] t_r6_c1_0;
  wire [7:0] t_r6_c1_1;
  wire [7:0] t_r6_c1_2;
  wire [7:0] t_r6_c1_3;
  wire [7:0] t_r6_c1_4;
  wire [7:0] t_r6_c1_5;
  wire [7:0] t_r6_c1_6;
  wire [7:0] t_r6_c1_7;
  wire [7:0] t_r6_c1_8;
  wire [7:0] t_r6_c1_9;
  wire [7:0] t_r6_c1_10;
  wire [7:0] t_r6_c1_11;
  wire [7:0] t_r6_c1_12;
  wire [7:0] t_r6_c2_0;
  wire [7:0] t_r6_c2_1;
  wire [7:0] t_r6_c2_2;
  wire [7:0] t_r6_c2_3;
  wire [7:0] t_r6_c2_4;
  wire [7:0] t_r6_c2_5;
  wire [7:0] t_r6_c2_6;
  wire [7:0] t_r6_c2_7;
  wire [7:0] t_r6_c2_8;
  wire [7:0] t_r6_c2_9;
  wire [7:0] t_r6_c2_10;
  wire [7:0] t_r6_c2_11;
  wire [7:0] t_r6_c2_12;
  wire [7:0] t_r6_c3_0;
  wire [7:0] t_r6_c3_1;
  wire [7:0] t_r6_c3_2;
  wire [7:0] t_r6_c3_3;
  wire [7:0] t_r6_c3_4;
  wire [7:0] t_r6_c3_5;
  wire [7:0] t_r6_c3_6;
  wire [7:0] t_r6_c3_7;
  wire [7:0] t_r6_c3_8;
  wire [7:0] t_r6_c3_9;
  wire [7:0] t_r6_c3_10;
  wire [7:0] t_r6_c3_11;
  wire [7:0] t_r6_c3_12;
  wire [7:0] t_r6_c4_0;
  wire [7:0] t_r6_c4_1;
  wire [7:0] t_r6_c4_2;
  wire [7:0] t_r6_c4_3;
  wire [7:0] t_r6_c4_4;
  wire [7:0] t_r6_c4_5;
  wire [7:0] t_r6_c4_6;
  wire [7:0] t_r6_c4_7;
  wire [7:0] t_r6_c4_8;
  wire [7:0] t_r6_c4_9;
  wire [7:0] t_r6_c4_10;
  wire [7:0] t_r6_c4_11;
  wire [7:0] t_r6_c4_12;
  wire [7:0] t_r6_c5_0;
  wire [7:0] t_r6_c5_1;
  wire [7:0] t_r6_c5_2;
  wire [7:0] t_r6_c5_3;
  wire [7:0] t_r6_c5_4;
  wire [7:0] t_r6_c5_5;
  wire [7:0] t_r6_c5_6;
  wire [7:0] t_r6_c5_7;
  wire [7:0] t_r6_c5_8;
  wire [7:0] t_r6_c5_9;
  wire [7:0] t_r6_c5_10;
  wire [7:0] t_r6_c5_11;
  wire [7:0] t_r6_c5_12;
  wire [7:0] t_r6_c6_0;
  wire [7:0] t_r6_c6_1;
  wire [7:0] t_r6_c6_2;
  wire [7:0] t_r6_c6_3;
  wire [7:0] t_r6_c6_4;
  wire [7:0] t_r6_c6_5;
  wire [7:0] t_r6_c6_6;
  wire [7:0] t_r6_c6_7;
  wire [7:0] t_r6_c6_8;
  wire [7:0] t_r6_c6_9;
  wire [7:0] t_r6_c6_10;
  wire [7:0] t_r6_c6_11;
  wire [7:0] t_r6_c6_12;
  wire [7:0] t_r6_c7_0;
  wire [7:0] t_r6_c7_1;
  wire [7:0] t_r6_c7_2;
  wire [7:0] t_r6_c7_3;
  wire [7:0] t_r6_c7_4;
  wire [7:0] t_r6_c7_5;
  wire [7:0] t_r6_c7_6;
  wire [7:0] t_r6_c7_7;
  wire [7:0] t_r6_c7_8;
  wire [7:0] t_r6_c7_9;
  wire [7:0] t_r6_c7_10;
  wire [7:0] t_r6_c7_11;
  wire [7:0] t_r6_c7_12;
  wire [7:0] t_r6_c8_0;
  wire [7:0] t_r6_c8_1;
  wire [7:0] t_r6_c8_2;
  wire [7:0] t_r6_c8_3;
  wire [7:0] t_r6_c8_4;
  wire [7:0] t_r6_c8_5;
  wire [7:0] t_r6_c8_6;
  wire [7:0] t_r6_c8_7;
  wire [7:0] t_r6_c8_8;
  wire [7:0] t_r6_c8_9;
  wire [7:0] t_r6_c8_10;
  wire [7:0] t_r6_c8_11;
  wire [7:0] t_r6_c8_12;
  wire [7:0] t_r6_c9_0;
  wire [7:0] t_r6_c9_1;
  wire [7:0] t_r6_c9_2;
  wire [7:0] t_r6_c9_3;
  wire [7:0] t_r6_c9_4;
  wire [7:0] t_r6_c9_5;
  wire [7:0] t_r6_c9_6;
  wire [7:0] t_r6_c9_7;
  wire [7:0] t_r6_c9_8;
  wire [7:0] t_r6_c9_9;
  wire [7:0] t_r6_c9_10;
  wire [7:0] t_r6_c9_11;
  wire [7:0] t_r6_c9_12;
  wire [7:0] t_r6_c10_0;
  wire [7:0] t_r6_c10_1;
  wire [7:0] t_r6_c10_2;
  wire [7:0] t_r6_c10_3;
  wire [7:0] t_r6_c10_4;
  wire [7:0] t_r6_c10_5;
  wire [7:0] t_r6_c10_6;
  wire [7:0] t_r6_c10_7;
  wire [7:0] t_r6_c10_8;
  wire [7:0] t_r6_c10_9;
  wire [7:0] t_r6_c10_10;
  wire [7:0] t_r6_c10_11;
  wire [7:0] t_r6_c10_12;
  wire [7:0] t_r6_c11_0;
  wire [7:0] t_r6_c11_1;
  wire [7:0] t_r6_c11_2;
  wire [7:0] t_r6_c11_3;
  wire [7:0] t_r6_c11_4;
  wire [7:0] t_r6_c11_5;
  wire [7:0] t_r6_c11_6;
  wire [7:0] t_r6_c11_7;
  wire [7:0] t_r6_c11_8;
  wire [7:0] t_r6_c11_9;
  wire [7:0] t_r6_c11_10;
  wire [7:0] t_r6_c11_11;
  wire [7:0] t_r6_c11_12;
  wire [7:0] t_r6_c12_0;
  wire [7:0] t_r6_c12_1;
  wire [7:0] t_r6_c12_2;
  wire [7:0] t_r6_c12_3;
  wire [7:0] t_r6_c12_4;
  wire [7:0] t_r6_c12_5;
  wire [7:0] t_r6_c12_6;
  wire [7:0] t_r6_c12_7;
  wire [7:0] t_r6_c12_8;
  wire [7:0] t_r6_c12_9;
  wire [7:0] t_r6_c12_10;
  wire [7:0] t_r6_c12_11;
  wire [7:0] t_r6_c12_12;
  wire [7:0] t_r6_c13_0;
  wire [7:0] t_r6_c13_1;
  wire [7:0] t_r6_c13_2;
  wire [7:0] t_r6_c13_3;
  wire [7:0] t_r6_c13_4;
  wire [7:0] t_r6_c13_5;
  wire [7:0] t_r6_c13_6;
  wire [7:0] t_r6_c13_7;
  wire [7:0] t_r6_c13_8;
  wire [7:0] t_r6_c13_9;
  wire [7:0] t_r6_c13_10;
  wire [7:0] t_r6_c13_11;
  wire [7:0] t_r6_c13_12;
  wire [7:0] t_r6_c14_0;
  wire [7:0] t_r6_c14_1;
  wire [7:0] t_r6_c14_2;
  wire [7:0] t_r6_c14_3;
  wire [7:0] t_r6_c14_4;
  wire [7:0] t_r6_c14_5;
  wire [7:0] t_r6_c14_6;
  wire [7:0] t_r6_c14_7;
  wire [7:0] t_r6_c14_8;
  wire [7:0] t_r6_c14_9;
  wire [7:0] t_r6_c14_10;
  wire [7:0] t_r6_c14_11;
  wire [7:0] t_r6_c14_12;
  wire [7:0] t_r6_c15_0;
  wire [7:0] t_r6_c15_1;
  wire [7:0] t_r6_c15_2;
  wire [7:0] t_r6_c15_3;
  wire [7:0] t_r6_c15_4;
  wire [7:0] t_r6_c15_5;
  wire [7:0] t_r6_c15_6;
  wire [7:0] t_r6_c15_7;
  wire [7:0] t_r6_c15_8;
  wire [7:0] t_r6_c15_9;
  wire [7:0] t_r6_c15_10;
  wire [7:0] t_r6_c15_11;
  wire [7:0] t_r6_c15_12;
  wire [7:0] t_r6_c16_0;
  wire [7:0] t_r6_c16_1;
  wire [7:0] t_r6_c16_2;
  wire [7:0] t_r6_c16_3;
  wire [7:0] t_r6_c16_4;
  wire [7:0] t_r6_c16_5;
  wire [7:0] t_r6_c16_6;
  wire [7:0] t_r6_c16_7;
  wire [7:0] t_r6_c16_8;
  wire [7:0] t_r6_c16_9;
  wire [7:0] t_r6_c16_10;
  wire [7:0] t_r6_c16_11;
  wire [7:0] t_r6_c16_12;
  wire [7:0] t_r6_c17_0;
  wire [7:0] t_r6_c17_1;
  wire [7:0] t_r6_c17_2;
  wire [7:0] t_r6_c17_3;
  wire [7:0] t_r6_c17_4;
  wire [7:0] t_r6_c17_5;
  wire [7:0] t_r6_c17_6;
  wire [7:0] t_r6_c17_7;
  wire [7:0] t_r6_c17_8;
  wire [7:0] t_r6_c17_9;
  wire [7:0] t_r6_c17_10;
  wire [7:0] t_r6_c17_11;
  wire [7:0] t_r6_c17_12;
  wire [7:0] t_r6_c18_0;
  wire [7:0] t_r6_c18_1;
  wire [7:0] t_r6_c18_2;
  wire [7:0] t_r6_c18_3;
  wire [7:0] t_r6_c18_4;
  wire [7:0] t_r6_c18_5;
  wire [7:0] t_r6_c18_6;
  wire [7:0] t_r6_c18_7;
  wire [7:0] t_r6_c18_8;
  wire [7:0] t_r6_c18_9;
  wire [7:0] t_r6_c18_10;
  wire [7:0] t_r6_c18_11;
  wire [7:0] t_r6_c18_12;
  wire [7:0] t_r6_c19_0;
  wire [7:0] t_r6_c19_1;
  wire [7:0] t_r6_c19_2;
  wire [7:0] t_r6_c19_3;
  wire [7:0] t_r6_c19_4;
  wire [7:0] t_r6_c19_5;
  wire [7:0] t_r6_c19_6;
  wire [7:0] t_r6_c19_7;
  wire [7:0] t_r6_c19_8;
  wire [7:0] t_r6_c19_9;
  wire [7:0] t_r6_c19_10;
  wire [7:0] t_r6_c19_11;
  wire [7:0] t_r6_c19_12;
  wire [7:0] t_r6_c20_0;
  wire [7:0] t_r6_c20_1;
  wire [7:0] t_r6_c20_2;
  wire [7:0] t_r6_c20_3;
  wire [7:0] t_r6_c20_4;
  wire [7:0] t_r6_c20_5;
  wire [7:0] t_r6_c20_6;
  wire [7:0] t_r6_c20_7;
  wire [7:0] t_r6_c20_8;
  wire [7:0] t_r6_c20_9;
  wire [7:0] t_r6_c20_10;
  wire [7:0] t_r6_c20_11;
  wire [7:0] t_r6_c20_12;
  wire [7:0] t_r6_c21_0;
  wire [7:0] t_r6_c21_1;
  wire [7:0] t_r6_c21_2;
  wire [7:0] t_r6_c21_3;
  wire [7:0] t_r6_c21_4;
  wire [7:0] t_r6_c21_5;
  wire [7:0] t_r6_c21_6;
  wire [7:0] t_r6_c21_7;
  wire [7:0] t_r6_c21_8;
  wire [7:0] t_r6_c21_9;
  wire [7:0] t_r6_c21_10;
  wire [7:0] t_r6_c21_11;
  wire [7:0] t_r6_c21_12;
  wire [7:0] t_r6_c22_0;
  wire [7:0] t_r6_c22_1;
  wire [7:0] t_r6_c22_2;
  wire [7:0] t_r6_c22_3;
  wire [7:0] t_r6_c22_4;
  wire [7:0] t_r6_c22_5;
  wire [7:0] t_r6_c22_6;
  wire [7:0] t_r6_c22_7;
  wire [7:0] t_r6_c22_8;
  wire [7:0] t_r6_c22_9;
  wire [7:0] t_r6_c22_10;
  wire [7:0] t_r6_c22_11;
  wire [7:0] t_r6_c22_12;
  wire [7:0] t_r6_c23_0;
  wire [7:0] t_r6_c23_1;
  wire [7:0] t_r6_c23_2;
  wire [7:0] t_r6_c23_3;
  wire [7:0] t_r6_c23_4;
  wire [7:0] t_r6_c23_5;
  wire [7:0] t_r6_c23_6;
  wire [7:0] t_r6_c23_7;
  wire [7:0] t_r6_c23_8;
  wire [7:0] t_r6_c23_9;
  wire [7:0] t_r6_c23_10;
  wire [7:0] t_r6_c23_11;
  wire [7:0] t_r6_c23_12;
  wire [7:0] t_r6_c24_0;
  wire [7:0] t_r6_c24_1;
  wire [7:0] t_r6_c24_2;
  wire [7:0] t_r6_c24_3;
  wire [7:0] t_r6_c24_4;
  wire [7:0] t_r6_c24_5;
  wire [7:0] t_r6_c24_6;
  wire [7:0] t_r6_c24_7;
  wire [7:0] t_r6_c24_8;
  wire [7:0] t_r6_c24_9;
  wire [7:0] t_r6_c24_10;
  wire [7:0] t_r6_c24_11;
  wire [7:0] t_r6_c24_12;
  wire [7:0] t_r6_c25_0;
  wire [7:0] t_r6_c25_1;
  wire [7:0] t_r6_c25_2;
  wire [7:0] t_r6_c25_3;
  wire [7:0] t_r6_c25_4;
  wire [7:0] t_r6_c25_5;
  wire [7:0] t_r6_c25_6;
  wire [7:0] t_r6_c25_7;
  wire [7:0] t_r6_c25_8;
  wire [7:0] t_r6_c25_9;
  wire [7:0] t_r6_c25_10;
  wire [7:0] t_r6_c25_11;
  wire [7:0] t_r6_c25_12;
  wire [7:0] t_r6_c26_0;
  wire [7:0] t_r6_c26_1;
  wire [7:0] t_r6_c26_2;
  wire [7:0] t_r6_c26_3;
  wire [7:0] t_r6_c26_4;
  wire [7:0] t_r6_c26_5;
  wire [7:0] t_r6_c26_6;
  wire [7:0] t_r6_c26_7;
  wire [7:0] t_r6_c26_8;
  wire [7:0] t_r6_c26_9;
  wire [7:0] t_r6_c26_10;
  wire [7:0] t_r6_c26_11;
  wire [7:0] t_r6_c26_12;
  wire [7:0] t_r6_c27_0;
  wire [7:0] t_r6_c27_1;
  wire [7:0] t_r6_c27_2;
  wire [7:0] t_r6_c27_3;
  wire [7:0] t_r6_c27_4;
  wire [7:0] t_r6_c27_5;
  wire [7:0] t_r6_c27_6;
  wire [7:0] t_r6_c27_7;
  wire [7:0] t_r6_c27_8;
  wire [7:0] t_r6_c27_9;
  wire [7:0] t_r6_c27_10;
  wire [7:0] t_r6_c27_11;
  wire [7:0] t_r6_c27_12;
  wire [7:0] t_r6_c28_0;
  wire [7:0] t_r6_c28_1;
  wire [7:0] t_r6_c28_2;
  wire [7:0] t_r6_c28_3;
  wire [7:0] t_r6_c28_4;
  wire [7:0] t_r6_c28_5;
  wire [7:0] t_r6_c28_6;
  wire [7:0] t_r6_c28_7;
  wire [7:0] t_r6_c28_8;
  wire [7:0] t_r6_c28_9;
  wire [7:0] t_r6_c28_10;
  wire [7:0] t_r6_c28_11;
  wire [7:0] t_r6_c28_12;
  wire [7:0] t_r6_c29_0;
  wire [7:0] t_r6_c29_1;
  wire [7:0] t_r6_c29_2;
  wire [7:0] t_r6_c29_3;
  wire [7:0] t_r6_c29_4;
  wire [7:0] t_r6_c29_5;
  wire [7:0] t_r6_c29_6;
  wire [7:0] t_r6_c29_7;
  wire [7:0] t_r6_c29_8;
  wire [7:0] t_r6_c29_9;
  wire [7:0] t_r6_c29_10;
  wire [7:0] t_r6_c29_11;
  wire [7:0] t_r6_c29_12;
  wire [7:0] t_r6_c30_0;
  wire [7:0] t_r6_c30_1;
  wire [7:0] t_r6_c30_2;
  wire [7:0] t_r6_c30_3;
  wire [7:0] t_r6_c30_4;
  wire [7:0] t_r6_c30_5;
  wire [7:0] t_r6_c30_6;
  wire [7:0] t_r6_c30_7;
  wire [7:0] t_r6_c30_8;
  wire [7:0] t_r6_c30_9;
  wire [7:0] t_r6_c30_10;
  wire [7:0] t_r6_c30_11;
  wire [7:0] t_r6_c30_12;
  wire [7:0] t_r6_c31_0;
  wire [7:0] t_r6_c31_1;
  wire [7:0] t_r6_c31_2;
  wire [7:0] t_r6_c31_3;
  wire [7:0] t_r6_c31_4;
  wire [7:0] t_r6_c31_5;
  wire [7:0] t_r6_c31_6;
  wire [7:0] t_r6_c31_7;
  wire [7:0] t_r6_c31_8;
  wire [7:0] t_r6_c31_9;
  wire [7:0] t_r6_c31_10;
  wire [7:0] t_r6_c31_11;
  wire [7:0] t_r6_c31_12;
  wire [7:0] t_r6_c32_0;
  wire [7:0] t_r6_c32_1;
  wire [7:0] t_r6_c32_2;
  wire [7:0] t_r6_c32_3;
  wire [7:0] t_r6_c32_4;
  wire [7:0] t_r6_c32_5;
  wire [7:0] t_r6_c32_6;
  wire [7:0] t_r6_c32_7;
  wire [7:0] t_r6_c32_8;
  wire [7:0] t_r6_c32_9;
  wire [7:0] t_r6_c32_10;
  wire [7:0] t_r6_c32_11;
  wire [7:0] t_r6_c32_12;
  wire [7:0] t_r6_c33_0;
  wire [7:0] t_r6_c33_1;
  wire [7:0] t_r6_c33_2;
  wire [7:0] t_r6_c33_3;
  wire [7:0] t_r6_c33_4;
  wire [7:0] t_r6_c33_5;
  wire [7:0] t_r6_c33_6;
  wire [7:0] t_r6_c33_7;
  wire [7:0] t_r6_c33_8;
  wire [7:0] t_r6_c33_9;
  wire [7:0] t_r6_c33_10;
  wire [7:0] t_r6_c33_11;
  wire [7:0] t_r6_c33_12;
  wire [7:0] t_r6_c34_0;
  wire [7:0] t_r6_c34_1;
  wire [7:0] t_r6_c34_2;
  wire [7:0] t_r6_c34_3;
  wire [7:0] t_r6_c34_4;
  wire [7:0] t_r6_c34_5;
  wire [7:0] t_r6_c34_6;
  wire [7:0] t_r6_c34_7;
  wire [7:0] t_r6_c34_8;
  wire [7:0] t_r6_c34_9;
  wire [7:0] t_r6_c34_10;
  wire [7:0] t_r6_c34_11;
  wire [7:0] t_r6_c34_12;
  wire [7:0] t_r6_c35_0;
  wire [7:0] t_r6_c35_1;
  wire [7:0] t_r6_c35_2;
  wire [7:0] t_r6_c35_3;
  wire [7:0] t_r6_c35_4;
  wire [7:0] t_r6_c35_5;
  wire [7:0] t_r6_c35_6;
  wire [7:0] t_r6_c35_7;
  wire [7:0] t_r6_c35_8;
  wire [7:0] t_r6_c35_9;
  wire [7:0] t_r6_c35_10;
  wire [7:0] t_r6_c35_11;
  wire [7:0] t_r6_c35_12;
  wire [7:0] t_r6_c36_0;
  wire [7:0] t_r6_c36_1;
  wire [7:0] t_r6_c36_2;
  wire [7:0] t_r6_c36_3;
  wire [7:0] t_r6_c36_4;
  wire [7:0] t_r6_c36_5;
  wire [7:0] t_r6_c36_6;
  wire [7:0] t_r6_c36_7;
  wire [7:0] t_r6_c36_8;
  wire [7:0] t_r6_c36_9;
  wire [7:0] t_r6_c36_10;
  wire [7:0] t_r6_c36_11;
  wire [7:0] t_r6_c36_12;
  wire [7:0] t_r6_c37_0;
  wire [7:0] t_r6_c37_1;
  wire [7:0] t_r6_c37_2;
  wire [7:0] t_r6_c37_3;
  wire [7:0] t_r6_c37_4;
  wire [7:0] t_r6_c37_5;
  wire [7:0] t_r6_c37_6;
  wire [7:0] t_r6_c37_7;
  wire [7:0] t_r6_c37_8;
  wire [7:0] t_r6_c37_9;
  wire [7:0] t_r6_c37_10;
  wire [7:0] t_r6_c37_11;
  wire [7:0] t_r6_c37_12;
  wire [7:0] t_r6_c38_0;
  wire [7:0] t_r6_c38_1;
  wire [7:0] t_r6_c38_2;
  wire [7:0] t_r6_c38_3;
  wire [7:0] t_r6_c38_4;
  wire [7:0] t_r6_c38_5;
  wire [7:0] t_r6_c38_6;
  wire [7:0] t_r6_c38_7;
  wire [7:0] t_r6_c38_8;
  wire [7:0] t_r6_c38_9;
  wire [7:0] t_r6_c38_10;
  wire [7:0] t_r6_c38_11;
  wire [7:0] t_r6_c38_12;
  wire [7:0] t_r6_c39_0;
  wire [7:0] t_r6_c39_1;
  wire [7:0] t_r6_c39_2;
  wire [7:0] t_r6_c39_3;
  wire [7:0] t_r6_c39_4;
  wire [7:0] t_r6_c39_5;
  wire [7:0] t_r6_c39_6;
  wire [7:0] t_r6_c39_7;
  wire [7:0] t_r6_c39_8;
  wire [7:0] t_r6_c39_9;
  wire [7:0] t_r6_c39_10;
  wire [7:0] t_r6_c39_11;
  wire [7:0] t_r6_c39_12;
  wire [7:0] t_r6_c40_0;
  wire [7:0] t_r6_c40_1;
  wire [7:0] t_r6_c40_2;
  wire [7:0] t_r6_c40_3;
  wire [7:0] t_r6_c40_4;
  wire [7:0] t_r6_c40_5;
  wire [7:0] t_r6_c40_6;
  wire [7:0] t_r6_c40_7;
  wire [7:0] t_r6_c40_8;
  wire [7:0] t_r6_c40_9;
  wire [7:0] t_r6_c40_10;
  wire [7:0] t_r6_c40_11;
  wire [7:0] t_r6_c40_12;
  wire [7:0] t_r6_c41_0;
  wire [7:0] t_r6_c41_1;
  wire [7:0] t_r6_c41_2;
  wire [7:0] t_r6_c41_3;
  wire [7:0] t_r6_c41_4;
  wire [7:0] t_r6_c41_5;
  wire [7:0] t_r6_c41_6;
  wire [7:0] t_r6_c41_7;
  wire [7:0] t_r6_c41_8;
  wire [7:0] t_r6_c41_9;
  wire [7:0] t_r6_c41_10;
  wire [7:0] t_r6_c41_11;
  wire [7:0] t_r6_c41_12;
  wire [7:0] t_r6_c42_0;
  wire [7:0] t_r6_c42_1;
  wire [7:0] t_r6_c42_2;
  wire [7:0] t_r6_c42_3;
  wire [7:0] t_r6_c42_4;
  wire [7:0] t_r6_c42_5;
  wire [7:0] t_r6_c42_6;
  wire [7:0] t_r6_c42_7;
  wire [7:0] t_r6_c42_8;
  wire [7:0] t_r6_c42_9;
  wire [7:0] t_r6_c42_10;
  wire [7:0] t_r6_c42_11;
  wire [7:0] t_r6_c42_12;
  wire [7:0] t_r6_c43_0;
  wire [7:0] t_r6_c43_1;
  wire [7:0] t_r6_c43_2;
  wire [7:0] t_r6_c43_3;
  wire [7:0] t_r6_c43_4;
  wire [7:0] t_r6_c43_5;
  wire [7:0] t_r6_c43_6;
  wire [7:0] t_r6_c43_7;
  wire [7:0] t_r6_c43_8;
  wire [7:0] t_r6_c43_9;
  wire [7:0] t_r6_c43_10;
  wire [7:0] t_r6_c43_11;
  wire [7:0] t_r6_c43_12;
  wire [7:0] t_r6_c44_0;
  wire [7:0] t_r6_c44_1;
  wire [7:0] t_r6_c44_2;
  wire [7:0] t_r6_c44_3;
  wire [7:0] t_r6_c44_4;
  wire [7:0] t_r6_c44_5;
  wire [7:0] t_r6_c44_6;
  wire [7:0] t_r6_c44_7;
  wire [7:0] t_r6_c44_8;
  wire [7:0] t_r6_c44_9;
  wire [7:0] t_r6_c44_10;
  wire [7:0] t_r6_c44_11;
  wire [7:0] t_r6_c44_12;
  wire [7:0] t_r6_c45_0;
  wire [7:0] t_r6_c45_1;
  wire [7:0] t_r6_c45_2;
  wire [7:0] t_r6_c45_3;
  wire [7:0] t_r6_c45_4;
  wire [7:0] t_r6_c45_5;
  wire [7:0] t_r6_c45_6;
  wire [7:0] t_r6_c45_7;
  wire [7:0] t_r6_c45_8;
  wire [7:0] t_r6_c45_9;
  wire [7:0] t_r6_c45_10;
  wire [7:0] t_r6_c45_11;
  wire [7:0] t_r6_c45_12;
  wire [7:0] t_r6_c46_0;
  wire [7:0] t_r6_c46_1;
  wire [7:0] t_r6_c46_2;
  wire [7:0] t_r6_c46_3;
  wire [7:0] t_r6_c46_4;
  wire [7:0] t_r6_c46_5;
  wire [7:0] t_r6_c46_6;
  wire [7:0] t_r6_c46_7;
  wire [7:0] t_r6_c46_8;
  wire [7:0] t_r6_c46_9;
  wire [7:0] t_r6_c46_10;
  wire [7:0] t_r6_c46_11;
  wire [7:0] t_r6_c46_12;
  wire [7:0] t_r6_c47_0;
  wire [7:0] t_r6_c47_1;
  wire [7:0] t_r6_c47_2;
  wire [7:0] t_r6_c47_3;
  wire [7:0] t_r6_c47_4;
  wire [7:0] t_r6_c47_5;
  wire [7:0] t_r6_c47_6;
  wire [7:0] t_r6_c47_7;
  wire [7:0] t_r6_c47_8;
  wire [7:0] t_r6_c47_9;
  wire [7:0] t_r6_c47_10;
  wire [7:0] t_r6_c47_11;
  wire [7:0] t_r6_c47_12;
  wire [7:0] t_r6_c48_0;
  wire [7:0] t_r6_c48_1;
  wire [7:0] t_r6_c48_2;
  wire [7:0] t_r6_c48_3;
  wire [7:0] t_r6_c48_4;
  wire [7:0] t_r6_c48_5;
  wire [7:0] t_r6_c48_6;
  wire [7:0] t_r6_c48_7;
  wire [7:0] t_r6_c48_8;
  wire [7:0] t_r6_c48_9;
  wire [7:0] t_r6_c48_10;
  wire [7:0] t_r6_c48_11;
  wire [7:0] t_r6_c48_12;
  wire [7:0] t_r6_c49_0;
  wire [7:0] t_r6_c49_1;
  wire [7:0] t_r6_c49_2;
  wire [7:0] t_r6_c49_3;
  wire [7:0] t_r6_c49_4;
  wire [7:0] t_r6_c49_5;
  wire [7:0] t_r6_c49_6;
  wire [7:0] t_r6_c49_7;
  wire [7:0] t_r6_c49_8;
  wire [7:0] t_r6_c49_9;
  wire [7:0] t_r6_c49_10;
  wire [7:0] t_r6_c49_11;
  wire [7:0] t_r6_c49_12;
  wire [7:0] t_r6_c50_0;
  wire [7:0] t_r6_c50_1;
  wire [7:0] t_r6_c50_2;
  wire [7:0] t_r6_c50_3;
  wire [7:0] t_r6_c50_4;
  wire [7:0] t_r6_c50_5;
  wire [7:0] t_r6_c50_6;
  wire [7:0] t_r6_c50_7;
  wire [7:0] t_r6_c50_8;
  wire [7:0] t_r6_c50_9;
  wire [7:0] t_r6_c50_10;
  wire [7:0] t_r6_c50_11;
  wire [7:0] t_r6_c50_12;
  wire [7:0] t_r6_c51_0;
  wire [7:0] t_r6_c51_1;
  wire [7:0] t_r6_c51_2;
  wire [7:0] t_r6_c51_3;
  wire [7:0] t_r6_c51_4;
  wire [7:0] t_r6_c51_5;
  wire [7:0] t_r6_c51_6;
  wire [7:0] t_r6_c51_7;
  wire [7:0] t_r6_c51_8;
  wire [7:0] t_r6_c51_9;
  wire [7:0] t_r6_c51_10;
  wire [7:0] t_r6_c51_11;
  wire [7:0] t_r6_c51_12;
  wire [7:0] t_r6_c52_0;
  wire [7:0] t_r6_c52_1;
  wire [7:0] t_r6_c52_2;
  wire [7:0] t_r6_c52_3;
  wire [7:0] t_r6_c52_4;
  wire [7:0] t_r6_c52_5;
  wire [7:0] t_r6_c52_6;
  wire [7:0] t_r6_c52_7;
  wire [7:0] t_r6_c52_8;
  wire [7:0] t_r6_c52_9;
  wire [7:0] t_r6_c52_10;
  wire [7:0] t_r6_c52_11;
  wire [7:0] t_r6_c52_12;
  wire [7:0] t_r6_c53_0;
  wire [7:0] t_r6_c53_1;
  wire [7:0] t_r6_c53_2;
  wire [7:0] t_r6_c53_3;
  wire [7:0] t_r6_c53_4;
  wire [7:0] t_r6_c53_5;
  wire [7:0] t_r6_c53_6;
  wire [7:0] t_r6_c53_7;
  wire [7:0] t_r6_c53_8;
  wire [7:0] t_r6_c53_9;
  wire [7:0] t_r6_c53_10;
  wire [7:0] t_r6_c53_11;
  wire [7:0] t_r6_c53_12;
  wire [7:0] t_r6_c54_0;
  wire [7:0] t_r6_c54_1;
  wire [7:0] t_r6_c54_2;
  wire [7:0] t_r6_c54_3;
  wire [7:0] t_r6_c54_4;
  wire [7:0] t_r6_c54_5;
  wire [7:0] t_r6_c54_6;
  wire [7:0] t_r6_c54_7;
  wire [7:0] t_r6_c54_8;
  wire [7:0] t_r6_c54_9;
  wire [7:0] t_r6_c54_10;
  wire [7:0] t_r6_c54_11;
  wire [7:0] t_r6_c54_12;
  wire [7:0] t_r6_c55_0;
  wire [7:0] t_r6_c55_1;
  wire [7:0] t_r6_c55_2;
  wire [7:0] t_r6_c55_3;
  wire [7:0] t_r6_c55_4;
  wire [7:0] t_r6_c55_5;
  wire [7:0] t_r6_c55_6;
  wire [7:0] t_r6_c55_7;
  wire [7:0] t_r6_c55_8;
  wire [7:0] t_r6_c55_9;
  wire [7:0] t_r6_c55_10;
  wire [7:0] t_r6_c55_11;
  wire [7:0] t_r6_c55_12;
  wire [7:0] t_r6_c56_0;
  wire [7:0] t_r6_c56_1;
  wire [7:0] t_r6_c56_2;
  wire [7:0] t_r6_c56_3;
  wire [7:0] t_r6_c56_4;
  wire [7:0] t_r6_c56_5;
  wire [7:0] t_r6_c56_6;
  wire [7:0] t_r6_c56_7;
  wire [7:0] t_r6_c56_8;
  wire [7:0] t_r6_c56_9;
  wire [7:0] t_r6_c56_10;
  wire [7:0] t_r6_c56_11;
  wire [7:0] t_r6_c56_12;
  wire [7:0] t_r6_c57_0;
  wire [7:0] t_r6_c57_1;
  wire [7:0] t_r6_c57_2;
  wire [7:0] t_r6_c57_3;
  wire [7:0] t_r6_c57_4;
  wire [7:0] t_r6_c57_5;
  wire [7:0] t_r6_c57_6;
  wire [7:0] t_r6_c57_7;
  wire [7:0] t_r6_c57_8;
  wire [7:0] t_r6_c57_9;
  wire [7:0] t_r6_c57_10;
  wire [7:0] t_r6_c57_11;
  wire [7:0] t_r6_c57_12;
  wire [7:0] t_r6_c58_0;
  wire [7:0] t_r6_c58_1;
  wire [7:0] t_r6_c58_2;
  wire [7:0] t_r6_c58_3;
  wire [7:0] t_r6_c58_4;
  wire [7:0] t_r6_c58_5;
  wire [7:0] t_r6_c58_6;
  wire [7:0] t_r6_c58_7;
  wire [7:0] t_r6_c58_8;
  wire [7:0] t_r6_c58_9;
  wire [7:0] t_r6_c58_10;
  wire [7:0] t_r6_c58_11;
  wire [7:0] t_r6_c58_12;
  wire [7:0] t_r6_c59_0;
  wire [7:0] t_r6_c59_1;
  wire [7:0] t_r6_c59_2;
  wire [7:0] t_r6_c59_3;
  wire [7:0] t_r6_c59_4;
  wire [7:0] t_r6_c59_5;
  wire [7:0] t_r6_c59_6;
  wire [7:0] t_r6_c59_7;
  wire [7:0] t_r6_c59_8;
  wire [7:0] t_r6_c59_9;
  wire [7:0] t_r6_c59_10;
  wire [7:0] t_r6_c59_11;
  wire [7:0] t_r6_c59_12;
  wire [7:0] t_r6_c60_0;
  wire [7:0] t_r6_c60_1;
  wire [7:0] t_r6_c60_2;
  wire [7:0] t_r6_c60_3;
  wire [7:0] t_r6_c60_4;
  wire [7:0] t_r6_c60_5;
  wire [7:0] t_r6_c60_6;
  wire [7:0] t_r6_c60_7;
  wire [7:0] t_r6_c60_8;
  wire [7:0] t_r6_c60_9;
  wire [7:0] t_r6_c60_10;
  wire [7:0] t_r6_c60_11;
  wire [7:0] t_r6_c60_12;
  wire [7:0] t_r6_c61_0;
  wire [7:0] t_r6_c61_1;
  wire [7:0] t_r6_c61_2;
  wire [7:0] t_r6_c61_3;
  wire [7:0] t_r6_c61_4;
  wire [7:0] t_r6_c61_5;
  wire [7:0] t_r6_c61_6;
  wire [7:0] t_r6_c61_7;
  wire [7:0] t_r6_c61_8;
  wire [7:0] t_r6_c61_9;
  wire [7:0] t_r6_c61_10;
  wire [7:0] t_r6_c61_11;
  wire [7:0] t_r6_c61_12;
  wire [7:0] t_r6_c62_0;
  wire [7:0] t_r6_c62_1;
  wire [7:0] t_r6_c62_2;
  wire [7:0] t_r6_c62_3;
  wire [7:0] t_r6_c62_4;
  wire [7:0] t_r6_c62_5;
  wire [7:0] t_r6_c62_6;
  wire [7:0] t_r6_c62_7;
  wire [7:0] t_r6_c62_8;
  wire [7:0] t_r6_c62_9;
  wire [7:0] t_r6_c62_10;
  wire [7:0] t_r6_c62_11;
  wire [7:0] t_r6_c62_12;
  wire [7:0] t_r6_c63_0;
  wire [7:0] t_r6_c63_1;
  wire [7:0] t_r6_c63_2;
  wire [7:0] t_r6_c63_3;
  wire [7:0] t_r6_c63_4;
  wire [7:0] t_r6_c63_5;
  wire [7:0] t_r6_c63_6;
  wire [7:0] t_r6_c63_7;
  wire [7:0] t_r6_c63_8;
  wire [7:0] t_r6_c63_9;
  wire [7:0] t_r6_c63_10;
  wire [7:0] t_r6_c63_11;
  wire [7:0] t_r6_c63_12;
  wire [7:0] t_r6_c64_0;
  wire [7:0] t_r6_c64_1;
  wire [7:0] t_r6_c64_2;
  wire [7:0] t_r6_c64_3;
  wire [7:0] t_r6_c64_4;
  wire [7:0] t_r6_c64_5;
  wire [7:0] t_r6_c64_6;
  wire [7:0] t_r6_c64_7;
  wire [7:0] t_r6_c64_8;
  wire [7:0] t_r6_c64_9;
  wire [7:0] t_r6_c64_10;
  wire [7:0] t_r6_c64_11;
  wire [7:0] t_r6_c64_12;
  wire [7:0] t_r6_c65_0;
  wire [7:0] t_r6_c65_1;
  wire [7:0] t_r6_c65_2;
  wire [7:0] t_r6_c65_3;
  wire [7:0] t_r6_c65_4;
  wire [7:0] t_r6_c65_5;
  wire [7:0] t_r6_c65_6;
  wire [7:0] t_r6_c65_7;
  wire [7:0] t_r6_c65_8;
  wire [7:0] t_r6_c65_9;
  wire [7:0] t_r6_c65_10;
  wire [7:0] t_r6_c65_11;
  wire [7:0] t_r6_c65_12;
  wire [7:0] t_r7_c0_0;
  wire [7:0] t_r7_c0_1;
  wire [7:0] t_r7_c0_2;
  wire [7:0] t_r7_c0_3;
  wire [7:0] t_r7_c0_4;
  wire [7:0] t_r7_c0_5;
  wire [7:0] t_r7_c0_6;
  wire [7:0] t_r7_c0_7;
  wire [7:0] t_r7_c0_8;
  wire [7:0] t_r7_c0_9;
  wire [7:0] t_r7_c0_10;
  wire [7:0] t_r7_c0_11;
  wire [7:0] t_r7_c0_12;
  wire [7:0] t_r7_c1_0;
  wire [7:0] t_r7_c1_1;
  wire [7:0] t_r7_c1_2;
  wire [7:0] t_r7_c1_3;
  wire [7:0] t_r7_c1_4;
  wire [7:0] t_r7_c1_5;
  wire [7:0] t_r7_c1_6;
  wire [7:0] t_r7_c1_7;
  wire [7:0] t_r7_c1_8;
  wire [7:0] t_r7_c1_9;
  wire [7:0] t_r7_c1_10;
  wire [7:0] t_r7_c1_11;
  wire [7:0] t_r7_c1_12;
  wire [7:0] t_r7_c2_0;
  wire [7:0] t_r7_c2_1;
  wire [7:0] t_r7_c2_2;
  wire [7:0] t_r7_c2_3;
  wire [7:0] t_r7_c2_4;
  wire [7:0] t_r7_c2_5;
  wire [7:0] t_r7_c2_6;
  wire [7:0] t_r7_c2_7;
  wire [7:0] t_r7_c2_8;
  wire [7:0] t_r7_c2_9;
  wire [7:0] t_r7_c2_10;
  wire [7:0] t_r7_c2_11;
  wire [7:0] t_r7_c2_12;
  wire [7:0] t_r7_c3_0;
  wire [7:0] t_r7_c3_1;
  wire [7:0] t_r7_c3_2;
  wire [7:0] t_r7_c3_3;
  wire [7:0] t_r7_c3_4;
  wire [7:0] t_r7_c3_5;
  wire [7:0] t_r7_c3_6;
  wire [7:0] t_r7_c3_7;
  wire [7:0] t_r7_c3_8;
  wire [7:0] t_r7_c3_9;
  wire [7:0] t_r7_c3_10;
  wire [7:0] t_r7_c3_11;
  wire [7:0] t_r7_c3_12;
  wire [7:0] t_r7_c4_0;
  wire [7:0] t_r7_c4_1;
  wire [7:0] t_r7_c4_2;
  wire [7:0] t_r7_c4_3;
  wire [7:0] t_r7_c4_4;
  wire [7:0] t_r7_c4_5;
  wire [7:0] t_r7_c4_6;
  wire [7:0] t_r7_c4_7;
  wire [7:0] t_r7_c4_8;
  wire [7:0] t_r7_c4_9;
  wire [7:0] t_r7_c4_10;
  wire [7:0] t_r7_c4_11;
  wire [7:0] t_r7_c4_12;
  wire [7:0] t_r7_c5_0;
  wire [7:0] t_r7_c5_1;
  wire [7:0] t_r7_c5_2;
  wire [7:0] t_r7_c5_3;
  wire [7:0] t_r7_c5_4;
  wire [7:0] t_r7_c5_5;
  wire [7:0] t_r7_c5_6;
  wire [7:0] t_r7_c5_7;
  wire [7:0] t_r7_c5_8;
  wire [7:0] t_r7_c5_9;
  wire [7:0] t_r7_c5_10;
  wire [7:0] t_r7_c5_11;
  wire [7:0] t_r7_c5_12;
  wire [7:0] t_r7_c6_0;
  wire [7:0] t_r7_c6_1;
  wire [7:0] t_r7_c6_2;
  wire [7:0] t_r7_c6_3;
  wire [7:0] t_r7_c6_4;
  wire [7:0] t_r7_c6_5;
  wire [7:0] t_r7_c6_6;
  wire [7:0] t_r7_c6_7;
  wire [7:0] t_r7_c6_8;
  wire [7:0] t_r7_c6_9;
  wire [7:0] t_r7_c6_10;
  wire [7:0] t_r7_c6_11;
  wire [7:0] t_r7_c6_12;
  wire [7:0] t_r7_c7_0;
  wire [7:0] t_r7_c7_1;
  wire [7:0] t_r7_c7_2;
  wire [7:0] t_r7_c7_3;
  wire [7:0] t_r7_c7_4;
  wire [7:0] t_r7_c7_5;
  wire [7:0] t_r7_c7_6;
  wire [7:0] t_r7_c7_7;
  wire [7:0] t_r7_c7_8;
  wire [7:0] t_r7_c7_9;
  wire [7:0] t_r7_c7_10;
  wire [7:0] t_r7_c7_11;
  wire [7:0] t_r7_c7_12;
  wire [7:0] t_r7_c8_0;
  wire [7:0] t_r7_c8_1;
  wire [7:0] t_r7_c8_2;
  wire [7:0] t_r7_c8_3;
  wire [7:0] t_r7_c8_4;
  wire [7:0] t_r7_c8_5;
  wire [7:0] t_r7_c8_6;
  wire [7:0] t_r7_c8_7;
  wire [7:0] t_r7_c8_8;
  wire [7:0] t_r7_c8_9;
  wire [7:0] t_r7_c8_10;
  wire [7:0] t_r7_c8_11;
  wire [7:0] t_r7_c8_12;
  wire [7:0] t_r7_c9_0;
  wire [7:0] t_r7_c9_1;
  wire [7:0] t_r7_c9_2;
  wire [7:0] t_r7_c9_3;
  wire [7:0] t_r7_c9_4;
  wire [7:0] t_r7_c9_5;
  wire [7:0] t_r7_c9_6;
  wire [7:0] t_r7_c9_7;
  wire [7:0] t_r7_c9_8;
  wire [7:0] t_r7_c9_9;
  wire [7:0] t_r7_c9_10;
  wire [7:0] t_r7_c9_11;
  wire [7:0] t_r7_c9_12;
  wire [7:0] t_r7_c10_0;
  wire [7:0] t_r7_c10_1;
  wire [7:0] t_r7_c10_2;
  wire [7:0] t_r7_c10_3;
  wire [7:0] t_r7_c10_4;
  wire [7:0] t_r7_c10_5;
  wire [7:0] t_r7_c10_6;
  wire [7:0] t_r7_c10_7;
  wire [7:0] t_r7_c10_8;
  wire [7:0] t_r7_c10_9;
  wire [7:0] t_r7_c10_10;
  wire [7:0] t_r7_c10_11;
  wire [7:0] t_r7_c10_12;
  wire [7:0] t_r7_c11_0;
  wire [7:0] t_r7_c11_1;
  wire [7:0] t_r7_c11_2;
  wire [7:0] t_r7_c11_3;
  wire [7:0] t_r7_c11_4;
  wire [7:0] t_r7_c11_5;
  wire [7:0] t_r7_c11_6;
  wire [7:0] t_r7_c11_7;
  wire [7:0] t_r7_c11_8;
  wire [7:0] t_r7_c11_9;
  wire [7:0] t_r7_c11_10;
  wire [7:0] t_r7_c11_11;
  wire [7:0] t_r7_c11_12;
  wire [7:0] t_r7_c12_0;
  wire [7:0] t_r7_c12_1;
  wire [7:0] t_r7_c12_2;
  wire [7:0] t_r7_c12_3;
  wire [7:0] t_r7_c12_4;
  wire [7:0] t_r7_c12_5;
  wire [7:0] t_r7_c12_6;
  wire [7:0] t_r7_c12_7;
  wire [7:0] t_r7_c12_8;
  wire [7:0] t_r7_c12_9;
  wire [7:0] t_r7_c12_10;
  wire [7:0] t_r7_c12_11;
  wire [7:0] t_r7_c12_12;
  wire [7:0] t_r7_c13_0;
  wire [7:0] t_r7_c13_1;
  wire [7:0] t_r7_c13_2;
  wire [7:0] t_r7_c13_3;
  wire [7:0] t_r7_c13_4;
  wire [7:0] t_r7_c13_5;
  wire [7:0] t_r7_c13_6;
  wire [7:0] t_r7_c13_7;
  wire [7:0] t_r7_c13_8;
  wire [7:0] t_r7_c13_9;
  wire [7:0] t_r7_c13_10;
  wire [7:0] t_r7_c13_11;
  wire [7:0] t_r7_c13_12;
  wire [7:0] t_r7_c14_0;
  wire [7:0] t_r7_c14_1;
  wire [7:0] t_r7_c14_2;
  wire [7:0] t_r7_c14_3;
  wire [7:0] t_r7_c14_4;
  wire [7:0] t_r7_c14_5;
  wire [7:0] t_r7_c14_6;
  wire [7:0] t_r7_c14_7;
  wire [7:0] t_r7_c14_8;
  wire [7:0] t_r7_c14_9;
  wire [7:0] t_r7_c14_10;
  wire [7:0] t_r7_c14_11;
  wire [7:0] t_r7_c14_12;
  wire [7:0] t_r7_c15_0;
  wire [7:0] t_r7_c15_1;
  wire [7:0] t_r7_c15_2;
  wire [7:0] t_r7_c15_3;
  wire [7:0] t_r7_c15_4;
  wire [7:0] t_r7_c15_5;
  wire [7:0] t_r7_c15_6;
  wire [7:0] t_r7_c15_7;
  wire [7:0] t_r7_c15_8;
  wire [7:0] t_r7_c15_9;
  wire [7:0] t_r7_c15_10;
  wire [7:0] t_r7_c15_11;
  wire [7:0] t_r7_c15_12;
  wire [7:0] t_r7_c16_0;
  wire [7:0] t_r7_c16_1;
  wire [7:0] t_r7_c16_2;
  wire [7:0] t_r7_c16_3;
  wire [7:0] t_r7_c16_4;
  wire [7:0] t_r7_c16_5;
  wire [7:0] t_r7_c16_6;
  wire [7:0] t_r7_c16_7;
  wire [7:0] t_r7_c16_8;
  wire [7:0] t_r7_c16_9;
  wire [7:0] t_r7_c16_10;
  wire [7:0] t_r7_c16_11;
  wire [7:0] t_r7_c16_12;
  wire [7:0] t_r7_c17_0;
  wire [7:0] t_r7_c17_1;
  wire [7:0] t_r7_c17_2;
  wire [7:0] t_r7_c17_3;
  wire [7:0] t_r7_c17_4;
  wire [7:0] t_r7_c17_5;
  wire [7:0] t_r7_c17_6;
  wire [7:0] t_r7_c17_7;
  wire [7:0] t_r7_c17_8;
  wire [7:0] t_r7_c17_9;
  wire [7:0] t_r7_c17_10;
  wire [7:0] t_r7_c17_11;
  wire [7:0] t_r7_c17_12;
  wire [7:0] t_r7_c18_0;
  wire [7:0] t_r7_c18_1;
  wire [7:0] t_r7_c18_2;
  wire [7:0] t_r7_c18_3;
  wire [7:0] t_r7_c18_4;
  wire [7:0] t_r7_c18_5;
  wire [7:0] t_r7_c18_6;
  wire [7:0] t_r7_c18_7;
  wire [7:0] t_r7_c18_8;
  wire [7:0] t_r7_c18_9;
  wire [7:0] t_r7_c18_10;
  wire [7:0] t_r7_c18_11;
  wire [7:0] t_r7_c18_12;
  wire [7:0] t_r7_c19_0;
  wire [7:0] t_r7_c19_1;
  wire [7:0] t_r7_c19_2;
  wire [7:0] t_r7_c19_3;
  wire [7:0] t_r7_c19_4;
  wire [7:0] t_r7_c19_5;
  wire [7:0] t_r7_c19_6;
  wire [7:0] t_r7_c19_7;
  wire [7:0] t_r7_c19_8;
  wire [7:0] t_r7_c19_9;
  wire [7:0] t_r7_c19_10;
  wire [7:0] t_r7_c19_11;
  wire [7:0] t_r7_c19_12;
  wire [7:0] t_r7_c20_0;
  wire [7:0] t_r7_c20_1;
  wire [7:0] t_r7_c20_2;
  wire [7:0] t_r7_c20_3;
  wire [7:0] t_r7_c20_4;
  wire [7:0] t_r7_c20_5;
  wire [7:0] t_r7_c20_6;
  wire [7:0] t_r7_c20_7;
  wire [7:0] t_r7_c20_8;
  wire [7:0] t_r7_c20_9;
  wire [7:0] t_r7_c20_10;
  wire [7:0] t_r7_c20_11;
  wire [7:0] t_r7_c20_12;
  wire [7:0] t_r7_c21_0;
  wire [7:0] t_r7_c21_1;
  wire [7:0] t_r7_c21_2;
  wire [7:0] t_r7_c21_3;
  wire [7:0] t_r7_c21_4;
  wire [7:0] t_r7_c21_5;
  wire [7:0] t_r7_c21_6;
  wire [7:0] t_r7_c21_7;
  wire [7:0] t_r7_c21_8;
  wire [7:0] t_r7_c21_9;
  wire [7:0] t_r7_c21_10;
  wire [7:0] t_r7_c21_11;
  wire [7:0] t_r7_c21_12;
  wire [7:0] t_r7_c22_0;
  wire [7:0] t_r7_c22_1;
  wire [7:0] t_r7_c22_2;
  wire [7:0] t_r7_c22_3;
  wire [7:0] t_r7_c22_4;
  wire [7:0] t_r7_c22_5;
  wire [7:0] t_r7_c22_6;
  wire [7:0] t_r7_c22_7;
  wire [7:0] t_r7_c22_8;
  wire [7:0] t_r7_c22_9;
  wire [7:0] t_r7_c22_10;
  wire [7:0] t_r7_c22_11;
  wire [7:0] t_r7_c22_12;
  wire [7:0] t_r7_c23_0;
  wire [7:0] t_r7_c23_1;
  wire [7:0] t_r7_c23_2;
  wire [7:0] t_r7_c23_3;
  wire [7:0] t_r7_c23_4;
  wire [7:0] t_r7_c23_5;
  wire [7:0] t_r7_c23_6;
  wire [7:0] t_r7_c23_7;
  wire [7:0] t_r7_c23_8;
  wire [7:0] t_r7_c23_9;
  wire [7:0] t_r7_c23_10;
  wire [7:0] t_r7_c23_11;
  wire [7:0] t_r7_c23_12;
  wire [7:0] t_r7_c24_0;
  wire [7:0] t_r7_c24_1;
  wire [7:0] t_r7_c24_2;
  wire [7:0] t_r7_c24_3;
  wire [7:0] t_r7_c24_4;
  wire [7:0] t_r7_c24_5;
  wire [7:0] t_r7_c24_6;
  wire [7:0] t_r7_c24_7;
  wire [7:0] t_r7_c24_8;
  wire [7:0] t_r7_c24_9;
  wire [7:0] t_r7_c24_10;
  wire [7:0] t_r7_c24_11;
  wire [7:0] t_r7_c24_12;
  wire [7:0] t_r7_c25_0;
  wire [7:0] t_r7_c25_1;
  wire [7:0] t_r7_c25_2;
  wire [7:0] t_r7_c25_3;
  wire [7:0] t_r7_c25_4;
  wire [7:0] t_r7_c25_5;
  wire [7:0] t_r7_c25_6;
  wire [7:0] t_r7_c25_7;
  wire [7:0] t_r7_c25_8;
  wire [7:0] t_r7_c25_9;
  wire [7:0] t_r7_c25_10;
  wire [7:0] t_r7_c25_11;
  wire [7:0] t_r7_c25_12;
  wire [7:0] t_r7_c26_0;
  wire [7:0] t_r7_c26_1;
  wire [7:0] t_r7_c26_2;
  wire [7:0] t_r7_c26_3;
  wire [7:0] t_r7_c26_4;
  wire [7:0] t_r7_c26_5;
  wire [7:0] t_r7_c26_6;
  wire [7:0] t_r7_c26_7;
  wire [7:0] t_r7_c26_8;
  wire [7:0] t_r7_c26_9;
  wire [7:0] t_r7_c26_10;
  wire [7:0] t_r7_c26_11;
  wire [7:0] t_r7_c26_12;
  wire [7:0] t_r7_c27_0;
  wire [7:0] t_r7_c27_1;
  wire [7:0] t_r7_c27_2;
  wire [7:0] t_r7_c27_3;
  wire [7:0] t_r7_c27_4;
  wire [7:0] t_r7_c27_5;
  wire [7:0] t_r7_c27_6;
  wire [7:0] t_r7_c27_7;
  wire [7:0] t_r7_c27_8;
  wire [7:0] t_r7_c27_9;
  wire [7:0] t_r7_c27_10;
  wire [7:0] t_r7_c27_11;
  wire [7:0] t_r7_c27_12;
  wire [7:0] t_r7_c28_0;
  wire [7:0] t_r7_c28_1;
  wire [7:0] t_r7_c28_2;
  wire [7:0] t_r7_c28_3;
  wire [7:0] t_r7_c28_4;
  wire [7:0] t_r7_c28_5;
  wire [7:0] t_r7_c28_6;
  wire [7:0] t_r7_c28_7;
  wire [7:0] t_r7_c28_8;
  wire [7:0] t_r7_c28_9;
  wire [7:0] t_r7_c28_10;
  wire [7:0] t_r7_c28_11;
  wire [7:0] t_r7_c28_12;
  wire [7:0] t_r7_c29_0;
  wire [7:0] t_r7_c29_1;
  wire [7:0] t_r7_c29_2;
  wire [7:0] t_r7_c29_3;
  wire [7:0] t_r7_c29_4;
  wire [7:0] t_r7_c29_5;
  wire [7:0] t_r7_c29_6;
  wire [7:0] t_r7_c29_7;
  wire [7:0] t_r7_c29_8;
  wire [7:0] t_r7_c29_9;
  wire [7:0] t_r7_c29_10;
  wire [7:0] t_r7_c29_11;
  wire [7:0] t_r7_c29_12;
  wire [7:0] t_r7_c30_0;
  wire [7:0] t_r7_c30_1;
  wire [7:0] t_r7_c30_2;
  wire [7:0] t_r7_c30_3;
  wire [7:0] t_r7_c30_4;
  wire [7:0] t_r7_c30_5;
  wire [7:0] t_r7_c30_6;
  wire [7:0] t_r7_c30_7;
  wire [7:0] t_r7_c30_8;
  wire [7:0] t_r7_c30_9;
  wire [7:0] t_r7_c30_10;
  wire [7:0] t_r7_c30_11;
  wire [7:0] t_r7_c30_12;
  wire [7:0] t_r7_c31_0;
  wire [7:0] t_r7_c31_1;
  wire [7:0] t_r7_c31_2;
  wire [7:0] t_r7_c31_3;
  wire [7:0] t_r7_c31_4;
  wire [7:0] t_r7_c31_5;
  wire [7:0] t_r7_c31_6;
  wire [7:0] t_r7_c31_7;
  wire [7:0] t_r7_c31_8;
  wire [7:0] t_r7_c31_9;
  wire [7:0] t_r7_c31_10;
  wire [7:0] t_r7_c31_11;
  wire [7:0] t_r7_c31_12;
  wire [7:0] t_r7_c32_0;
  wire [7:0] t_r7_c32_1;
  wire [7:0] t_r7_c32_2;
  wire [7:0] t_r7_c32_3;
  wire [7:0] t_r7_c32_4;
  wire [7:0] t_r7_c32_5;
  wire [7:0] t_r7_c32_6;
  wire [7:0] t_r7_c32_7;
  wire [7:0] t_r7_c32_8;
  wire [7:0] t_r7_c32_9;
  wire [7:0] t_r7_c32_10;
  wire [7:0] t_r7_c32_11;
  wire [7:0] t_r7_c32_12;
  wire [7:0] t_r7_c33_0;
  wire [7:0] t_r7_c33_1;
  wire [7:0] t_r7_c33_2;
  wire [7:0] t_r7_c33_3;
  wire [7:0] t_r7_c33_4;
  wire [7:0] t_r7_c33_5;
  wire [7:0] t_r7_c33_6;
  wire [7:0] t_r7_c33_7;
  wire [7:0] t_r7_c33_8;
  wire [7:0] t_r7_c33_9;
  wire [7:0] t_r7_c33_10;
  wire [7:0] t_r7_c33_11;
  wire [7:0] t_r7_c33_12;
  wire [7:0] t_r7_c34_0;
  wire [7:0] t_r7_c34_1;
  wire [7:0] t_r7_c34_2;
  wire [7:0] t_r7_c34_3;
  wire [7:0] t_r7_c34_4;
  wire [7:0] t_r7_c34_5;
  wire [7:0] t_r7_c34_6;
  wire [7:0] t_r7_c34_7;
  wire [7:0] t_r7_c34_8;
  wire [7:0] t_r7_c34_9;
  wire [7:0] t_r7_c34_10;
  wire [7:0] t_r7_c34_11;
  wire [7:0] t_r7_c34_12;
  wire [7:0] t_r7_c35_0;
  wire [7:0] t_r7_c35_1;
  wire [7:0] t_r7_c35_2;
  wire [7:0] t_r7_c35_3;
  wire [7:0] t_r7_c35_4;
  wire [7:0] t_r7_c35_5;
  wire [7:0] t_r7_c35_6;
  wire [7:0] t_r7_c35_7;
  wire [7:0] t_r7_c35_8;
  wire [7:0] t_r7_c35_9;
  wire [7:0] t_r7_c35_10;
  wire [7:0] t_r7_c35_11;
  wire [7:0] t_r7_c35_12;
  wire [7:0] t_r7_c36_0;
  wire [7:0] t_r7_c36_1;
  wire [7:0] t_r7_c36_2;
  wire [7:0] t_r7_c36_3;
  wire [7:0] t_r7_c36_4;
  wire [7:0] t_r7_c36_5;
  wire [7:0] t_r7_c36_6;
  wire [7:0] t_r7_c36_7;
  wire [7:0] t_r7_c36_8;
  wire [7:0] t_r7_c36_9;
  wire [7:0] t_r7_c36_10;
  wire [7:0] t_r7_c36_11;
  wire [7:0] t_r7_c36_12;
  wire [7:0] t_r7_c37_0;
  wire [7:0] t_r7_c37_1;
  wire [7:0] t_r7_c37_2;
  wire [7:0] t_r7_c37_3;
  wire [7:0] t_r7_c37_4;
  wire [7:0] t_r7_c37_5;
  wire [7:0] t_r7_c37_6;
  wire [7:0] t_r7_c37_7;
  wire [7:0] t_r7_c37_8;
  wire [7:0] t_r7_c37_9;
  wire [7:0] t_r7_c37_10;
  wire [7:0] t_r7_c37_11;
  wire [7:0] t_r7_c37_12;
  wire [7:0] t_r7_c38_0;
  wire [7:0] t_r7_c38_1;
  wire [7:0] t_r7_c38_2;
  wire [7:0] t_r7_c38_3;
  wire [7:0] t_r7_c38_4;
  wire [7:0] t_r7_c38_5;
  wire [7:0] t_r7_c38_6;
  wire [7:0] t_r7_c38_7;
  wire [7:0] t_r7_c38_8;
  wire [7:0] t_r7_c38_9;
  wire [7:0] t_r7_c38_10;
  wire [7:0] t_r7_c38_11;
  wire [7:0] t_r7_c38_12;
  wire [7:0] t_r7_c39_0;
  wire [7:0] t_r7_c39_1;
  wire [7:0] t_r7_c39_2;
  wire [7:0] t_r7_c39_3;
  wire [7:0] t_r7_c39_4;
  wire [7:0] t_r7_c39_5;
  wire [7:0] t_r7_c39_6;
  wire [7:0] t_r7_c39_7;
  wire [7:0] t_r7_c39_8;
  wire [7:0] t_r7_c39_9;
  wire [7:0] t_r7_c39_10;
  wire [7:0] t_r7_c39_11;
  wire [7:0] t_r7_c39_12;
  wire [7:0] t_r7_c40_0;
  wire [7:0] t_r7_c40_1;
  wire [7:0] t_r7_c40_2;
  wire [7:0] t_r7_c40_3;
  wire [7:0] t_r7_c40_4;
  wire [7:0] t_r7_c40_5;
  wire [7:0] t_r7_c40_6;
  wire [7:0] t_r7_c40_7;
  wire [7:0] t_r7_c40_8;
  wire [7:0] t_r7_c40_9;
  wire [7:0] t_r7_c40_10;
  wire [7:0] t_r7_c40_11;
  wire [7:0] t_r7_c40_12;
  wire [7:0] t_r7_c41_0;
  wire [7:0] t_r7_c41_1;
  wire [7:0] t_r7_c41_2;
  wire [7:0] t_r7_c41_3;
  wire [7:0] t_r7_c41_4;
  wire [7:0] t_r7_c41_5;
  wire [7:0] t_r7_c41_6;
  wire [7:0] t_r7_c41_7;
  wire [7:0] t_r7_c41_8;
  wire [7:0] t_r7_c41_9;
  wire [7:0] t_r7_c41_10;
  wire [7:0] t_r7_c41_11;
  wire [7:0] t_r7_c41_12;
  wire [7:0] t_r7_c42_0;
  wire [7:0] t_r7_c42_1;
  wire [7:0] t_r7_c42_2;
  wire [7:0] t_r7_c42_3;
  wire [7:0] t_r7_c42_4;
  wire [7:0] t_r7_c42_5;
  wire [7:0] t_r7_c42_6;
  wire [7:0] t_r7_c42_7;
  wire [7:0] t_r7_c42_8;
  wire [7:0] t_r7_c42_9;
  wire [7:0] t_r7_c42_10;
  wire [7:0] t_r7_c42_11;
  wire [7:0] t_r7_c42_12;
  wire [7:0] t_r7_c43_0;
  wire [7:0] t_r7_c43_1;
  wire [7:0] t_r7_c43_2;
  wire [7:0] t_r7_c43_3;
  wire [7:0] t_r7_c43_4;
  wire [7:0] t_r7_c43_5;
  wire [7:0] t_r7_c43_6;
  wire [7:0] t_r7_c43_7;
  wire [7:0] t_r7_c43_8;
  wire [7:0] t_r7_c43_9;
  wire [7:0] t_r7_c43_10;
  wire [7:0] t_r7_c43_11;
  wire [7:0] t_r7_c43_12;
  wire [7:0] t_r7_c44_0;
  wire [7:0] t_r7_c44_1;
  wire [7:0] t_r7_c44_2;
  wire [7:0] t_r7_c44_3;
  wire [7:0] t_r7_c44_4;
  wire [7:0] t_r7_c44_5;
  wire [7:0] t_r7_c44_6;
  wire [7:0] t_r7_c44_7;
  wire [7:0] t_r7_c44_8;
  wire [7:0] t_r7_c44_9;
  wire [7:0] t_r7_c44_10;
  wire [7:0] t_r7_c44_11;
  wire [7:0] t_r7_c44_12;
  wire [7:0] t_r7_c45_0;
  wire [7:0] t_r7_c45_1;
  wire [7:0] t_r7_c45_2;
  wire [7:0] t_r7_c45_3;
  wire [7:0] t_r7_c45_4;
  wire [7:0] t_r7_c45_5;
  wire [7:0] t_r7_c45_6;
  wire [7:0] t_r7_c45_7;
  wire [7:0] t_r7_c45_8;
  wire [7:0] t_r7_c45_9;
  wire [7:0] t_r7_c45_10;
  wire [7:0] t_r7_c45_11;
  wire [7:0] t_r7_c45_12;
  wire [7:0] t_r7_c46_0;
  wire [7:0] t_r7_c46_1;
  wire [7:0] t_r7_c46_2;
  wire [7:0] t_r7_c46_3;
  wire [7:0] t_r7_c46_4;
  wire [7:0] t_r7_c46_5;
  wire [7:0] t_r7_c46_6;
  wire [7:0] t_r7_c46_7;
  wire [7:0] t_r7_c46_8;
  wire [7:0] t_r7_c46_9;
  wire [7:0] t_r7_c46_10;
  wire [7:0] t_r7_c46_11;
  wire [7:0] t_r7_c46_12;
  wire [7:0] t_r7_c47_0;
  wire [7:0] t_r7_c47_1;
  wire [7:0] t_r7_c47_2;
  wire [7:0] t_r7_c47_3;
  wire [7:0] t_r7_c47_4;
  wire [7:0] t_r7_c47_5;
  wire [7:0] t_r7_c47_6;
  wire [7:0] t_r7_c47_7;
  wire [7:0] t_r7_c47_8;
  wire [7:0] t_r7_c47_9;
  wire [7:0] t_r7_c47_10;
  wire [7:0] t_r7_c47_11;
  wire [7:0] t_r7_c47_12;
  wire [7:0] t_r7_c48_0;
  wire [7:0] t_r7_c48_1;
  wire [7:0] t_r7_c48_2;
  wire [7:0] t_r7_c48_3;
  wire [7:0] t_r7_c48_4;
  wire [7:0] t_r7_c48_5;
  wire [7:0] t_r7_c48_6;
  wire [7:0] t_r7_c48_7;
  wire [7:0] t_r7_c48_8;
  wire [7:0] t_r7_c48_9;
  wire [7:0] t_r7_c48_10;
  wire [7:0] t_r7_c48_11;
  wire [7:0] t_r7_c48_12;
  wire [7:0] t_r7_c49_0;
  wire [7:0] t_r7_c49_1;
  wire [7:0] t_r7_c49_2;
  wire [7:0] t_r7_c49_3;
  wire [7:0] t_r7_c49_4;
  wire [7:0] t_r7_c49_5;
  wire [7:0] t_r7_c49_6;
  wire [7:0] t_r7_c49_7;
  wire [7:0] t_r7_c49_8;
  wire [7:0] t_r7_c49_9;
  wire [7:0] t_r7_c49_10;
  wire [7:0] t_r7_c49_11;
  wire [7:0] t_r7_c49_12;
  wire [7:0] t_r7_c50_0;
  wire [7:0] t_r7_c50_1;
  wire [7:0] t_r7_c50_2;
  wire [7:0] t_r7_c50_3;
  wire [7:0] t_r7_c50_4;
  wire [7:0] t_r7_c50_5;
  wire [7:0] t_r7_c50_6;
  wire [7:0] t_r7_c50_7;
  wire [7:0] t_r7_c50_8;
  wire [7:0] t_r7_c50_9;
  wire [7:0] t_r7_c50_10;
  wire [7:0] t_r7_c50_11;
  wire [7:0] t_r7_c50_12;
  wire [7:0] t_r7_c51_0;
  wire [7:0] t_r7_c51_1;
  wire [7:0] t_r7_c51_2;
  wire [7:0] t_r7_c51_3;
  wire [7:0] t_r7_c51_4;
  wire [7:0] t_r7_c51_5;
  wire [7:0] t_r7_c51_6;
  wire [7:0] t_r7_c51_7;
  wire [7:0] t_r7_c51_8;
  wire [7:0] t_r7_c51_9;
  wire [7:0] t_r7_c51_10;
  wire [7:0] t_r7_c51_11;
  wire [7:0] t_r7_c51_12;
  wire [7:0] t_r7_c52_0;
  wire [7:0] t_r7_c52_1;
  wire [7:0] t_r7_c52_2;
  wire [7:0] t_r7_c52_3;
  wire [7:0] t_r7_c52_4;
  wire [7:0] t_r7_c52_5;
  wire [7:0] t_r7_c52_6;
  wire [7:0] t_r7_c52_7;
  wire [7:0] t_r7_c52_8;
  wire [7:0] t_r7_c52_9;
  wire [7:0] t_r7_c52_10;
  wire [7:0] t_r7_c52_11;
  wire [7:0] t_r7_c52_12;
  wire [7:0] t_r7_c53_0;
  wire [7:0] t_r7_c53_1;
  wire [7:0] t_r7_c53_2;
  wire [7:0] t_r7_c53_3;
  wire [7:0] t_r7_c53_4;
  wire [7:0] t_r7_c53_5;
  wire [7:0] t_r7_c53_6;
  wire [7:0] t_r7_c53_7;
  wire [7:0] t_r7_c53_8;
  wire [7:0] t_r7_c53_9;
  wire [7:0] t_r7_c53_10;
  wire [7:0] t_r7_c53_11;
  wire [7:0] t_r7_c53_12;
  wire [7:0] t_r7_c54_0;
  wire [7:0] t_r7_c54_1;
  wire [7:0] t_r7_c54_2;
  wire [7:0] t_r7_c54_3;
  wire [7:0] t_r7_c54_4;
  wire [7:0] t_r7_c54_5;
  wire [7:0] t_r7_c54_6;
  wire [7:0] t_r7_c54_7;
  wire [7:0] t_r7_c54_8;
  wire [7:0] t_r7_c54_9;
  wire [7:0] t_r7_c54_10;
  wire [7:0] t_r7_c54_11;
  wire [7:0] t_r7_c54_12;
  wire [7:0] t_r7_c55_0;
  wire [7:0] t_r7_c55_1;
  wire [7:0] t_r7_c55_2;
  wire [7:0] t_r7_c55_3;
  wire [7:0] t_r7_c55_4;
  wire [7:0] t_r7_c55_5;
  wire [7:0] t_r7_c55_6;
  wire [7:0] t_r7_c55_7;
  wire [7:0] t_r7_c55_8;
  wire [7:0] t_r7_c55_9;
  wire [7:0] t_r7_c55_10;
  wire [7:0] t_r7_c55_11;
  wire [7:0] t_r7_c55_12;
  wire [7:0] t_r7_c56_0;
  wire [7:0] t_r7_c56_1;
  wire [7:0] t_r7_c56_2;
  wire [7:0] t_r7_c56_3;
  wire [7:0] t_r7_c56_4;
  wire [7:0] t_r7_c56_5;
  wire [7:0] t_r7_c56_6;
  wire [7:0] t_r7_c56_7;
  wire [7:0] t_r7_c56_8;
  wire [7:0] t_r7_c56_9;
  wire [7:0] t_r7_c56_10;
  wire [7:0] t_r7_c56_11;
  wire [7:0] t_r7_c56_12;
  wire [7:0] t_r7_c57_0;
  wire [7:0] t_r7_c57_1;
  wire [7:0] t_r7_c57_2;
  wire [7:0] t_r7_c57_3;
  wire [7:0] t_r7_c57_4;
  wire [7:0] t_r7_c57_5;
  wire [7:0] t_r7_c57_6;
  wire [7:0] t_r7_c57_7;
  wire [7:0] t_r7_c57_8;
  wire [7:0] t_r7_c57_9;
  wire [7:0] t_r7_c57_10;
  wire [7:0] t_r7_c57_11;
  wire [7:0] t_r7_c57_12;
  wire [7:0] t_r7_c58_0;
  wire [7:0] t_r7_c58_1;
  wire [7:0] t_r7_c58_2;
  wire [7:0] t_r7_c58_3;
  wire [7:0] t_r7_c58_4;
  wire [7:0] t_r7_c58_5;
  wire [7:0] t_r7_c58_6;
  wire [7:0] t_r7_c58_7;
  wire [7:0] t_r7_c58_8;
  wire [7:0] t_r7_c58_9;
  wire [7:0] t_r7_c58_10;
  wire [7:0] t_r7_c58_11;
  wire [7:0] t_r7_c58_12;
  wire [7:0] t_r7_c59_0;
  wire [7:0] t_r7_c59_1;
  wire [7:0] t_r7_c59_2;
  wire [7:0] t_r7_c59_3;
  wire [7:0] t_r7_c59_4;
  wire [7:0] t_r7_c59_5;
  wire [7:0] t_r7_c59_6;
  wire [7:0] t_r7_c59_7;
  wire [7:0] t_r7_c59_8;
  wire [7:0] t_r7_c59_9;
  wire [7:0] t_r7_c59_10;
  wire [7:0] t_r7_c59_11;
  wire [7:0] t_r7_c59_12;
  wire [7:0] t_r7_c60_0;
  wire [7:0] t_r7_c60_1;
  wire [7:0] t_r7_c60_2;
  wire [7:0] t_r7_c60_3;
  wire [7:0] t_r7_c60_4;
  wire [7:0] t_r7_c60_5;
  wire [7:0] t_r7_c60_6;
  wire [7:0] t_r7_c60_7;
  wire [7:0] t_r7_c60_8;
  wire [7:0] t_r7_c60_9;
  wire [7:0] t_r7_c60_10;
  wire [7:0] t_r7_c60_11;
  wire [7:0] t_r7_c60_12;
  wire [7:0] t_r7_c61_0;
  wire [7:0] t_r7_c61_1;
  wire [7:0] t_r7_c61_2;
  wire [7:0] t_r7_c61_3;
  wire [7:0] t_r7_c61_4;
  wire [7:0] t_r7_c61_5;
  wire [7:0] t_r7_c61_6;
  wire [7:0] t_r7_c61_7;
  wire [7:0] t_r7_c61_8;
  wire [7:0] t_r7_c61_9;
  wire [7:0] t_r7_c61_10;
  wire [7:0] t_r7_c61_11;
  wire [7:0] t_r7_c61_12;
  wire [7:0] t_r7_c62_0;
  wire [7:0] t_r7_c62_1;
  wire [7:0] t_r7_c62_2;
  wire [7:0] t_r7_c62_3;
  wire [7:0] t_r7_c62_4;
  wire [7:0] t_r7_c62_5;
  wire [7:0] t_r7_c62_6;
  wire [7:0] t_r7_c62_7;
  wire [7:0] t_r7_c62_8;
  wire [7:0] t_r7_c62_9;
  wire [7:0] t_r7_c62_10;
  wire [7:0] t_r7_c62_11;
  wire [7:0] t_r7_c62_12;
  wire [7:0] t_r7_c63_0;
  wire [7:0] t_r7_c63_1;
  wire [7:0] t_r7_c63_2;
  wire [7:0] t_r7_c63_3;
  wire [7:0] t_r7_c63_4;
  wire [7:0] t_r7_c63_5;
  wire [7:0] t_r7_c63_6;
  wire [7:0] t_r7_c63_7;
  wire [7:0] t_r7_c63_8;
  wire [7:0] t_r7_c63_9;
  wire [7:0] t_r7_c63_10;
  wire [7:0] t_r7_c63_11;
  wire [7:0] t_r7_c63_12;
  wire [7:0] t_r7_c64_0;
  wire [7:0] t_r7_c64_1;
  wire [7:0] t_r7_c64_2;
  wire [7:0] t_r7_c64_3;
  wire [7:0] t_r7_c64_4;
  wire [7:0] t_r7_c64_5;
  wire [7:0] t_r7_c64_6;
  wire [7:0] t_r7_c64_7;
  wire [7:0] t_r7_c64_8;
  wire [7:0] t_r7_c64_9;
  wire [7:0] t_r7_c64_10;
  wire [7:0] t_r7_c64_11;
  wire [7:0] t_r7_c64_12;
  wire [7:0] t_r7_c65_0;
  wire [7:0] t_r7_c65_1;
  wire [7:0] t_r7_c65_2;
  wire [7:0] t_r7_c65_3;
  wire [7:0] t_r7_c65_4;
  wire [7:0] t_r7_c65_5;
  wire [7:0] t_r7_c65_6;
  wire [7:0] t_r7_c65_7;
  wire [7:0] t_r7_c65_8;
  wire [7:0] t_r7_c65_9;
  wire [7:0] t_r7_c65_10;
  wire [7:0] t_r7_c65_11;
  wire [7:0] t_r7_c65_12;
  wire [7:0] t_r8_c0_0;
  wire [7:0] t_r8_c0_1;
  wire [7:0] t_r8_c0_2;
  wire [7:0] t_r8_c0_3;
  wire [7:0] t_r8_c0_4;
  wire [7:0] t_r8_c0_5;
  wire [7:0] t_r8_c0_6;
  wire [7:0] t_r8_c0_7;
  wire [7:0] t_r8_c0_8;
  wire [7:0] t_r8_c0_9;
  wire [7:0] t_r8_c0_10;
  wire [7:0] t_r8_c0_11;
  wire [7:0] t_r8_c0_12;
  wire [7:0] t_r8_c1_0;
  wire [7:0] t_r8_c1_1;
  wire [7:0] t_r8_c1_2;
  wire [7:0] t_r8_c1_3;
  wire [7:0] t_r8_c1_4;
  wire [7:0] t_r8_c1_5;
  wire [7:0] t_r8_c1_6;
  wire [7:0] t_r8_c1_7;
  wire [7:0] t_r8_c1_8;
  wire [7:0] t_r8_c1_9;
  wire [7:0] t_r8_c1_10;
  wire [7:0] t_r8_c1_11;
  wire [7:0] t_r8_c1_12;
  wire [7:0] t_r8_c2_0;
  wire [7:0] t_r8_c2_1;
  wire [7:0] t_r8_c2_2;
  wire [7:0] t_r8_c2_3;
  wire [7:0] t_r8_c2_4;
  wire [7:0] t_r8_c2_5;
  wire [7:0] t_r8_c2_6;
  wire [7:0] t_r8_c2_7;
  wire [7:0] t_r8_c2_8;
  wire [7:0] t_r8_c2_9;
  wire [7:0] t_r8_c2_10;
  wire [7:0] t_r8_c2_11;
  wire [7:0] t_r8_c2_12;
  wire [7:0] t_r8_c3_0;
  wire [7:0] t_r8_c3_1;
  wire [7:0] t_r8_c3_2;
  wire [7:0] t_r8_c3_3;
  wire [7:0] t_r8_c3_4;
  wire [7:0] t_r8_c3_5;
  wire [7:0] t_r8_c3_6;
  wire [7:0] t_r8_c3_7;
  wire [7:0] t_r8_c3_8;
  wire [7:0] t_r8_c3_9;
  wire [7:0] t_r8_c3_10;
  wire [7:0] t_r8_c3_11;
  wire [7:0] t_r8_c3_12;
  wire [7:0] t_r8_c4_0;
  wire [7:0] t_r8_c4_1;
  wire [7:0] t_r8_c4_2;
  wire [7:0] t_r8_c4_3;
  wire [7:0] t_r8_c4_4;
  wire [7:0] t_r8_c4_5;
  wire [7:0] t_r8_c4_6;
  wire [7:0] t_r8_c4_7;
  wire [7:0] t_r8_c4_8;
  wire [7:0] t_r8_c4_9;
  wire [7:0] t_r8_c4_10;
  wire [7:0] t_r8_c4_11;
  wire [7:0] t_r8_c4_12;
  wire [7:0] t_r8_c5_0;
  wire [7:0] t_r8_c5_1;
  wire [7:0] t_r8_c5_2;
  wire [7:0] t_r8_c5_3;
  wire [7:0] t_r8_c5_4;
  wire [7:0] t_r8_c5_5;
  wire [7:0] t_r8_c5_6;
  wire [7:0] t_r8_c5_7;
  wire [7:0] t_r8_c5_8;
  wire [7:0] t_r8_c5_9;
  wire [7:0] t_r8_c5_10;
  wire [7:0] t_r8_c5_11;
  wire [7:0] t_r8_c5_12;
  wire [7:0] t_r8_c6_0;
  wire [7:0] t_r8_c6_1;
  wire [7:0] t_r8_c6_2;
  wire [7:0] t_r8_c6_3;
  wire [7:0] t_r8_c6_4;
  wire [7:0] t_r8_c6_5;
  wire [7:0] t_r8_c6_6;
  wire [7:0] t_r8_c6_7;
  wire [7:0] t_r8_c6_8;
  wire [7:0] t_r8_c6_9;
  wire [7:0] t_r8_c6_10;
  wire [7:0] t_r8_c6_11;
  wire [7:0] t_r8_c6_12;
  wire [7:0] t_r8_c7_0;
  wire [7:0] t_r8_c7_1;
  wire [7:0] t_r8_c7_2;
  wire [7:0] t_r8_c7_3;
  wire [7:0] t_r8_c7_4;
  wire [7:0] t_r8_c7_5;
  wire [7:0] t_r8_c7_6;
  wire [7:0] t_r8_c7_7;
  wire [7:0] t_r8_c7_8;
  wire [7:0] t_r8_c7_9;
  wire [7:0] t_r8_c7_10;
  wire [7:0] t_r8_c7_11;
  wire [7:0] t_r8_c7_12;
  wire [7:0] t_r8_c8_0;
  wire [7:0] t_r8_c8_1;
  wire [7:0] t_r8_c8_2;
  wire [7:0] t_r8_c8_3;
  wire [7:0] t_r8_c8_4;
  wire [7:0] t_r8_c8_5;
  wire [7:0] t_r8_c8_6;
  wire [7:0] t_r8_c8_7;
  wire [7:0] t_r8_c8_8;
  wire [7:0] t_r8_c8_9;
  wire [7:0] t_r8_c8_10;
  wire [7:0] t_r8_c8_11;
  wire [7:0] t_r8_c8_12;
  wire [7:0] t_r8_c9_0;
  wire [7:0] t_r8_c9_1;
  wire [7:0] t_r8_c9_2;
  wire [7:0] t_r8_c9_3;
  wire [7:0] t_r8_c9_4;
  wire [7:0] t_r8_c9_5;
  wire [7:0] t_r8_c9_6;
  wire [7:0] t_r8_c9_7;
  wire [7:0] t_r8_c9_8;
  wire [7:0] t_r8_c9_9;
  wire [7:0] t_r8_c9_10;
  wire [7:0] t_r8_c9_11;
  wire [7:0] t_r8_c9_12;
  wire [7:0] t_r8_c10_0;
  wire [7:0] t_r8_c10_1;
  wire [7:0] t_r8_c10_2;
  wire [7:0] t_r8_c10_3;
  wire [7:0] t_r8_c10_4;
  wire [7:0] t_r8_c10_5;
  wire [7:0] t_r8_c10_6;
  wire [7:0] t_r8_c10_7;
  wire [7:0] t_r8_c10_8;
  wire [7:0] t_r8_c10_9;
  wire [7:0] t_r8_c10_10;
  wire [7:0] t_r8_c10_11;
  wire [7:0] t_r8_c10_12;
  wire [7:0] t_r8_c11_0;
  wire [7:0] t_r8_c11_1;
  wire [7:0] t_r8_c11_2;
  wire [7:0] t_r8_c11_3;
  wire [7:0] t_r8_c11_4;
  wire [7:0] t_r8_c11_5;
  wire [7:0] t_r8_c11_6;
  wire [7:0] t_r8_c11_7;
  wire [7:0] t_r8_c11_8;
  wire [7:0] t_r8_c11_9;
  wire [7:0] t_r8_c11_10;
  wire [7:0] t_r8_c11_11;
  wire [7:0] t_r8_c11_12;
  wire [7:0] t_r8_c12_0;
  wire [7:0] t_r8_c12_1;
  wire [7:0] t_r8_c12_2;
  wire [7:0] t_r8_c12_3;
  wire [7:0] t_r8_c12_4;
  wire [7:0] t_r8_c12_5;
  wire [7:0] t_r8_c12_6;
  wire [7:0] t_r8_c12_7;
  wire [7:0] t_r8_c12_8;
  wire [7:0] t_r8_c12_9;
  wire [7:0] t_r8_c12_10;
  wire [7:0] t_r8_c12_11;
  wire [7:0] t_r8_c12_12;
  wire [7:0] t_r8_c13_0;
  wire [7:0] t_r8_c13_1;
  wire [7:0] t_r8_c13_2;
  wire [7:0] t_r8_c13_3;
  wire [7:0] t_r8_c13_4;
  wire [7:0] t_r8_c13_5;
  wire [7:0] t_r8_c13_6;
  wire [7:0] t_r8_c13_7;
  wire [7:0] t_r8_c13_8;
  wire [7:0] t_r8_c13_9;
  wire [7:0] t_r8_c13_10;
  wire [7:0] t_r8_c13_11;
  wire [7:0] t_r8_c13_12;
  wire [7:0] t_r8_c14_0;
  wire [7:0] t_r8_c14_1;
  wire [7:0] t_r8_c14_2;
  wire [7:0] t_r8_c14_3;
  wire [7:0] t_r8_c14_4;
  wire [7:0] t_r8_c14_5;
  wire [7:0] t_r8_c14_6;
  wire [7:0] t_r8_c14_7;
  wire [7:0] t_r8_c14_8;
  wire [7:0] t_r8_c14_9;
  wire [7:0] t_r8_c14_10;
  wire [7:0] t_r8_c14_11;
  wire [7:0] t_r8_c14_12;
  wire [7:0] t_r8_c15_0;
  wire [7:0] t_r8_c15_1;
  wire [7:0] t_r8_c15_2;
  wire [7:0] t_r8_c15_3;
  wire [7:0] t_r8_c15_4;
  wire [7:0] t_r8_c15_5;
  wire [7:0] t_r8_c15_6;
  wire [7:0] t_r8_c15_7;
  wire [7:0] t_r8_c15_8;
  wire [7:0] t_r8_c15_9;
  wire [7:0] t_r8_c15_10;
  wire [7:0] t_r8_c15_11;
  wire [7:0] t_r8_c15_12;
  wire [7:0] t_r8_c16_0;
  wire [7:0] t_r8_c16_1;
  wire [7:0] t_r8_c16_2;
  wire [7:0] t_r8_c16_3;
  wire [7:0] t_r8_c16_4;
  wire [7:0] t_r8_c16_5;
  wire [7:0] t_r8_c16_6;
  wire [7:0] t_r8_c16_7;
  wire [7:0] t_r8_c16_8;
  wire [7:0] t_r8_c16_9;
  wire [7:0] t_r8_c16_10;
  wire [7:0] t_r8_c16_11;
  wire [7:0] t_r8_c16_12;
  wire [7:0] t_r8_c17_0;
  wire [7:0] t_r8_c17_1;
  wire [7:0] t_r8_c17_2;
  wire [7:0] t_r8_c17_3;
  wire [7:0] t_r8_c17_4;
  wire [7:0] t_r8_c17_5;
  wire [7:0] t_r8_c17_6;
  wire [7:0] t_r8_c17_7;
  wire [7:0] t_r8_c17_8;
  wire [7:0] t_r8_c17_9;
  wire [7:0] t_r8_c17_10;
  wire [7:0] t_r8_c17_11;
  wire [7:0] t_r8_c17_12;
  wire [7:0] t_r8_c18_0;
  wire [7:0] t_r8_c18_1;
  wire [7:0] t_r8_c18_2;
  wire [7:0] t_r8_c18_3;
  wire [7:0] t_r8_c18_4;
  wire [7:0] t_r8_c18_5;
  wire [7:0] t_r8_c18_6;
  wire [7:0] t_r8_c18_7;
  wire [7:0] t_r8_c18_8;
  wire [7:0] t_r8_c18_9;
  wire [7:0] t_r8_c18_10;
  wire [7:0] t_r8_c18_11;
  wire [7:0] t_r8_c18_12;
  wire [7:0] t_r8_c19_0;
  wire [7:0] t_r8_c19_1;
  wire [7:0] t_r8_c19_2;
  wire [7:0] t_r8_c19_3;
  wire [7:0] t_r8_c19_4;
  wire [7:0] t_r8_c19_5;
  wire [7:0] t_r8_c19_6;
  wire [7:0] t_r8_c19_7;
  wire [7:0] t_r8_c19_8;
  wire [7:0] t_r8_c19_9;
  wire [7:0] t_r8_c19_10;
  wire [7:0] t_r8_c19_11;
  wire [7:0] t_r8_c19_12;
  wire [7:0] t_r8_c20_0;
  wire [7:0] t_r8_c20_1;
  wire [7:0] t_r8_c20_2;
  wire [7:0] t_r8_c20_3;
  wire [7:0] t_r8_c20_4;
  wire [7:0] t_r8_c20_5;
  wire [7:0] t_r8_c20_6;
  wire [7:0] t_r8_c20_7;
  wire [7:0] t_r8_c20_8;
  wire [7:0] t_r8_c20_9;
  wire [7:0] t_r8_c20_10;
  wire [7:0] t_r8_c20_11;
  wire [7:0] t_r8_c20_12;
  wire [7:0] t_r8_c21_0;
  wire [7:0] t_r8_c21_1;
  wire [7:0] t_r8_c21_2;
  wire [7:0] t_r8_c21_3;
  wire [7:0] t_r8_c21_4;
  wire [7:0] t_r8_c21_5;
  wire [7:0] t_r8_c21_6;
  wire [7:0] t_r8_c21_7;
  wire [7:0] t_r8_c21_8;
  wire [7:0] t_r8_c21_9;
  wire [7:0] t_r8_c21_10;
  wire [7:0] t_r8_c21_11;
  wire [7:0] t_r8_c21_12;
  wire [7:0] t_r8_c22_0;
  wire [7:0] t_r8_c22_1;
  wire [7:0] t_r8_c22_2;
  wire [7:0] t_r8_c22_3;
  wire [7:0] t_r8_c22_4;
  wire [7:0] t_r8_c22_5;
  wire [7:0] t_r8_c22_6;
  wire [7:0] t_r8_c22_7;
  wire [7:0] t_r8_c22_8;
  wire [7:0] t_r8_c22_9;
  wire [7:0] t_r8_c22_10;
  wire [7:0] t_r8_c22_11;
  wire [7:0] t_r8_c22_12;
  wire [7:0] t_r8_c23_0;
  wire [7:0] t_r8_c23_1;
  wire [7:0] t_r8_c23_2;
  wire [7:0] t_r8_c23_3;
  wire [7:0] t_r8_c23_4;
  wire [7:0] t_r8_c23_5;
  wire [7:0] t_r8_c23_6;
  wire [7:0] t_r8_c23_7;
  wire [7:0] t_r8_c23_8;
  wire [7:0] t_r8_c23_9;
  wire [7:0] t_r8_c23_10;
  wire [7:0] t_r8_c23_11;
  wire [7:0] t_r8_c23_12;
  wire [7:0] t_r8_c24_0;
  wire [7:0] t_r8_c24_1;
  wire [7:0] t_r8_c24_2;
  wire [7:0] t_r8_c24_3;
  wire [7:0] t_r8_c24_4;
  wire [7:0] t_r8_c24_5;
  wire [7:0] t_r8_c24_6;
  wire [7:0] t_r8_c24_7;
  wire [7:0] t_r8_c24_8;
  wire [7:0] t_r8_c24_9;
  wire [7:0] t_r8_c24_10;
  wire [7:0] t_r8_c24_11;
  wire [7:0] t_r8_c24_12;
  wire [7:0] t_r8_c25_0;
  wire [7:0] t_r8_c25_1;
  wire [7:0] t_r8_c25_2;
  wire [7:0] t_r8_c25_3;
  wire [7:0] t_r8_c25_4;
  wire [7:0] t_r8_c25_5;
  wire [7:0] t_r8_c25_6;
  wire [7:0] t_r8_c25_7;
  wire [7:0] t_r8_c25_8;
  wire [7:0] t_r8_c25_9;
  wire [7:0] t_r8_c25_10;
  wire [7:0] t_r8_c25_11;
  wire [7:0] t_r8_c25_12;
  wire [7:0] t_r8_c26_0;
  wire [7:0] t_r8_c26_1;
  wire [7:0] t_r8_c26_2;
  wire [7:0] t_r8_c26_3;
  wire [7:0] t_r8_c26_4;
  wire [7:0] t_r8_c26_5;
  wire [7:0] t_r8_c26_6;
  wire [7:0] t_r8_c26_7;
  wire [7:0] t_r8_c26_8;
  wire [7:0] t_r8_c26_9;
  wire [7:0] t_r8_c26_10;
  wire [7:0] t_r8_c26_11;
  wire [7:0] t_r8_c26_12;
  wire [7:0] t_r8_c27_0;
  wire [7:0] t_r8_c27_1;
  wire [7:0] t_r8_c27_2;
  wire [7:0] t_r8_c27_3;
  wire [7:0] t_r8_c27_4;
  wire [7:0] t_r8_c27_5;
  wire [7:0] t_r8_c27_6;
  wire [7:0] t_r8_c27_7;
  wire [7:0] t_r8_c27_8;
  wire [7:0] t_r8_c27_9;
  wire [7:0] t_r8_c27_10;
  wire [7:0] t_r8_c27_11;
  wire [7:0] t_r8_c27_12;
  wire [7:0] t_r8_c28_0;
  wire [7:0] t_r8_c28_1;
  wire [7:0] t_r8_c28_2;
  wire [7:0] t_r8_c28_3;
  wire [7:0] t_r8_c28_4;
  wire [7:0] t_r8_c28_5;
  wire [7:0] t_r8_c28_6;
  wire [7:0] t_r8_c28_7;
  wire [7:0] t_r8_c28_8;
  wire [7:0] t_r8_c28_9;
  wire [7:0] t_r8_c28_10;
  wire [7:0] t_r8_c28_11;
  wire [7:0] t_r8_c28_12;
  wire [7:0] t_r8_c29_0;
  wire [7:0] t_r8_c29_1;
  wire [7:0] t_r8_c29_2;
  wire [7:0] t_r8_c29_3;
  wire [7:0] t_r8_c29_4;
  wire [7:0] t_r8_c29_5;
  wire [7:0] t_r8_c29_6;
  wire [7:0] t_r8_c29_7;
  wire [7:0] t_r8_c29_8;
  wire [7:0] t_r8_c29_9;
  wire [7:0] t_r8_c29_10;
  wire [7:0] t_r8_c29_11;
  wire [7:0] t_r8_c29_12;
  wire [7:0] t_r8_c30_0;
  wire [7:0] t_r8_c30_1;
  wire [7:0] t_r8_c30_2;
  wire [7:0] t_r8_c30_3;
  wire [7:0] t_r8_c30_4;
  wire [7:0] t_r8_c30_5;
  wire [7:0] t_r8_c30_6;
  wire [7:0] t_r8_c30_7;
  wire [7:0] t_r8_c30_8;
  wire [7:0] t_r8_c30_9;
  wire [7:0] t_r8_c30_10;
  wire [7:0] t_r8_c30_11;
  wire [7:0] t_r8_c30_12;
  wire [7:0] t_r8_c31_0;
  wire [7:0] t_r8_c31_1;
  wire [7:0] t_r8_c31_2;
  wire [7:0] t_r8_c31_3;
  wire [7:0] t_r8_c31_4;
  wire [7:0] t_r8_c31_5;
  wire [7:0] t_r8_c31_6;
  wire [7:0] t_r8_c31_7;
  wire [7:0] t_r8_c31_8;
  wire [7:0] t_r8_c31_9;
  wire [7:0] t_r8_c31_10;
  wire [7:0] t_r8_c31_11;
  wire [7:0] t_r8_c31_12;
  wire [7:0] t_r8_c32_0;
  wire [7:0] t_r8_c32_1;
  wire [7:0] t_r8_c32_2;
  wire [7:0] t_r8_c32_3;
  wire [7:0] t_r8_c32_4;
  wire [7:0] t_r8_c32_5;
  wire [7:0] t_r8_c32_6;
  wire [7:0] t_r8_c32_7;
  wire [7:0] t_r8_c32_8;
  wire [7:0] t_r8_c32_9;
  wire [7:0] t_r8_c32_10;
  wire [7:0] t_r8_c32_11;
  wire [7:0] t_r8_c32_12;
  wire [7:0] t_r8_c33_0;
  wire [7:0] t_r8_c33_1;
  wire [7:0] t_r8_c33_2;
  wire [7:0] t_r8_c33_3;
  wire [7:0] t_r8_c33_4;
  wire [7:0] t_r8_c33_5;
  wire [7:0] t_r8_c33_6;
  wire [7:0] t_r8_c33_7;
  wire [7:0] t_r8_c33_8;
  wire [7:0] t_r8_c33_9;
  wire [7:0] t_r8_c33_10;
  wire [7:0] t_r8_c33_11;
  wire [7:0] t_r8_c33_12;
  wire [7:0] t_r8_c34_0;
  wire [7:0] t_r8_c34_1;
  wire [7:0] t_r8_c34_2;
  wire [7:0] t_r8_c34_3;
  wire [7:0] t_r8_c34_4;
  wire [7:0] t_r8_c34_5;
  wire [7:0] t_r8_c34_6;
  wire [7:0] t_r8_c34_7;
  wire [7:0] t_r8_c34_8;
  wire [7:0] t_r8_c34_9;
  wire [7:0] t_r8_c34_10;
  wire [7:0] t_r8_c34_11;
  wire [7:0] t_r8_c34_12;
  wire [7:0] t_r8_c35_0;
  wire [7:0] t_r8_c35_1;
  wire [7:0] t_r8_c35_2;
  wire [7:0] t_r8_c35_3;
  wire [7:0] t_r8_c35_4;
  wire [7:0] t_r8_c35_5;
  wire [7:0] t_r8_c35_6;
  wire [7:0] t_r8_c35_7;
  wire [7:0] t_r8_c35_8;
  wire [7:0] t_r8_c35_9;
  wire [7:0] t_r8_c35_10;
  wire [7:0] t_r8_c35_11;
  wire [7:0] t_r8_c35_12;
  wire [7:0] t_r8_c36_0;
  wire [7:0] t_r8_c36_1;
  wire [7:0] t_r8_c36_2;
  wire [7:0] t_r8_c36_3;
  wire [7:0] t_r8_c36_4;
  wire [7:0] t_r8_c36_5;
  wire [7:0] t_r8_c36_6;
  wire [7:0] t_r8_c36_7;
  wire [7:0] t_r8_c36_8;
  wire [7:0] t_r8_c36_9;
  wire [7:0] t_r8_c36_10;
  wire [7:0] t_r8_c36_11;
  wire [7:0] t_r8_c36_12;
  wire [7:0] t_r8_c37_0;
  wire [7:0] t_r8_c37_1;
  wire [7:0] t_r8_c37_2;
  wire [7:0] t_r8_c37_3;
  wire [7:0] t_r8_c37_4;
  wire [7:0] t_r8_c37_5;
  wire [7:0] t_r8_c37_6;
  wire [7:0] t_r8_c37_7;
  wire [7:0] t_r8_c37_8;
  wire [7:0] t_r8_c37_9;
  wire [7:0] t_r8_c37_10;
  wire [7:0] t_r8_c37_11;
  wire [7:0] t_r8_c37_12;
  wire [7:0] t_r8_c38_0;
  wire [7:0] t_r8_c38_1;
  wire [7:0] t_r8_c38_2;
  wire [7:0] t_r8_c38_3;
  wire [7:0] t_r8_c38_4;
  wire [7:0] t_r8_c38_5;
  wire [7:0] t_r8_c38_6;
  wire [7:0] t_r8_c38_7;
  wire [7:0] t_r8_c38_8;
  wire [7:0] t_r8_c38_9;
  wire [7:0] t_r8_c38_10;
  wire [7:0] t_r8_c38_11;
  wire [7:0] t_r8_c38_12;
  wire [7:0] t_r8_c39_0;
  wire [7:0] t_r8_c39_1;
  wire [7:0] t_r8_c39_2;
  wire [7:0] t_r8_c39_3;
  wire [7:0] t_r8_c39_4;
  wire [7:0] t_r8_c39_5;
  wire [7:0] t_r8_c39_6;
  wire [7:0] t_r8_c39_7;
  wire [7:0] t_r8_c39_8;
  wire [7:0] t_r8_c39_9;
  wire [7:0] t_r8_c39_10;
  wire [7:0] t_r8_c39_11;
  wire [7:0] t_r8_c39_12;
  wire [7:0] t_r8_c40_0;
  wire [7:0] t_r8_c40_1;
  wire [7:0] t_r8_c40_2;
  wire [7:0] t_r8_c40_3;
  wire [7:0] t_r8_c40_4;
  wire [7:0] t_r8_c40_5;
  wire [7:0] t_r8_c40_6;
  wire [7:0] t_r8_c40_7;
  wire [7:0] t_r8_c40_8;
  wire [7:0] t_r8_c40_9;
  wire [7:0] t_r8_c40_10;
  wire [7:0] t_r8_c40_11;
  wire [7:0] t_r8_c40_12;
  wire [7:0] t_r8_c41_0;
  wire [7:0] t_r8_c41_1;
  wire [7:0] t_r8_c41_2;
  wire [7:0] t_r8_c41_3;
  wire [7:0] t_r8_c41_4;
  wire [7:0] t_r8_c41_5;
  wire [7:0] t_r8_c41_6;
  wire [7:0] t_r8_c41_7;
  wire [7:0] t_r8_c41_8;
  wire [7:0] t_r8_c41_9;
  wire [7:0] t_r8_c41_10;
  wire [7:0] t_r8_c41_11;
  wire [7:0] t_r8_c41_12;
  wire [7:0] t_r8_c42_0;
  wire [7:0] t_r8_c42_1;
  wire [7:0] t_r8_c42_2;
  wire [7:0] t_r8_c42_3;
  wire [7:0] t_r8_c42_4;
  wire [7:0] t_r8_c42_5;
  wire [7:0] t_r8_c42_6;
  wire [7:0] t_r8_c42_7;
  wire [7:0] t_r8_c42_8;
  wire [7:0] t_r8_c42_9;
  wire [7:0] t_r8_c42_10;
  wire [7:0] t_r8_c42_11;
  wire [7:0] t_r8_c42_12;
  wire [7:0] t_r8_c43_0;
  wire [7:0] t_r8_c43_1;
  wire [7:0] t_r8_c43_2;
  wire [7:0] t_r8_c43_3;
  wire [7:0] t_r8_c43_4;
  wire [7:0] t_r8_c43_5;
  wire [7:0] t_r8_c43_6;
  wire [7:0] t_r8_c43_7;
  wire [7:0] t_r8_c43_8;
  wire [7:0] t_r8_c43_9;
  wire [7:0] t_r8_c43_10;
  wire [7:0] t_r8_c43_11;
  wire [7:0] t_r8_c43_12;
  wire [7:0] t_r8_c44_0;
  wire [7:0] t_r8_c44_1;
  wire [7:0] t_r8_c44_2;
  wire [7:0] t_r8_c44_3;
  wire [7:0] t_r8_c44_4;
  wire [7:0] t_r8_c44_5;
  wire [7:0] t_r8_c44_6;
  wire [7:0] t_r8_c44_7;
  wire [7:0] t_r8_c44_8;
  wire [7:0] t_r8_c44_9;
  wire [7:0] t_r8_c44_10;
  wire [7:0] t_r8_c44_11;
  wire [7:0] t_r8_c44_12;
  wire [7:0] t_r8_c45_0;
  wire [7:0] t_r8_c45_1;
  wire [7:0] t_r8_c45_2;
  wire [7:0] t_r8_c45_3;
  wire [7:0] t_r8_c45_4;
  wire [7:0] t_r8_c45_5;
  wire [7:0] t_r8_c45_6;
  wire [7:0] t_r8_c45_7;
  wire [7:0] t_r8_c45_8;
  wire [7:0] t_r8_c45_9;
  wire [7:0] t_r8_c45_10;
  wire [7:0] t_r8_c45_11;
  wire [7:0] t_r8_c45_12;
  wire [7:0] t_r8_c46_0;
  wire [7:0] t_r8_c46_1;
  wire [7:0] t_r8_c46_2;
  wire [7:0] t_r8_c46_3;
  wire [7:0] t_r8_c46_4;
  wire [7:0] t_r8_c46_5;
  wire [7:0] t_r8_c46_6;
  wire [7:0] t_r8_c46_7;
  wire [7:0] t_r8_c46_8;
  wire [7:0] t_r8_c46_9;
  wire [7:0] t_r8_c46_10;
  wire [7:0] t_r8_c46_11;
  wire [7:0] t_r8_c46_12;
  wire [7:0] t_r8_c47_0;
  wire [7:0] t_r8_c47_1;
  wire [7:0] t_r8_c47_2;
  wire [7:0] t_r8_c47_3;
  wire [7:0] t_r8_c47_4;
  wire [7:0] t_r8_c47_5;
  wire [7:0] t_r8_c47_6;
  wire [7:0] t_r8_c47_7;
  wire [7:0] t_r8_c47_8;
  wire [7:0] t_r8_c47_9;
  wire [7:0] t_r8_c47_10;
  wire [7:0] t_r8_c47_11;
  wire [7:0] t_r8_c47_12;
  wire [7:0] t_r8_c48_0;
  wire [7:0] t_r8_c48_1;
  wire [7:0] t_r8_c48_2;
  wire [7:0] t_r8_c48_3;
  wire [7:0] t_r8_c48_4;
  wire [7:0] t_r8_c48_5;
  wire [7:0] t_r8_c48_6;
  wire [7:0] t_r8_c48_7;
  wire [7:0] t_r8_c48_8;
  wire [7:0] t_r8_c48_9;
  wire [7:0] t_r8_c48_10;
  wire [7:0] t_r8_c48_11;
  wire [7:0] t_r8_c48_12;
  wire [7:0] t_r8_c49_0;
  wire [7:0] t_r8_c49_1;
  wire [7:0] t_r8_c49_2;
  wire [7:0] t_r8_c49_3;
  wire [7:0] t_r8_c49_4;
  wire [7:0] t_r8_c49_5;
  wire [7:0] t_r8_c49_6;
  wire [7:0] t_r8_c49_7;
  wire [7:0] t_r8_c49_8;
  wire [7:0] t_r8_c49_9;
  wire [7:0] t_r8_c49_10;
  wire [7:0] t_r8_c49_11;
  wire [7:0] t_r8_c49_12;
  wire [7:0] t_r8_c50_0;
  wire [7:0] t_r8_c50_1;
  wire [7:0] t_r8_c50_2;
  wire [7:0] t_r8_c50_3;
  wire [7:0] t_r8_c50_4;
  wire [7:0] t_r8_c50_5;
  wire [7:0] t_r8_c50_6;
  wire [7:0] t_r8_c50_7;
  wire [7:0] t_r8_c50_8;
  wire [7:0] t_r8_c50_9;
  wire [7:0] t_r8_c50_10;
  wire [7:0] t_r8_c50_11;
  wire [7:0] t_r8_c50_12;
  wire [7:0] t_r8_c51_0;
  wire [7:0] t_r8_c51_1;
  wire [7:0] t_r8_c51_2;
  wire [7:0] t_r8_c51_3;
  wire [7:0] t_r8_c51_4;
  wire [7:0] t_r8_c51_5;
  wire [7:0] t_r8_c51_6;
  wire [7:0] t_r8_c51_7;
  wire [7:0] t_r8_c51_8;
  wire [7:0] t_r8_c51_9;
  wire [7:0] t_r8_c51_10;
  wire [7:0] t_r8_c51_11;
  wire [7:0] t_r8_c51_12;
  wire [7:0] t_r8_c52_0;
  wire [7:0] t_r8_c52_1;
  wire [7:0] t_r8_c52_2;
  wire [7:0] t_r8_c52_3;
  wire [7:0] t_r8_c52_4;
  wire [7:0] t_r8_c52_5;
  wire [7:0] t_r8_c52_6;
  wire [7:0] t_r8_c52_7;
  wire [7:0] t_r8_c52_8;
  wire [7:0] t_r8_c52_9;
  wire [7:0] t_r8_c52_10;
  wire [7:0] t_r8_c52_11;
  wire [7:0] t_r8_c52_12;
  wire [7:0] t_r8_c53_0;
  wire [7:0] t_r8_c53_1;
  wire [7:0] t_r8_c53_2;
  wire [7:0] t_r8_c53_3;
  wire [7:0] t_r8_c53_4;
  wire [7:0] t_r8_c53_5;
  wire [7:0] t_r8_c53_6;
  wire [7:0] t_r8_c53_7;
  wire [7:0] t_r8_c53_8;
  wire [7:0] t_r8_c53_9;
  wire [7:0] t_r8_c53_10;
  wire [7:0] t_r8_c53_11;
  wire [7:0] t_r8_c53_12;
  wire [7:0] t_r8_c54_0;
  wire [7:0] t_r8_c54_1;
  wire [7:0] t_r8_c54_2;
  wire [7:0] t_r8_c54_3;
  wire [7:0] t_r8_c54_4;
  wire [7:0] t_r8_c54_5;
  wire [7:0] t_r8_c54_6;
  wire [7:0] t_r8_c54_7;
  wire [7:0] t_r8_c54_8;
  wire [7:0] t_r8_c54_9;
  wire [7:0] t_r8_c54_10;
  wire [7:0] t_r8_c54_11;
  wire [7:0] t_r8_c54_12;
  wire [7:0] t_r8_c55_0;
  wire [7:0] t_r8_c55_1;
  wire [7:0] t_r8_c55_2;
  wire [7:0] t_r8_c55_3;
  wire [7:0] t_r8_c55_4;
  wire [7:0] t_r8_c55_5;
  wire [7:0] t_r8_c55_6;
  wire [7:0] t_r8_c55_7;
  wire [7:0] t_r8_c55_8;
  wire [7:0] t_r8_c55_9;
  wire [7:0] t_r8_c55_10;
  wire [7:0] t_r8_c55_11;
  wire [7:0] t_r8_c55_12;
  wire [7:0] t_r8_c56_0;
  wire [7:0] t_r8_c56_1;
  wire [7:0] t_r8_c56_2;
  wire [7:0] t_r8_c56_3;
  wire [7:0] t_r8_c56_4;
  wire [7:0] t_r8_c56_5;
  wire [7:0] t_r8_c56_6;
  wire [7:0] t_r8_c56_7;
  wire [7:0] t_r8_c56_8;
  wire [7:0] t_r8_c56_9;
  wire [7:0] t_r8_c56_10;
  wire [7:0] t_r8_c56_11;
  wire [7:0] t_r8_c56_12;
  wire [7:0] t_r8_c57_0;
  wire [7:0] t_r8_c57_1;
  wire [7:0] t_r8_c57_2;
  wire [7:0] t_r8_c57_3;
  wire [7:0] t_r8_c57_4;
  wire [7:0] t_r8_c57_5;
  wire [7:0] t_r8_c57_6;
  wire [7:0] t_r8_c57_7;
  wire [7:0] t_r8_c57_8;
  wire [7:0] t_r8_c57_9;
  wire [7:0] t_r8_c57_10;
  wire [7:0] t_r8_c57_11;
  wire [7:0] t_r8_c57_12;
  wire [7:0] t_r8_c58_0;
  wire [7:0] t_r8_c58_1;
  wire [7:0] t_r8_c58_2;
  wire [7:0] t_r8_c58_3;
  wire [7:0] t_r8_c58_4;
  wire [7:0] t_r8_c58_5;
  wire [7:0] t_r8_c58_6;
  wire [7:0] t_r8_c58_7;
  wire [7:0] t_r8_c58_8;
  wire [7:0] t_r8_c58_9;
  wire [7:0] t_r8_c58_10;
  wire [7:0] t_r8_c58_11;
  wire [7:0] t_r8_c58_12;
  wire [7:0] t_r8_c59_0;
  wire [7:0] t_r8_c59_1;
  wire [7:0] t_r8_c59_2;
  wire [7:0] t_r8_c59_3;
  wire [7:0] t_r8_c59_4;
  wire [7:0] t_r8_c59_5;
  wire [7:0] t_r8_c59_6;
  wire [7:0] t_r8_c59_7;
  wire [7:0] t_r8_c59_8;
  wire [7:0] t_r8_c59_9;
  wire [7:0] t_r8_c59_10;
  wire [7:0] t_r8_c59_11;
  wire [7:0] t_r8_c59_12;
  wire [7:0] t_r8_c60_0;
  wire [7:0] t_r8_c60_1;
  wire [7:0] t_r8_c60_2;
  wire [7:0] t_r8_c60_3;
  wire [7:0] t_r8_c60_4;
  wire [7:0] t_r8_c60_5;
  wire [7:0] t_r8_c60_6;
  wire [7:0] t_r8_c60_7;
  wire [7:0] t_r8_c60_8;
  wire [7:0] t_r8_c60_9;
  wire [7:0] t_r8_c60_10;
  wire [7:0] t_r8_c60_11;
  wire [7:0] t_r8_c60_12;
  wire [7:0] t_r8_c61_0;
  wire [7:0] t_r8_c61_1;
  wire [7:0] t_r8_c61_2;
  wire [7:0] t_r8_c61_3;
  wire [7:0] t_r8_c61_4;
  wire [7:0] t_r8_c61_5;
  wire [7:0] t_r8_c61_6;
  wire [7:0] t_r8_c61_7;
  wire [7:0] t_r8_c61_8;
  wire [7:0] t_r8_c61_9;
  wire [7:0] t_r8_c61_10;
  wire [7:0] t_r8_c61_11;
  wire [7:0] t_r8_c61_12;
  wire [7:0] t_r8_c62_0;
  wire [7:0] t_r8_c62_1;
  wire [7:0] t_r8_c62_2;
  wire [7:0] t_r8_c62_3;
  wire [7:0] t_r8_c62_4;
  wire [7:0] t_r8_c62_5;
  wire [7:0] t_r8_c62_6;
  wire [7:0] t_r8_c62_7;
  wire [7:0] t_r8_c62_8;
  wire [7:0] t_r8_c62_9;
  wire [7:0] t_r8_c62_10;
  wire [7:0] t_r8_c62_11;
  wire [7:0] t_r8_c62_12;
  wire [7:0] t_r8_c63_0;
  wire [7:0] t_r8_c63_1;
  wire [7:0] t_r8_c63_2;
  wire [7:0] t_r8_c63_3;
  wire [7:0] t_r8_c63_4;
  wire [7:0] t_r8_c63_5;
  wire [7:0] t_r8_c63_6;
  wire [7:0] t_r8_c63_7;
  wire [7:0] t_r8_c63_8;
  wire [7:0] t_r8_c63_9;
  wire [7:0] t_r8_c63_10;
  wire [7:0] t_r8_c63_11;
  wire [7:0] t_r8_c63_12;
  wire [7:0] t_r8_c64_0;
  wire [7:0] t_r8_c64_1;
  wire [7:0] t_r8_c64_2;
  wire [7:0] t_r8_c64_3;
  wire [7:0] t_r8_c64_4;
  wire [7:0] t_r8_c64_5;
  wire [7:0] t_r8_c64_6;
  wire [7:0] t_r8_c64_7;
  wire [7:0] t_r8_c64_8;
  wire [7:0] t_r8_c64_9;
  wire [7:0] t_r8_c64_10;
  wire [7:0] t_r8_c64_11;
  wire [7:0] t_r8_c64_12;
  wire [7:0] t_r8_c65_0;
  wire [7:0] t_r8_c65_1;
  wire [7:0] t_r8_c65_2;
  wire [7:0] t_r8_c65_3;
  wire [7:0] t_r8_c65_4;
  wire [7:0] t_r8_c65_5;
  wire [7:0] t_r8_c65_6;
  wire [7:0] t_r8_c65_7;
  wire [7:0] t_r8_c65_8;
  wire [7:0] t_r8_c65_9;
  wire [7:0] t_r8_c65_10;
  wire [7:0] t_r8_c65_11;
  wire [7:0] t_r8_c65_12;
  wire [7:0] t_r9_c0_0;
  wire [7:0] t_r9_c0_1;
  wire [7:0] t_r9_c0_2;
  wire [7:0] t_r9_c0_3;
  wire [7:0] t_r9_c0_4;
  wire [7:0] t_r9_c0_5;
  wire [7:0] t_r9_c0_6;
  wire [7:0] t_r9_c0_7;
  wire [7:0] t_r9_c0_8;
  wire [7:0] t_r9_c0_9;
  wire [7:0] t_r9_c0_10;
  wire [7:0] t_r9_c0_11;
  wire [7:0] t_r9_c0_12;
  wire [7:0] t_r9_c1_0;
  wire [7:0] t_r9_c1_1;
  wire [7:0] t_r9_c1_2;
  wire [7:0] t_r9_c1_3;
  wire [7:0] t_r9_c1_4;
  wire [7:0] t_r9_c1_5;
  wire [7:0] t_r9_c1_6;
  wire [7:0] t_r9_c1_7;
  wire [7:0] t_r9_c1_8;
  wire [7:0] t_r9_c1_9;
  wire [7:0] t_r9_c1_10;
  wire [7:0] t_r9_c1_11;
  wire [7:0] t_r9_c1_12;
  wire [7:0] t_r9_c2_0;
  wire [7:0] t_r9_c2_1;
  wire [7:0] t_r9_c2_2;
  wire [7:0] t_r9_c2_3;
  wire [7:0] t_r9_c2_4;
  wire [7:0] t_r9_c2_5;
  wire [7:0] t_r9_c2_6;
  wire [7:0] t_r9_c2_7;
  wire [7:0] t_r9_c2_8;
  wire [7:0] t_r9_c2_9;
  wire [7:0] t_r9_c2_10;
  wire [7:0] t_r9_c2_11;
  wire [7:0] t_r9_c2_12;
  wire [7:0] t_r9_c3_0;
  wire [7:0] t_r9_c3_1;
  wire [7:0] t_r9_c3_2;
  wire [7:0] t_r9_c3_3;
  wire [7:0] t_r9_c3_4;
  wire [7:0] t_r9_c3_5;
  wire [7:0] t_r9_c3_6;
  wire [7:0] t_r9_c3_7;
  wire [7:0] t_r9_c3_8;
  wire [7:0] t_r9_c3_9;
  wire [7:0] t_r9_c3_10;
  wire [7:0] t_r9_c3_11;
  wire [7:0] t_r9_c3_12;
  wire [7:0] t_r9_c4_0;
  wire [7:0] t_r9_c4_1;
  wire [7:0] t_r9_c4_2;
  wire [7:0] t_r9_c4_3;
  wire [7:0] t_r9_c4_4;
  wire [7:0] t_r9_c4_5;
  wire [7:0] t_r9_c4_6;
  wire [7:0] t_r9_c4_7;
  wire [7:0] t_r9_c4_8;
  wire [7:0] t_r9_c4_9;
  wire [7:0] t_r9_c4_10;
  wire [7:0] t_r9_c4_11;
  wire [7:0] t_r9_c4_12;
  wire [7:0] t_r9_c5_0;
  wire [7:0] t_r9_c5_1;
  wire [7:0] t_r9_c5_2;
  wire [7:0] t_r9_c5_3;
  wire [7:0] t_r9_c5_4;
  wire [7:0] t_r9_c5_5;
  wire [7:0] t_r9_c5_6;
  wire [7:0] t_r9_c5_7;
  wire [7:0] t_r9_c5_8;
  wire [7:0] t_r9_c5_9;
  wire [7:0] t_r9_c5_10;
  wire [7:0] t_r9_c5_11;
  wire [7:0] t_r9_c5_12;
  wire [7:0] t_r9_c6_0;
  wire [7:0] t_r9_c6_1;
  wire [7:0] t_r9_c6_2;
  wire [7:0] t_r9_c6_3;
  wire [7:0] t_r9_c6_4;
  wire [7:0] t_r9_c6_5;
  wire [7:0] t_r9_c6_6;
  wire [7:0] t_r9_c6_7;
  wire [7:0] t_r9_c6_8;
  wire [7:0] t_r9_c6_9;
  wire [7:0] t_r9_c6_10;
  wire [7:0] t_r9_c6_11;
  wire [7:0] t_r9_c6_12;
  wire [7:0] t_r9_c7_0;
  wire [7:0] t_r9_c7_1;
  wire [7:0] t_r9_c7_2;
  wire [7:0] t_r9_c7_3;
  wire [7:0] t_r9_c7_4;
  wire [7:0] t_r9_c7_5;
  wire [7:0] t_r9_c7_6;
  wire [7:0] t_r9_c7_7;
  wire [7:0] t_r9_c7_8;
  wire [7:0] t_r9_c7_9;
  wire [7:0] t_r9_c7_10;
  wire [7:0] t_r9_c7_11;
  wire [7:0] t_r9_c7_12;
  wire [7:0] t_r9_c8_0;
  wire [7:0] t_r9_c8_1;
  wire [7:0] t_r9_c8_2;
  wire [7:0] t_r9_c8_3;
  wire [7:0] t_r9_c8_4;
  wire [7:0] t_r9_c8_5;
  wire [7:0] t_r9_c8_6;
  wire [7:0] t_r9_c8_7;
  wire [7:0] t_r9_c8_8;
  wire [7:0] t_r9_c8_9;
  wire [7:0] t_r9_c8_10;
  wire [7:0] t_r9_c8_11;
  wire [7:0] t_r9_c8_12;
  wire [7:0] t_r9_c9_0;
  wire [7:0] t_r9_c9_1;
  wire [7:0] t_r9_c9_2;
  wire [7:0] t_r9_c9_3;
  wire [7:0] t_r9_c9_4;
  wire [7:0] t_r9_c9_5;
  wire [7:0] t_r9_c9_6;
  wire [7:0] t_r9_c9_7;
  wire [7:0] t_r9_c9_8;
  wire [7:0] t_r9_c9_9;
  wire [7:0] t_r9_c9_10;
  wire [7:0] t_r9_c9_11;
  wire [7:0] t_r9_c9_12;
  wire [7:0] t_r9_c10_0;
  wire [7:0] t_r9_c10_1;
  wire [7:0] t_r9_c10_2;
  wire [7:0] t_r9_c10_3;
  wire [7:0] t_r9_c10_4;
  wire [7:0] t_r9_c10_5;
  wire [7:0] t_r9_c10_6;
  wire [7:0] t_r9_c10_7;
  wire [7:0] t_r9_c10_8;
  wire [7:0] t_r9_c10_9;
  wire [7:0] t_r9_c10_10;
  wire [7:0] t_r9_c10_11;
  wire [7:0] t_r9_c10_12;
  wire [7:0] t_r9_c11_0;
  wire [7:0] t_r9_c11_1;
  wire [7:0] t_r9_c11_2;
  wire [7:0] t_r9_c11_3;
  wire [7:0] t_r9_c11_4;
  wire [7:0] t_r9_c11_5;
  wire [7:0] t_r9_c11_6;
  wire [7:0] t_r9_c11_7;
  wire [7:0] t_r9_c11_8;
  wire [7:0] t_r9_c11_9;
  wire [7:0] t_r9_c11_10;
  wire [7:0] t_r9_c11_11;
  wire [7:0] t_r9_c11_12;
  wire [7:0] t_r9_c12_0;
  wire [7:0] t_r9_c12_1;
  wire [7:0] t_r9_c12_2;
  wire [7:0] t_r9_c12_3;
  wire [7:0] t_r9_c12_4;
  wire [7:0] t_r9_c12_5;
  wire [7:0] t_r9_c12_6;
  wire [7:0] t_r9_c12_7;
  wire [7:0] t_r9_c12_8;
  wire [7:0] t_r9_c12_9;
  wire [7:0] t_r9_c12_10;
  wire [7:0] t_r9_c12_11;
  wire [7:0] t_r9_c12_12;
  wire [7:0] t_r9_c13_0;
  wire [7:0] t_r9_c13_1;
  wire [7:0] t_r9_c13_2;
  wire [7:0] t_r9_c13_3;
  wire [7:0] t_r9_c13_4;
  wire [7:0] t_r9_c13_5;
  wire [7:0] t_r9_c13_6;
  wire [7:0] t_r9_c13_7;
  wire [7:0] t_r9_c13_8;
  wire [7:0] t_r9_c13_9;
  wire [7:0] t_r9_c13_10;
  wire [7:0] t_r9_c13_11;
  wire [7:0] t_r9_c13_12;
  wire [7:0] t_r9_c14_0;
  wire [7:0] t_r9_c14_1;
  wire [7:0] t_r9_c14_2;
  wire [7:0] t_r9_c14_3;
  wire [7:0] t_r9_c14_4;
  wire [7:0] t_r9_c14_5;
  wire [7:0] t_r9_c14_6;
  wire [7:0] t_r9_c14_7;
  wire [7:0] t_r9_c14_8;
  wire [7:0] t_r9_c14_9;
  wire [7:0] t_r9_c14_10;
  wire [7:0] t_r9_c14_11;
  wire [7:0] t_r9_c14_12;
  wire [7:0] t_r9_c15_0;
  wire [7:0] t_r9_c15_1;
  wire [7:0] t_r9_c15_2;
  wire [7:0] t_r9_c15_3;
  wire [7:0] t_r9_c15_4;
  wire [7:0] t_r9_c15_5;
  wire [7:0] t_r9_c15_6;
  wire [7:0] t_r9_c15_7;
  wire [7:0] t_r9_c15_8;
  wire [7:0] t_r9_c15_9;
  wire [7:0] t_r9_c15_10;
  wire [7:0] t_r9_c15_11;
  wire [7:0] t_r9_c15_12;
  wire [7:0] t_r9_c16_0;
  wire [7:0] t_r9_c16_1;
  wire [7:0] t_r9_c16_2;
  wire [7:0] t_r9_c16_3;
  wire [7:0] t_r9_c16_4;
  wire [7:0] t_r9_c16_5;
  wire [7:0] t_r9_c16_6;
  wire [7:0] t_r9_c16_7;
  wire [7:0] t_r9_c16_8;
  wire [7:0] t_r9_c16_9;
  wire [7:0] t_r9_c16_10;
  wire [7:0] t_r9_c16_11;
  wire [7:0] t_r9_c16_12;
  wire [7:0] t_r9_c17_0;
  wire [7:0] t_r9_c17_1;
  wire [7:0] t_r9_c17_2;
  wire [7:0] t_r9_c17_3;
  wire [7:0] t_r9_c17_4;
  wire [7:0] t_r9_c17_5;
  wire [7:0] t_r9_c17_6;
  wire [7:0] t_r9_c17_7;
  wire [7:0] t_r9_c17_8;
  wire [7:0] t_r9_c17_9;
  wire [7:0] t_r9_c17_10;
  wire [7:0] t_r9_c17_11;
  wire [7:0] t_r9_c17_12;
  wire [7:0] t_r9_c18_0;
  wire [7:0] t_r9_c18_1;
  wire [7:0] t_r9_c18_2;
  wire [7:0] t_r9_c18_3;
  wire [7:0] t_r9_c18_4;
  wire [7:0] t_r9_c18_5;
  wire [7:0] t_r9_c18_6;
  wire [7:0] t_r9_c18_7;
  wire [7:0] t_r9_c18_8;
  wire [7:0] t_r9_c18_9;
  wire [7:0] t_r9_c18_10;
  wire [7:0] t_r9_c18_11;
  wire [7:0] t_r9_c18_12;
  wire [7:0] t_r9_c19_0;
  wire [7:0] t_r9_c19_1;
  wire [7:0] t_r9_c19_2;
  wire [7:0] t_r9_c19_3;
  wire [7:0] t_r9_c19_4;
  wire [7:0] t_r9_c19_5;
  wire [7:0] t_r9_c19_6;
  wire [7:0] t_r9_c19_7;
  wire [7:0] t_r9_c19_8;
  wire [7:0] t_r9_c19_9;
  wire [7:0] t_r9_c19_10;
  wire [7:0] t_r9_c19_11;
  wire [7:0] t_r9_c19_12;
  wire [7:0] t_r9_c20_0;
  wire [7:0] t_r9_c20_1;
  wire [7:0] t_r9_c20_2;
  wire [7:0] t_r9_c20_3;
  wire [7:0] t_r9_c20_4;
  wire [7:0] t_r9_c20_5;
  wire [7:0] t_r9_c20_6;
  wire [7:0] t_r9_c20_7;
  wire [7:0] t_r9_c20_8;
  wire [7:0] t_r9_c20_9;
  wire [7:0] t_r9_c20_10;
  wire [7:0] t_r9_c20_11;
  wire [7:0] t_r9_c20_12;
  wire [7:0] t_r9_c21_0;
  wire [7:0] t_r9_c21_1;
  wire [7:0] t_r9_c21_2;
  wire [7:0] t_r9_c21_3;
  wire [7:0] t_r9_c21_4;
  wire [7:0] t_r9_c21_5;
  wire [7:0] t_r9_c21_6;
  wire [7:0] t_r9_c21_7;
  wire [7:0] t_r9_c21_8;
  wire [7:0] t_r9_c21_9;
  wire [7:0] t_r9_c21_10;
  wire [7:0] t_r9_c21_11;
  wire [7:0] t_r9_c21_12;
  wire [7:0] t_r9_c22_0;
  wire [7:0] t_r9_c22_1;
  wire [7:0] t_r9_c22_2;
  wire [7:0] t_r9_c22_3;
  wire [7:0] t_r9_c22_4;
  wire [7:0] t_r9_c22_5;
  wire [7:0] t_r9_c22_6;
  wire [7:0] t_r9_c22_7;
  wire [7:0] t_r9_c22_8;
  wire [7:0] t_r9_c22_9;
  wire [7:0] t_r9_c22_10;
  wire [7:0] t_r9_c22_11;
  wire [7:0] t_r9_c22_12;
  wire [7:0] t_r9_c23_0;
  wire [7:0] t_r9_c23_1;
  wire [7:0] t_r9_c23_2;
  wire [7:0] t_r9_c23_3;
  wire [7:0] t_r9_c23_4;
  wire [7:0] t_r9_c23_5;
  wire [7:0] t_r9_c23_6;
  wire [7:0] t_r9_c23_7;
  wire [7:0] t_r9_c23_8;
  wire [7:0] t_r9_c23_9;
  wire [7:0] t_r9_c23_10;
  wire [7:0] t_r9_c23_11;
  wire [7:0] t_r9_c23_12;
  wire [7:0] t_r9_c24_0;
  wire [7:0] t_r9_c24_1;
  wire [7:0] t_r9_c24_2;
  wire [7:0] t_r9_c24_3;
  wire [7:0] t_r9_c24_4;
  wire [7:0] t_r9_c24_5;
  wire [7:0] t_r9_c24_6;
  wire [7:0] t_r9_c24_7;
  wire [7:0] t_r9_c24_8;
  wire [7:0] t_r9_c24_9;
  wire [7:0] t_r9_c24_10;
  wire [7:0] t_r9_c24_11;
  wire [7:0] t_r9_c24_12;
  wire [7:0] t_r9_c25_0;
  wire [7:0] t_r9_c25_1;
  wire [7:0] t_r9_c25_2;
  wire [7:0] t_r9_c25_3;
  wire [7:0] t_r9_c25_4;
  wire [7:0] t_r9_c25_5;
  wire [7:0] t_r9_c25_6;
  wire [7:0] t_r9_c25_7;
  wire [7:0] t_r9_c25_8;
  wire [7:0] t_r9_c25_9;
  wire [7:0] t_r9_c25_10;
  wire [7:0] t_r9_c25_11;
  wire [7:0] t_r9_c25_12;
  wire [7:0] t_r9_c26_0;
  wire [7:0] t_r9_c26_1;
  wire [7:0] t_r9_c26_2;
  wire [7:0] t_r9_c26_3;
  wire [7:0] t_r9_c26_4;
  wire [7:0] t_r9_c26_5;
  wire [7:0] t_r9_c26_6;
  wire [7:0] t_r9_c26_7;
  wire [7:0] t_r9_c26_8;
  wire [7:0] t_r9_c26_9;
  wire [7:0] t_r9_c26_10;
  wire [7:0] t_r9_c26_11;
  wire [7:0] t_r9_c26_12;
  wire [7:0] t_r9_c27_0;
  wire [7:0] t_r9_c27_1;
  wire [7:0] t_r9_c27_2;
  wire [7:0] t_r9_c27_3;
  wire [7:0] t_r9_c27_4;
  wire [7:0] t_r9_c27_5;
  wire [7:0] t_r9_c27_6;
  wire [7:0] t_r9_c27_7;
  wire [7:0] t_r9_c27_8;
  wire [7:0] t_r9_c27_9;
  wire [7:0] t_r9_c27_10;
  wire [7:0] t_r9_c27_11;
  wire [7:0] t_r9_c27_12;
  wire [7:0] t_r9_c28_0;
  wire [7:0] t_r9_c28_1;
  wire [7:0] t_r9_c28_2;
  wire [7:0] t_r9_c28_3;
  wire [7:0] t_r9_c28_4;
  wire [7:0] t_r9_c28_5;
  wire [7:0] t_r9_c28_6;
  wire [7:0] t_r9_c28_7;
  wire [7:0] t_r9_c28_8;
  wire [7:0] t_r9_c28_9;
  wire [7:0] t_r9_c28_10;
  wire [7:0] t_r9_c28_11;
  wire [7:0] t_r9_c28_12;
  wire [7:0] t_r9_c29_0;
  wire [7:0] t_r9_c29_1;
  wire [7:0] t_r9_c29_2;
  wire [7:0] t_r9_c29_3;
  wire [7:0] t_r9_c29_4;
  wire [7:0] t_r9_c29_5;
  wire [7:0] t_r9_c29_6;
  wire [7:0] t_r9_c29_7;
  wire [7:0] t_r9_c29_8;
  wire [7:0] t_r9_c29_9;
  wire [7:0] t_r9_c29_10;
  wire [7:0] t_r9_c29_11;
  wire [7:0] t_r9_c29_12;
  wire [7:0] t_r9_c30_0;
  wire [7:0] t_r9_c30_1;
  wire [7:0] t_r9_c30_2;
  wire [7:0] t_r9_c30_3;
  wire [7:0] t_r9_c30_4;
  wire [7:0] t_r9_c30_5;
  wire [7:0] t_r9_c30_6;
  wire [7:0] t_r9_c30_7;
  wire [7:0] t_r9_c30_8;
  wire [7:0] t_r9_c30_9;
  wire [7:0] t_r9_c30_10;
  wire [7:0] t_r9_c30_11;
  wire [7:0] t_r9_c30_12;
  wire [7:0] t_r9_c31_0;
  wire [7:0] t_r9_c31_1;
  wire [7:0] t_r9_c31_2;
  wire [7:0] t_r9_c31_3;
  wire [7:0] t_r9_c31_4;
  wire [7:0] t_r9_c31_5;
  wire [7:0] t_r9_c31_6;
  wire [7:0] t_r9_c31_7;
  wire [7:0] t_r9_c31_8;
  wire [7:0] t_r9_c31_9;
  wire [7:0] t_r9_c31_10;
  wire [7:0] t_r9_c31_11;
  wire [7:0] t_r9_c31_12;
  wire [7:0] t_r9_c32_0;
  wire [7:0] t_r9_c32_1;
  wire [7:0] t_r9_c32_2;
  wire [7:0] t_r9_c32_3;
  wire [7:0] t_r9_c32_4;
  wire [7:0] t_r9_c32_5;
  wire [7:0] t_r9_c32_6;
  wire [7:0] t_r9_c32_7;
  wire [7:0] t_r9_c32_8;
  wire [7:0] t_r9_c32_9;
  wire [7:0] t_r9_c32_10;
  wire [7:0] t_r9_c32_11;
  wire [7:0] t_r9_c32_12;
  wire [7:0] t_r9_c33_0;
  wire [7:0] t_r9_c33_1;
  wire [7:0] t_r9_c33_2;
  wire [7:0] t_r9_c33_3;
  wire [7:0] t_r9_c33_4;
  wire [7:0] t_r9_c33_5;
  wire [7:0] t_r9_c33_6;
  wire [7:0] t_r9_c33_7;
  wire [7:0] t_r9_c33_8;
  wire [7:0] t_r9_c33_9;
  wire [7:0] t_r9_c33_10;
  wire [7:0] t_r9_c33_11;
  wire [7:0] t_r9_c33_12;
  wire [7:0] t_r9_c34_0;
  wire [7:0] t_r9_c34_1;
  wire [7:0] t_r9_c34_2;
  wire [7:0] t_r9_c34_3;
  wire [7:0] t_r9_c34_4;
  wire [7:0] t_r9_c34_5;
  wire [7:0] t_r9_c34_6;
  wire [7:0] t_r9_c34_7;
  wire [7:0] t_r9_c34_8;
  wire [7:0] t_r9_c34_9;
  wire [7:0] t_r9_c34_10;
  wire [7:0] t_r9_c34_11;
  wire [7:0] t_r9_c34_12;
  wire [7:0] t_r9_c35_0;
  wire [7:0] t_r9_c35_1;
  wire [7:0] t_r9_c35_2;
  wire [7:0] t_r9_c35_3;
  wire [7:0] t_r9_c35_4;
  wire [7:0] t_r9_c35_5;
  wire [7:0] t_r9_c35_6;
  wire [7:0] t_r9_c35_7;
  wire [7:0] t_r9_c35_8;
  wire [7:0] t_r9_c35_9;
  wire [7:0] t_r9_c35_10;
  wire [7:0] t_r9_c35_11;
  wire [7:0] t_r9_c35_12;
  wire [7:0] t_r9_c36_0;
  wire [7:0] t_r9_c36_1;
  wire [7:0] t_r9_c36_2;
  wire [7:0] t_r9_c36_3;
  wire [7:0] t_r9_c36_4;
  wire [7:0] t_r9_c36_5;
  wire [7:0] t_r9_c36_6;
  wire [7:0] t_r9_c36_7;
  wire [7:0] t_r9_c36_8;
  wire [7:0] t_r9_c36_9;
  wire [7:0] t_r9_c36_10;
  wire [7:0] t_r9_c36_11;
  wire [7:0] t_r9_c36_12;
  wire [7:0] t_r9_c37_0;
  wire [7:0] t_r9_c37_1;
  wire [7:0] t_r9_c37_2;
  wire [7:0] t_r9_c37_3;
  wire [7:0] t_r9_c37_4;
  wire [7:0] t_r9_c37_5;
  wire [7:0] t_r9_c37_6;
  wire [7:0] t_r9_c37_7;
  wire [7:0] t_r9_c37_8;
  wire [7:0] t_r9_c37_9;
  wire [7:0] t_r9_c37_10;
  wire [7:0] t_r9_c37_11;
  wire [7:0] t_r9_c37_12;
  wire [7:0] t_r9_c38_0;
  wire [7:0] t_r9_c38_1;
  wire [7:0] t_r9_c38_2;
  wire [7:0] t_r9_c38_3;
  wire [7:0] t_r9_c38_4;
  wire [7:0] t_r9_c38_5;
  wire [7:0] t_r9_c38_6;
  wire [7:0] t_r9_c38_7;
  wire [7:0] t_r9_c38_8;
  wire [7:0] t_r9_c38_9;
  wire [7:0] t_r9_c38_10;
  wire [7:0] t_r9_c38_11;
  wire [7:0] t_r9_c38_12;
  wire [7:0] t_r9_c39_0;
  wire [7:0] t_r9_c39_1;
  wire [7:0] t_r9_c39_2;
  wire [7:0] t_r9_c39_3;
  wire [7:0] t_r9_c39_4;
  wire [7:0] t_r9_c39_5;
  wire [7:0] t_r9_c39_6;
  wire [7:0] t_r9_c39_7;
  wire [7:0] t_r9_c39_8;
  wire [7:0] t_r9_c39_9;
  wire [7:0] t_r9_c39_10;
  wire [7:0] t_r9_c39_11;
  wire [7:0] t_r9_c39_12;
  wire [7:0] t_r9_c40_0;
  wire [7:0] t_r9_c40_1;
  wire [7:0] t_r9_c40_2;
  wire [7:0] t_r9_c40_3;
  wire [7:0] t_r9_c40_4;
  wire [7:0] t_r9_c40_5;
  wire [7:0] t_r9_c40_6;
  wire [7:0] t_r9_c40_7;
  wire [7:0] t_r9_c40_8;
  wire [7:0] t_r9_c40_9;
  wire [7:0] t_r9_c40_10;
  wire [7:0] t_r9_c40_11;
  wire [7:0] t_r9_c40_12;
  wire [7:0] t_r9_c41_0;
  wire [7:0] t_r9_c41_1;
  wire [7:0] t_r9_c41_2;
  wire [7:0] t_r9_c41_3;
  wire [7:0] t_r9_c41_4;
  wire [7:0] t_r9_c41_5;
  wire [7:0] t_r9_c41_6;
  wire [7:0] t_r9_c41_7;
  wire [7:0] t_r9_c41_8;
  wire [7:0] t_r9_c41_9;
  wire [7:0] t_r9_c41_10;
  wire [7:0] t_r9_c41_11;
  wire [7:0] t_r9_c41_12;
  wire [7:0] t_r9_c42_0;
  wire [7:0] t_r9_c42_1;
  wire [7:0] t_r9_c42_2;
  wire [7:0] t_r9_c42_3;
  wire [7:0] t_r9_c42_4;
  wire [7:0] t_r9_c42_5;
  wire [7:0] t_r9_c42_6;
  wire [7:0] t_r9_c42_7;
  wire [7:0] t_r9_c42_8;
  wire [7:0] t_r9_c42_9;
  wire [7:0] t_r9_c42_10;
  wire [7:0] t_r9_c42_11;
  wire [7:0] t_r9_c42_12;
  wire [7:0] t_r9_c43_0;
  wire [7:0] t_r9_c43_1;
  wire [7:0] t_r9_c43_2;
  wire [7:0] t_r9_c43_3;
  wire [7:0] t_r9_c43_4;
  wire [7:0] t_r9_c43_5;
  wire [7:0] t_r9_c43_6;
  wire [7:0] t_r9_c43_7;
  wire [7:0] t_r9_c43_8;
  wire [7:0] t_r9_c43_9;
  wire [7:0] t_r9_c43_10;
  wire [7:0] t_r9_c43_11;
  wire [7:0] t_r9_c43_12;
  wire [7:0] t_r9_c44_0;
  wire [7:0] t_r9_c44_1;
  wire [7:0] t_r9_c44_2;
  wire [7:0] t_r9_c44_3;
  wire [7:0] t_r9_c44_4;
  wire [7:0] t_r9_c44_5;
  wire [7:0] t_r9_c44_6;
  wire [7:0] t_r9_c44_7;
  wire [7:0] t_r9_c44_8;
  wire [7:0] t_r9_c44_9;
  wire [7:0] t_r9_c44_10;
  wire [7:0] t_r9_c44_11;
  wire [7:0] t_r9_c44_12;
  wire [7:0] t_r9_c45_0;
  wire [7:0] t_r9_c45_1;
  wire [7:0] t_r9_c45_2;
  wire [7:0] t_r9_c45_3;
  wire [7:0] t_r9_c45_4;
  wire [7:0] t_r9_c45_5;
  wire [7:0] t_r9_c45_6;
  wire [7:0] t_r9_c45_7;
  wire [7:0] t_r9_c45_8;
  wire [7:0] t_r9_c45_9;
  wire [7:0] t_r9_c45_10;
  wire [7:0] t_r9_c45_11;
  wire [7:0] t_r9_c45_12;
  wire [7:0] t_r9_c46_0;
  wire [7:0] t_r9_c46_1;
  wire [7:0] t_r9_c46_2;
  wire [7:0] t_r9_c46_3;
  wire [7:0] t_r9_c46_4;
  wire [7:0] t_r9_c46_5;
  wire [7:0] t_r9_c46_6;
  wire [7:0] t_r9_c46_7;
  wire [7:0] t_r9_c46_8;
  wire [7:0] t_r9_c46_9;
  wire [7:0] t_r9_c46_10;
  wire [7:0] t_r9_c46_11;
  wire [7:0] t_r9_c46_12;
  wire [7:0] t_r9_c47_0;
  wire [7:0] t_r9_c47_1;
  wire [7:0] t_r9_c47_2;
  wire [7:0] t_r9_c47_3;
  wire [7:0] t_r9_c47_4;
  wire [7:0] t_r9_c47_5;
  wire [7:0] t_r9_c47_6;
  wire [7:0] t_r9_c47_7;
  wire [7:0] t_r9_c47_8;
  wire [7:0] t_r9_c47_9;
  wire [7:0] t_r9_c47_10;
  wire [7:0] t_r9_c47_11;
  wire [7:0] t_r9_c47_12;
  wire [7:0] t_r9_c48_0;
  wire [7:0] t_r9_c48_1;
  wire [7:0] t_r9_c48_2;
  wire [7:0] t_r9_c48_3;
  wire [7:0] t_r9_c48_4;
  wire [7:0] t_r9_c48_5;
  wire [7:0] t_r9_c48_6;
  wire [7:0] t_r9_c48_7;
  wire [7:0] t_r9_c48_8;
  wire [7:0] t_r9_c48_9;
  wire [7:0] t_r9_c48_10;
  wire [7:0] t_r9_c48_11;
  wire [7:0] t_r9_c48_12;
  wire [7:0] t_r9_c49_0;
  wire [7:0] t_r9_c49_1;
  wire [7:0] t_r9_c49_2;
  wire [7:0] t_r9_c49_3;
  wire [7:0] t_r9_c49_4;
  wire [7:0] t_r9_c49_5;
  wire [7:0] t_r9_c49_6;
  wire [7:0] t_r9_c49_7;
  wire [7:0] t_r9_c49_8;
  wire [7:0] t_r9_c49_9;
  wire [7:0] t_r9_c49_10;
  wire [7:0] t_r9_c49_11;
  wire [7:0] t_r9_c49_12;
  wire [7:0] t_r9_c50_0;
  wire [7:0] t_r9_c50_1;
  wire [7:0] t_r9_c50_2;
  wire [7:0] t_r9_c50_3;
  wire [7:0] t_r9_c50_4;
  wire [7:0] t_r9_c50_5;
  wire [7:0] t_r9_c50_6;
  wire [7:0] t_r9_c50_7;
  wire [7:0] t_r9_c50_8;
  wire [7:0] t_r9_c50_9;
  wire [7:0] t_r9_c50_10;
  wire [7:0] t_r9_c50_11;
  wire [7:0] t_r9_c50_12;
  wire [7:0] t_r9_c51_0;
  wire [7:0] t_r9_c51_1;
  wire [7:0] t_r9_c51_2;
  wire [7:0] t_r9_c51_3;
  wire [7:0] t_r9_c51_4;
  wire [7:0] t_r9_c51_5;
  wire [7:0] t_r9_c51_6;
  wire [7:0] t_r9_c51_7;
  wire [7:0] t_r9_c51_8;
  wire [7:0] t_r9_c51_9;
  wire [7:0] t_r9_c51_10;
  wire [7:0] t_r9_c51_11;
  wire [7:0] t_r9_c51_12;
  wire [7:0] t_r9_c52_0;
  wire [7:0] t_r9_c52_1;
  wire [7:0] t_r9_c52_2;
  wire [7:0] t_r9_c52_3;
  wire [7:0] t_r9_c52_4;
  wire [7:0] t_r9_c52_5;
  wire [7:0] t_r9_c52_6;
  wire [7:0] t_r9_c52_7;
  wire [7:0] t_r9_c52_8;
  wire [7:0] t_r9_c52_9;
  wire [7:0] t_r9_c52_10;
  wire [7:0] t_r9_c52_11;
  wire [7:0] t_r9_c52_12;
  wire [7:0] t_r9_c53_0;
  wire [7:0] t_r9_c53_1;
  wire [7:0] t_r9_c53_2;
  wire [7:0] t_r9_c53_3;
  wire [7:0] t_r9_c53_4;
  wire [7:0] t_r9_c53_5;
  wire [7:0] t_r9_c53_6;
  wire [7:0] t_r9_c53_7;
  wire [7:0] t_r9_c53_8;
  wire [7:0] t_r9_c53_9;
  wire [7:0] t_r9_c53_10;
  wire [7:0] t_r9_c53_11;
  wire [7:0] t_r9_c53_12;
  wire [7:0] t_r9_c54_0;
  wire [7:0] t_r9_c54_1;
  wire [7:0] t_r9_c54_2;
  wire [7:0] t_r9_c54_3;
  wire [7:0] t_r9_c54_4;
  wire [7:0] t_r9_c54_5;
  wire [7:0] t_r9_c54_6;
  wire [7:0] t_r9_c54_7;
  wire [7:0] t_r9_c54_8;
  wire [7:0] t_r9_c54_9;
  wire [7:0] t_r9_c54_10;
  wire [7:0] t_r9_c54_11;
  wire [7:0] t_r9_c54_12;
  wire [7:0] t_r9_c55_0;
  wire [7:0] t_r9_c55_1;
  wire [7:0] t_r9_c55_2;
  wire [7:0] t_r9_c55_3;
  wire [7:0] t_r9_c55_4;
  wire [7:0] t_r9_c55_5;
  wire [7:0] t_r9_c55_6;
  wire [7:0] t_r9_c55_7;
  wire [7:0] t_r9_c55_8;
  wire [7:0] t_r9_c55_9;
  wire [7:0] t_r9_c55_10;
  wire [7:0] t_r9_c55_11;
  wire [7:0] t_r9_c55_12;
  wire [7:0] t_r9_c56_0;
  wire [7:0] t_r9_c56_1;
  wire [7:0] t_r9_c56_2;
  wire [7:0] t_r9_c56_3;
  wire [7:0] t_r9_c56_4;
  wire [7:0] t_r9_c56_5;
  wire [7:0] t_r9_c56_6;
  wire [7:0] t_r9_c56_7;
  wire [7:0] t_r9_c56_8;
  wire [7:0] t_r9_c56_9;
  wire [7:0] t_r9_c56_10;
  wire [7:0] t_r9_c56_11;
  wire [7:0] t_r9_c56_12;
  wire [7:0] t_r9_c57_0;
  wire [7:0] t_r9_c57_1;
  wire [7:0] t_r9_c57_2;
  wire [7:0] t_r9_c57_3;
  wire [7:0] t_r9_c57_4;
  wire [7:0] t_r9_c57_5;
  wire [7:0] t_r9_c57_6;
  wire [7:0] t_r9_c57_7;
  wire [7:0] t_r9_c57_8;
  wire [7:0] t_r9_c57_9;
  wire [7:0] t_r9_c57_10;
  wire [7:0] t_r9_c57_11;
  wire [7:0] t_r9_c57_12;
  wire [7:0] t_r9_c58_0;
  wire [7:0] t_r9_c58_1;
  wire [7:0] t_r9_c58_2;
  wire [7:0] t_r9_c58_3;
  wire [7:0] t_r9_c58_4;
  wire [7:0] t_r9_c58_5;
  wire [7:0] t_r9_c58_6;
  wire [7:0] t_r9_c58_7;
  wire [7:0] t_r9_c58_8;
  wire [7:0] t_r9_c58_9;
  wire [7:0] t_r9_c58_10;
  wire [7:0] t_r9_c58_11;
  wire [7:0] t_r9_c58_12;
  wire [7:0] t_r9_c59_0;
  wire [7:0] t_r9_c59_1;
  wire [7:0] t_r9_c59_2;
  wire [7:0] t_r9_c59_3;
  wire [7:0] t_r9_c59_4;
  wire [7:0] t_r9_c59_5;
  wire [7:0] t_r9_c59_6;
  wire [7:0] t_r9_c59_7;
  wire [7:0] t_r9_c59_8;
  wire [7:0] t_r9_c59_9;
  wire [7:0] t_r9_c59_10;
  wire [7:0] t_r9_c59_11;
  wire [7:0] t_r9_c59_12;
  wire [7:0] t_r9_c60_0;
  wire [7:0] t_r9_c60_1;
  wire [7:0] t_r9_c60_2;
  wire [7:0] t_r9_c60_3;
  wire [7:0] t_r9_c60_4;
  wire [7:0] t_r9_c60_5;
  wire [7:0] t_r9_c60_6;
  wire [7:0] t_r9_c60_7;
  wire [7:0] t_r9_c60_8;
  wire [7:0] t_r9_c60_9;
  wire [7:0] t_r9_c60_10;
  wire [7:0] t_r9_c60_11;
  wire [7:0] t_r9_c60_12;
  wire [7:0] t_r9_c61_0;
  wire [7:0] t_r9_c61_1;
  wire [7:0] t_r9_c61_2;
  wire [7:0] t_r9_c61_3;
  wire [7:0] t_r9_c61_4;
  wire [7:0] t_r9_c61_5;
  wire [7:0] t_r9_c61_6;
  wire [7:0] t_r9_c61_7;
  wire [7:0] t_r9_c61_8;
  wire [7:0] t_r9_c61_9;
  wire [7:0] t_r9_c61_10;
  wire [7:0] t_r9_c61_11;
  wire [7:0] t_r9_c61_12;
  wire [7:0] t_r9_c62_0;
  wire [7:0] t_r9_c62_1;
  wire [7:0] t_r9_c62_2;
  wire [7:0] t_r9_c62_3;
  wire [7:0] t_r9_c62_4;
  wire [7:0] t_r9_c62_5;
  wire [7:0] t_r9_c62_6;
  wire [7:0] t_r9_c62_7;
  wire [7:0] t_r9_c62_8;
  wire [7:0] t_r9_c62_9;
  wire [7:0] t_r9_c62_10;
  wire [7:0] t_r9_c62_11;
  wire [7:0] t_r9_c62_12;
  wire [7:0] t_r9_c63_0;
  wire [7:0] t_r9_c63_1;
  wire [7:0] t_r9_c63_2;
  wire [7:0] t_r9_c63_3;
  wire [7:0] t_r9_c63_4;
  wire [7:0] t_r9_c63_5;
  wire [7:0] t_r9_c63_6;
  wire [7:0] t_r9_c63_7;
  wire [7:0] t_r9_c63_8;
  wire [7:0] t_r9_c63_9;
  wire [7:0] t_r9_c63_10;
  wire [7:0] t_r9_c63_11;
  wire [7:0] t_r9_c63_12;
  wire [7:0] t_r9_c64_0;
  wire [7:0] t_r9_c64_1;
  wire [7:0] t_r9_c64_2;
  wire [7:0] t_r9_c64_3;
  wire [7:0] t_r9_c64_4;
  wire [7:0] t_r9_c64_5;
  wire [7:0] t_r9_c64_6;
  wire [7:0] t_r9_c64_7;
  wire [7:0] t_r9_c64_8;
  wire [7:0] t_r9_c64_9;
  wire [7:0] t_r9_c64_10;
  wire [7:0] t_r9_c64_11;
  wire [7:0] t_r9_c64_12;
  wire [7:0] t_r9_c65_0;
  wire [7:0] t_r9_c65_1;
  wire [7:0] t_r9_c65_2;
  wire [7:0] t_r9_c65_3;
  wire [7:0] t_r9_c65_4;
  wire [7:0] t_r9_c65_5;
  wire [7:0] t_r9_c65_6;
  wire [7:0] t_r9_c65_7;
  wire [7:0] t_r9_c65_8;
  wire [7:0] t_r9_c65_9;
  wire [7:0] t_r9_c65_10;
  wire [7:0] t_r9_c65_11;
  wire [7:0] t_r9_c65_12;
  wire [7:0] t_r10_c0_0;
  wire [7:0] t_r10_c0_1;
  wire [7:0] t_r10_c0_2;
  wire [7:0] t_r10_c0_3;
  wire [7:0] t_r10_c0_4;
  wire [7:0] t_r10_c0_5;
  wire [7:0] t_r10_c0_6;
  wire [7:0] t_r10_c0_7;
  wire [7:0] t_r10_c0_8;
  wire [7:0] t_r10_c0_9;
  wire [7:0] t_r10_c0_10;
  wire [7:0] t_r10_c0_11;
  wire [7:0] t_r10_c0_12;
  wire [7:0] t_r10_c1_0;
  wire [7:0] t_r10_c1_1;
  wire [7:0] t_r10_c1_2;
  wire [7:0] t_r10_c1_3;
  wire [7:0] t_r10_c1_4;
  wire [7:0] t_r10_c1_5;
  wire [7:0] t_r10_c1_6;
  wire [7:0] t_r10_c1_7;
  wire [7:0] t_r10_c1_8;
  wire [7:0] t_r10_c1_9;
  wire [7:0] t_r10_c1_10;
  wire [7:0] t_r10_c1_11;
  wire [7:0] t_r10_c1_12;
  wire [7:0] t_r10_c2_0;
  wire [7:0] t_r10_c2_1;
  wire [7:0] t_r10_c2_2;
  wire [7:0] t_r10_c2_3;
  wire [7:0] t_r10_c2_4;
  wire [7:0] t_r10_c2_5;
  wire [7:0] t_r10_c2_6;
  wire [7:0] t_r10_c2_7;
  wire [7:0] t_r10_c2_8;
  wire [7:0] t_r10_c2_9;
  wire [7:0] t_r10_c2_10;
  wire [7:0] t_r10_c2_11;
  wire [7:0] t_r10_c2_12;
  wire [7:0] t_r10_c3_0;
  wire [7:0] t_r10_c3_1;
  wire [7:0] t_r10_c3_2;
  wire [7:0] t_r10_c3_3;
  wire [7:0] t_r10_c3_4;
  wire [7:0] t_r10_c3_5;
  wire [7:0] t_r10_c3_6;
  wire [7:0] t_r10_c3_7;
  wire [7:0] t_r10_c3_8;
  wire [7:0] t_r10_c3_9;
  wire [7:0] t_r10_c3_10;
  wire [7:0] t_r10_c3_11;
  wire [7:0] t_r10_c3_12;
  wire [7:0] t_r10_c4_0;
  wire [7:0] t_r10_c4_1;
  wire [7:0] t_r10_c4_2;
  wire [7:0] t_r10_c4_3;
  wire [7:0] t_r10_c4_4;
  wire [7:0] t_r10_c4_5;
  wire [7:0] t_r10_c4_6;
  wire [7:0] t_r10_c4_7;
  wire [7:0] t_r10_c4_8;
  wire [7:0] t_r10_c4_9;
  wire [7:0] t_r10_c4_10;
  wire [7:0] t_r10_c4_11;
  wire [7:0] t_r10_c4_12;
  wire [7:0] t_r10_c5_0;
  wire [7:0] t_r10_c5_1;
  wire [7:0] t_r10_c5_2;
  wire [7:0] t_r10_c5_3;
  wire [7:0] t_r10_c5_4;
  wire [7:0] t_r10_c5_5;
  wire [7:0] t_r10_c5_6;
  wire [7:0] t_r10_c5_7;
  wire [7:0] t_r10_c5_8;
  wire [7:0] t_r10_c5_9;
  wire [7:0] t_r10_c5_10;
  wire [7:0] t_r10_c5_11;
  wire [7:0] t_r10_c5_12;
  wire [7:0] t_r10_c6_0;
  wire [7:0] t_r10_c6_1;
  wire [7:0] t_r10_c6_2;
  wire [7:0] t_r10_c6_3;
  wire [7:0] t_r10_c6_4;
  wire [7:0] t_r10_c6_5;
  wire [7:0] t_r10_c6_6;
  wire [7:0] t_r10_c6_7;
  wire [7:0] t_r10_c6_8;
  wire [7:0] t_r10_c6_9;
  wire [7:0] t_r10_c6_10;
  wire [7:0] t_r10_c6_11;
  wire [7:0] t_r10_c6_12;
  wire [7:0] t_r10_c7_0;
  wire [7:0] t_r10_c7_1;
  wire [7:0] t_r10_c7_2;
  wire [7:0] t_r10_c7_3;
  wire [7:0] t_r10_c7_4;
  wire [7:0] t_r10_c7_5;
  wire [7:0] t_r10_c7_6;
  wire [7:0] t_r10_c7_7;
  wire [7:0] t_r10_c7_8;
  wire [7:0] t_r10_c7_9;
  wire [7:0] t_r10_c7_10;
  wire [7:0] t_r10_c7_11;
  wire [7:0] t_r10_c7_12;
  wire [7:0] t_r10_c8_0;
  wire [7:0] t_r10_c8_1;
  wire [7:0] t_r10_c8_2;
  wire [7:0] t_r10_c8_3;
  wire [7:0] t_r10_c8_4;
  wire [7:0] t_r10_c8_5;
  wire [7:0] t_r10_c8_6;
  wire [7:0] t_r10_c8_7;
  wire [7:0] t_r10_c8_8;
  wire [7:0] t_r10_c8_9;
  wire [7:0] t_r10_c8_10;
  wire [7:0] t_r10_c8_11;
  wire [7:0] t_r10_c8_12;
  wire [7:0] t_r10_c9_0;
  wire [7:0] t_r10_c9_1;
  wire [7:0] t_r10_c9_2;
  wire [7:0] t_r10_c9_3;
  wire [7:0] t_r10_c9_4;
  wire [7:0] t_r10_c9_5;
  wire [7:0] t_r10_c9_6;
  wire [7:0] t_r10_c9_7;
  wire [7:0] t_r10_c9_8;
  wire [7:0] t_r10_c9_9;
  wire [7:0] t_r10_c9_10;
  wire [7:0] t_r10_c9_11;
  wire [7:0] t_r10_c9_12;
  wire [7:0] t_r10_c10_0;
  wire [7:0] t_r10_c10_1;
  wire [7:0] t_r10_c10_2;
  wire [7:0] t_r10_c10_3;
  wire [7:0] t_r10_c10_4;
  wire [7:0] t_r10_c10_5;
  wire [7:0] t_r10_c10_6;
  wire [7:0] t_r10_c10_7;
  wire [7:0] t_r10_c10_8;
  wire [7:0] t_r10_c10_9;
  wire [7:0] t_r10_c10_10;
  wire [7:0] t_r10_c10_11;
  wire [7:0] t_r10_c10_12;
  wire [7:0] t_r10_c11_0;
  wire [7:0] t_r10_c11_1;
  wire [7:0] t_r10_c11_2;
  wire [7:0] t_r10_c11_3;
  wire [7:0] t_r10_c11_4;
  wire [7:0] t_r10_c11_5;
  wire [7:0] t_r10_c11_6;
  wire [7:0] t_r10_c11_7;
  wire [7:0] t_r10_c11_8;
  wire [7:0] t_r10_c11_9;
  wire [7:0] t_r10_c11_10;
  wire [7:0] t_r10_c11_11;
  wire [7:0] t_r10_c11_12;
  wire [7:0] t_r10_c12_0;
  wire [7:0] t_r10_c12_1;
  wire [7:0] t_r10_c12_2;
  wire [7:0] t_r10_c12_3;
  wire [7:0] t_r10_c12_4;
  wire [7:0] t_r10_c12_5;
  wire [7:0] t_r10_c12_6;
  wire [7:0] t_r10_c12_7;
  wire [7:0] t_r10_c12_8;
  wire [7:0] t_r10_c12_9;
  wire [7:0] t_r10_c12_10;
  wire [7:0] t_r10_c12_11;
  wire [7:0] t_r10_c12_12;
  wire [7:0] t_r10_c13_0;
  wire [7:0] t_r10_c13_1;
  wire [7:0] t_r10_c13_2;
  wire [7:0] t_r10_c13_3;
  wire [7:0] t_r10_c13_4;
  wire [7:0] t_r10_c13_5;
  wire [7:0] t_r10_c13_6;
  wire [7:0] t_r10_c13_7;
  wire [7:0] t_r10_c13_8;
  wire [7:0] t_r10_c13_9;
  wire [7:0] t_r10_c13_10;
  wire [7:0] t_r10_c13_11;
  wire [7:0] t_r10_c13_12;
  wire [7:0] t_r10_c14_0;
  wire [7:0] t_r10_c14_1;
  wire [7:0] t_r10_c14_2;
  wire [7:0] t_r10_c14_3;
  wire [7:0] t_r10_c14_4;
  wire [7:0] t_r10_c14_5;
  wire [7:0] t_r10_c14_6;
  wire [7:0] t_r10_c14_7;
  wire [7:0] t_r10_c14_8;
  wire [7:0] t_r10_c14_9;
  wire [7:0] t_r10_c14_10;
  wire [7:0] t_r10_c14_11;
  wire [7:0] t_r10_c14_12;
  wire [7:0] t_r10_c15_0;
  wire [7:0] t_r10_c15_1;
  wire [7:0] t_r10_c15_2;
  wire [7:0] t_r10_c15_3;
  wire [7:0] t_r10_c15_4;
  wire [7:0] t_r10_c15_5;
  wire [7:0] t_r10_c15_6;
  wire [7:0] t_r10_c15_7;
  wire [7:0] t_r10_c15_8;
  wire [7:0] t_r10_c15_9;
  wire [7:0] t_r10_c15_10;
  wire [7:0] t_r10_c15_11;
  wire [7:0] t_r10_c15_12;
  wire [7:0] t_r10_c16_0;
  wire [7:0] t_r10_c16_1;
  wire [7:0] t_r10_c16_2;
  wire [7:0] t_r10_c16_3;
  wire [7:0] t_r10_c16_4;
  wire [7:0] t_r10_c16_5;
  wire [7:0] t_r10_c16_6;
  wire [7:0] t_r10_c16_7;
  wire [7:0] t_r10_c16_8;
  wire [7:0] t_r10_c16_9;
  wire [7:0] t_r10_c16_10;
  wire [7:0] t_r10_c16_11;
  wire [7:0] t_r10_c16_12;
  wire [7:0] t_r10_c17_0;
  wire [7:0] t_r10_c17_1;
  wire [7:0] t_r10_c17_2;
  wire [7:0] t_r10_c17_3;
  wire [7:0] t_r10_c17_4;
  wire [7:0] t_r10_c17_5;
  wire [7:0] t_r10_c17_6;
  wire [7:0] t_r10_c17_7;
  wire [7:0] t_r10_c17_8;
  wire [7:0] t_r10_c17_9;
  wire [7:0] t_r10_c17_10;
  wire [7:0] t_r10_c17_11;
  wire [7:0] t_r10_c17_12;
  wire [7:0] t_r10_c18_0;
  wire [7:0] t_r10_c18_1;
  wire [7:0] t_r10_c18_2;
  wire [7:0] t_r10_c18_3;
  wire [7:0] t_r10_c18_4;
  wire [7:0] t_r10_c18_5;
  wire [7:0] t_r10_c18_6;
  wire [7:0] t_r10_c18_7;
  wire [7:0] t_r10_c18_8;
  wire [7:0] t_r10_c18_9;
  wire [7:0] t_r10_c18_10;
  wire [7:0] t_r10_c18_11;
  wire [7:0] t_r10_c18_12;
  wire [7:0] t_r10_c19_0;
  wire [7:0] t_r10_c19_1;
  wire [7:0] t_r10_c19_2;
  wire [7:0] t_r10_c19_3;
  wire [7:0] t_r10_c19_4;
  wire [7:0] t_r10_c19_5;
  wire [7:0] t_r10_c19_6;
  wire [7:0] t_r10_c19_7;
  wire [7:0] t_r10_c19_8;
  wire [7:0] t_r10_c19_9;
  wire [7:0] t_r10_c19_10;
  wire [7:0] t_r10_c19_11;
  wire [7:0] t_r10_c19_12;
  wire [7:0] t_r10_c20_0;
  wire [7:0] t_r10_c20_1;
  wire [7:0] t_r10_c20_2;
  wire [7:0] t_r10_c20_3;
  wire [7:0] t_r10_c20_4;
  wire [7:0] t_r10_c20_5;
  wire [7:0] t_r10_c20_6;
  wire [7:0] t_r10_c20_7;
  wire [7:0] t_r10_c20_8;
  wire [7:0] t_r10_c20_9;
  wire [7:0] t_r10_c20_10;
  wire [7:0] t_r10_c20_11;
  wire [7:0] t_r10_c20_12;
  wire [7:0] t_r10_c21_0;
  wire [7:0] t_r10_c21_1;
  wire [7:0] t_r10_c21_2;
  wire [7:0] t_r10_c21_3;
  wire [7:0] t_r10_c21_4;
  wire [7:0] t_r10_c21_5;
  wire [7:0] t_r10_c21_6;
  wire [7:0] t_r10_c21_7;
  wire [7:0] t_r10_c21_8;
  wire [7:0] t_r10_c21_9;
  wire [7:0] t_r10_c21_10;
  wire [7:0] t_r10_c21_11;
  wire [7:0] t_r10_c21_12;
  wire [7:0] t_r10_c22_0;
  wire [7:0] t_r10_c22_1;
  wire [7:0] t_r10_c22_2;
  wire [7:0] t_r10_c22_3;
  wire [7:0] t_r10_c22_4;
  wire [7:0] t_r10_c22_5;
  wire [7:0] t_r10_c22_6;
  wire [7:0] t_r10_c22_7;
  wire [7:0] t_r10_c22_8;
  wire [7:0] t_r10_c22_9;
  wire [7:0] t_r10_c22_10;
  wire [7:0] t_r10_c22_11;
  wire [7:0] t_r10_c22_12;
  wire [7:0] t_r10_c23_0;
  wire [7:0] t_r10_c23_1;
  wire [7:0] t_r10_c23_2;
  wire [7:0] t_r10_c23_3;
  wire [7:0] t_r10_c23_4;
  wire [7:0] t_r10_c23_5;
  wire [7:0] t_r10_c23_6;
  wire [7:0] t_r10_c23_7;
  wire [7:0] t_r10_c23_8;
  wire [7:0] t_r10_c23_9;
  wire [7:0] t_r10_c23_10;
  wire [7:0] t_r10_c23_11;
  wire [7:0] t_r10_c23_12;
  wire [7:0] t_r10_c24_0;
  wire [7:0] t_r10_c24_1;
  wire [7:0] t_r10_c24_2;
  wire [7:0] t_r10_c24_3;
  wire [7:0] t_r10_c24_4;
  wire [7:0] t_r10_c24_5;
  wire [7:0] t_r10_c24_6;
  wire [7:0] t_r10_c24_7;
  wire [7:0] t_r10_c24_8;
  wire [7:0] t_r10_c24_9;
  wire [7:0] t_r10_c24_10;
  wire [7:0] t_r10_c24_11;
  wire [7:0] t_r10_c24_12;
  wire [7:0] t_r10_c25_0;
  wire [7:0] t_r10_c25_1;
  wire [7:0] t_r10_c25_2;
  wire [7:0] t_r10_c25_3;
  wire [7:0] t_r10_c25_4;
  wire [7:0] t_r10_c25_5;
  wire [7:0] t_r10_c25_6;
  wire [7:0] t_r10_c25_7;
  wire [7:0] t_r10_c25_8;
  wire [7:0] t_r10_c25_9;
  wire [7:0] t_r10_c25_10;
  wire [7:0] t_r10_c25_11;
  wire [7:0] t_r10_c25_12;
  wire [7:0] t_r10_c26_0;
  wire [7:0] t_r10_c26_1;
  wire [7:0] t_r10_c26_2;
  wire [7:0] t_r10_c26_3;
  wire [7:0] t_r10_c26_4;
  wire [7:0] t_r10_c26_5;
  wire [7:0] t_r10_c26_6;
  wire [7:0] t_r10_c26_7;
  wire [7:0] t_r10_c26_8;
  wire [7:0] t_r10_c26_9;
  wire [7:0] t_r10_c26_10;
  wire [7:0] t_r10_c26_11;
  wire [7:0] t_r10_c26_12;
  wire [7:0] t_r10_c27_0;
  wire [7:0] t_r10_c27_1;
  wire [7:0] t_r10_c27_2;
  wire [7:0] t_r10_c27_3;
  wire [7:0] t_r10_c27_4;
  wire [7:0] t_r10_c27_5;
  wire [7:0] t_r10_c27_6;
  wire [7:0] t_r10_c27_7;
  wire [7:0] t_r10_c27_8;
  wire [7:0] t_r10_c27_9;
  wire [7:0] t_r10_c27_10;
  wire [7:0] t_r10_c27_11;
  wire [7:0] t_r10_c27_12;
  wire [7:0] t_r10_c28_0;
  wire [7:0] t_r10_c28_1;
  wire [7:0] t_r10_c28_2;
  wire [7:0] t_r10_c28_3;
  wire [7:0] t_r10_c28_4;
  wire [7:0] t_r10_c28_5;
  wire [7:0] t_r10_c28_6;
  wire [7:0] t_r10_c28_7;
  wire [7:0] t_r10_c28_8;
  wire [7:0] t_r10_c28_9;
  wire [7:0] t_r10_c28_10;
  wire [7:0] t_r10_c28_11;
  wire [7:0] t_r10_c28_12;
  wire [7:0] t_r10_c29_0;
  wire [7:0] t_r10_c29_1;
  wire [7:0] t_r10_c29_2;
  wire [7:0] t_r10_c29_3;
  wire [7:0] t_r10_c29_4;
  wire [7:0] t_r10_c29_5;
  wire [7:0] t_r10_c29_6;
  wire [7:0] t_r10_c29_7;
  wire [7:0] t_r10_c29_8;
  wire [7:0] t_r10_c29_9;
  wire [7:0] t_r10_c29_10;
  wire [7:0] t_r10_c29_11;
  wire [7:0] t_r10_c29_12;
  wire [7:0] t_r10_c30_0;
  wire [7:0] t_r10_c30_1;
  wire [7:0] t_r10_c30_2;
  wire [7:0] t_r10_c30_3;
  wire [7:0] t_r10_c30_4;
  wire [7:0] t_r10_c30_5;
  wire [7:0] t_r10_c30_6;
  wire [7:0] t_r10_c30_7;
  wire [7:0] t_r10_c30_8;
  wire [7:0] t_r10_c30_9;
  wire [7:0] t_r10_c30_10;
  wire [7:0] t_r10_c30_11;
  wire [7:0] t_r10_c30_12;
  wire [7:0] t_r10_c31_0;
  wire [7:0] t_r10_c31_1;
  wire [7:0] t_r10_c31_2;
  wire [7:0] t_r10_c31_3;
  wire [7:0] t_r10_c31_4;
  wire [7:0] t_r10_c31_5;
  wire [7:0] t_r10_c31_6;
  wire [7:0] t_r10_c31_7;
  wire [7:0] t_r10_c31_8;
  wire [7:0] t_r10_c31_9;
  wire [7:0] t_r10_c31_10;
  wire [7:0] t_r10_c31_11;
  wire [7:0] t_r10_c31_12;
  wire [7:0] t_r10_c32_0;
  wire [7:0] t_r10_c32_1;
  wire [7:0] t_r10_c32_2;
  wire [7:0] t_r10_c32_3;
  wire [7:0] t_r10_c32_4;
  wire [7:0] t_r10_c32_5;
  wire [7:0] t_r10_c32_6;
  wire [7:0] t_r10_c32_7;
  wire [7:0] t_r10_c32_8;
  wire [7:0] t_r10_c32_9;
  wire [7:0] t_r10_c32_10;
  wire [7:0] t_r10_c32_11;
  wire [7:0] t_r10_c32_12;
  wire [7:0] t_r10_c33_0;
  wire [7:0] t_r10_c33_1;
  wire [7:0] t_r10_c33_2;
  wire [7:0] t_r10_c33_3;
  wire [7:0] t_r10_c33_4;
  wire [7:0] t_r10_c33_5;
  wire [7:0] t_r10_c33_6;
  wire [7:0] t_r10_c33_7;
  wire [7:0] t_r10_c33_8;
  wire [7:0] t_r10_c33_9;
  wire [7:0] t_r10_c33_10;
  wire [7:0] t_r10_c33_11;
  wire [7:0] t_r10_c33_12;
  wire [7:0] t_r10_c34_0;
  wire [7:0] t_r10_c34_1;
  wire [7:0] t_r10_c34_2;
  wire [7:0] t_r10_c34_3;
  wire [7:0] t_r10_c34_4;
  wire [7:0] t_r10_c34_5;
  wire [7:0] t_r10_c34_6;
  wire [7:0] t_r10_c34_7;
  wire [7:0] t_r10_c34_8;
  wire [7:0] t_r10_c34_9;
  wire [7:0] t_r10_c34_10;
  wire [7:0] t_r10_c34_11;
  wire [7:0] t_r10_c34_12;
  wire [7:0] t_r10_c35_0;
  wire [7:0] t_r10_c35_1;
  wire [7:0] t_r10_c35_2;
  wire [7:0] t_r10_c35_3;
  wire [7:0] t_r10_c35_4;
  wire [7:0] t_r10_c35_5;
  wire [7:0] t_r10_c35_6;
  wire [7:0] t_r10_c35_7;
  wire [7:0] t_r10_c35_8;
  wire [7:0] t_r10_c35_9;
  wire [7:0] t_r10_c35_10;
  wire [7:0] t_r10_c35_11;
  wire [7:0] t_r10_c35_12;
  wire [7:0] t_r10_c36_0;
  wire [7:0] t_r10_c36_1;
  wire [7:0] t_r10_c36_2;
  wire [7:0] t_r10_c36_3;
  wire [7:0] t_r10_c36_4;
  wire [7:0] t_r10_c36_5;
  wire [7:0] t_r10_c36_6;
  wire [7:0] t_r10_c36_7;
  wire [7:0] t_r10_c36_8;
  wire [7:0] t_r10_c36_9;
  wire [7:0] t_r10_c36_10;
  wire [7:0] t_r10_c36_11;
  wire [7:0] t_r10_c36_12;
  wire [7:0] t_r10_c37_0;
  wire [7:0] t_r10_c37_1;
  wire [7:0] t_r10_c37_2;
  wire [7:0] t_r10_c37_3;
  wire [7:0] t_r10_c37_4;
  wire [7:0] t_r10_c37_5;
  wire [7:0] t_r10_c37_6;
  wire [7:0] t_r10_c37_7;
  wire [7:0] t_r10_c37_8;
  wire [7:0] t_r10_c37_9;
  wire [7:0] t_r10_c37_10;
  wire [7:0] t_r10_c37_11;
  wire [7:0] t_r10_c37_12;
  wire [7:0] t_r10_c38_0;
  wire [7:0] t_r10_c38_1;
  wire [7:0] t_r10_c38_2;
  wire [7:0] t_r10_c38_3;
  wire [7:0] t_r10_c38_4;
  wire [7:0] t_r10_c38_5;
  wire [7:0] t_r10_c38_6;
  wire [7:0] t_r10_c38_7;
  wire [7:0] t_r10_c38_8;
  wire [7:0] t_r10_c38_9;
  wire [7:0] t_r10_c38_10;
  wire [7:0] t_r10_c38_11;
  wire [7:0] t_r10_c38_12;
  wire [7:0] t_r10_c39_0;
  wire [7:0] t_r10_c39_1;
  wire [7:0] t_r10_c39_2;
  wire [7:0] t_r10_c39_3;
  wire [7:0] t_r10_c39_4;
  wire [7:0] t_r10_c39_5;
  wire [7:0] t_r10_c39_6;
  wire [7:0] t_r10_c39_7;
  wire [7:0] t_r10_c39_8;
  wire [7:0] t_r10_c39_9;
  wire [7:0] t_r10_c39_10;
  wire [7:0] t_r10_c39_11;
  wire [7:0] t_r10_c39_12;
  wire [7:0] t_r10_c40_0;
  wire [7:0] t_r10_c40_1;
  wire [7:0] t_r10_c40_2;
  wire [7:0] t_r10_c40_3;
  wire [7:0] t_r10_c40_4;
  wire [7:0] t_r10_c40_5;
  wire [7:0] t_r10_c40_6;
  wire [7:0] t_r10_c40_7;
  wire [7:0] t_r10_c40_8;
  wire [7:0] t_r10_c40_9;
  wire [7:0] t_r10_c40_10;
  wire [7:0] t_r10_c40_11;
  wire [7:0] t_r10_c40_12;
  wire [7:0] t_r10_c41_0;
  wire [7:0] t_r10_c41_1;
  wire [7:0] t_r10_c41_2;
  wire [7:0] t_r10_c41_3;
  wire [7:0] t_r10_c41_4;
  wire [7:0] t_r10_c41_5;
  wire [7:0] t_r10_c41_6;
  wire [7:0] t_r10_c41_7;
  wire [7:0] t_r10_c41_8;
  wire [7:0] t_r10_c41_9;
  wire [7:0] t_r10_c41_10;
  wire [7:0] t_r10_c41_11;
  wire [7:0] t_r10_c41_12;
  wire [7:0] t_r10_c42_0;
  wire [7:0] t_r10_c42_1;
  wire [7:0] t_r10_c42_2;
  wire [7:0] t_r10_c42_3;
  wire [7:0] t_r10_c42_4;
  wire [7:0] t_r10_c42_5;
  wire [7:0] t_r10_c42_6;
  wire [7:0] t_r10_c42_7;
  wire [7:0] t_r10_c42_8;
  wire [7:0] t_r10_c42_9;
  wire [7:0] t_r10_c42_10;
  wire [7:0] t_r10_c42_11;
  wire [7:0] t_r10_c42_12;
  wire [7:0] t_r10_c43_0;
  wire [7:0] t_r10_c43_1;
  wire [7:0] t_r10_c43_2;
  wire [7:0] t_r10_c43_3;
  wire [7:0] t_r10_c43_4;
  wire [7:0] t_r10_c43_5;
  wire [7:0] t_r10_c43_6;
  wire [7:0] t_r10_c43_7;
  wire [7:0] t_r10_c43_8;
  wire [7:0] t_r10_c43_9;
  wire [7:0] t_r10_c43_10;
  wire [7:0] t_r10_c43_11;
  wire [7:0] t_r10_c43_12;
  wire [7:0] t_r10_c44_0;
  wire [7:0] t_r10_c44_1;
  wire [7:0] t_r10_c44_2;
  wire [7:0] t_r10_c44_3;
  wire [7:0] t_r10_c44_4;
  wire [7:0] t_r10_c44_5;
  wire [7:0] t_r10_c44_6;
  wire [7:0] t_r10_c44_7;
  wire [7:0] t_r10_c44_8;
  wire [7:0] t_r10_c44_9;
  wire [7:0] t_r10_c44_10;
  wire [7:0] t_r10_c44_11;
  wire [7:0] t_r10_c44_12;
  wire [7:0] t_r10_c45_0;
  wire [7:0] t_r10_c45_1;
  wire [7:0] t_r10_c45_2;
  wire [7:0] t_r10_c45_3;
  wire [7:0] t_r10_c45_4;
  wire [7:0] t_r10_c45_5;
  wire [7:0] t_r10_c45_6;
  wire [7:0] t_r10_c45_7;
  wire [7:0] t_r10_c45_8;
  wire [7:0] t_r10_c45_9;
  wire [7:0] t_r10_c45_10;
  wire [7:0] t_r10_c45_11;
  wire [7:0] t_r10_c45_12;
  wire [7:0] t_r10_c46_0;
  wire [7:0] t_r10_c46_1;
  wire [7:0] t_r10_c46_2;
  wire [7:0] t_r10_c46_3;
  wire [7:0] t_r10_c46_4;
  wire [7:0] t_r10_c46_5;
  wire [7:0] t_r10_c46_6;
  wire [7:0] t_r10_c46_7;
  wire [7:0] t_r10_c46_8;
  wire [7:0] t_r10_c46_9;
  wire [7:0] t_r10_c46_10;
  wire [7:0] t_r10_c46_11;
  wire [7:0] t_r10_c46_12;
  wire [7:0] t_r10_c47_0;
  wire [7:0] t_r10_c47_1;
  wire [7:0] t_r10_c47_2;
  wire [7:0] t_r10_c47_3;
  wire [7:0] t_r10_c47_4;
  wire [7:0] t_r10_c47_5;
  wire [7:0] t_r10_c47_6;
  wire [7:0] t_r10_c47_7;
  wire [7:0] t_r10_c47_8;
  wire [7:0] t_r10_c47_9;
  wire [7:0] t_r10_c47_10;
  wire [7:0] t_r10_c47_11;
  wire [7:0] t_r10_c47_12;
  wire [7:0] t_r10_c48_0;
  wire [7:0] t_r10_c48_1;
  wire [7:0] t_r10_c48_2;
  wire [7:0] t_r10_c48_3;
  wire [7:0] t_r10_c48_4;
  wire [7:0] t_r10_c48_5;
  wire [7:0] t_r10_c48_6;
  wire [7:0] t_r10_c48_7;
  wire [7:0] t_r10_c48_8;
  wire [7:0] t_r10_c48_9;
  wire [7:0] t_r10_c48_10;
  wire [7:0] t_r10_c48_11;
  wire [7:0] t_r10_c48_12;
  wire [7:0] t_r10_c49_0;
  wire [7:0] t_r10_c49_1;
  wire [7:0] t_r10_c49_2;
  wire [7:0] t_r10_c49_3;
  wire [7:0] t_r10_c49_4;
  wire [7:0] t_r10_c49_5;
  wire [7:0] t_r10_c49_6;
  wire [7:0] t_r10_c49_7;
  wire [7:0] t_r10_c49_8;
  wire [7:0] t_r10_c49_9;
  wire [7:0] t_r10_c49_10;
  wire [7:0] t_r10_c49_11;
  wire [7:0] t_r10_c49_12;
  wire [7:0] t_r10_c50_0;
  wire [7:0] t_r10_c50_1;
  wire [7:0] t_r10_c50_2;
  wire [7:0] t_r10_c50_3;
  wire [7:0] t_r10_c50_4;
  wire [7:0] t_r10_c50_5;
  wire [7:0] t_r10_c50_6;
  wire [7:0] t_r10_c50_7;
  wire [7:0] t_r10_c50_8;
  wire [7:0] t_r10_c50_9;
  wire [7:0] t_r10_c50_10;
  wire [7:0] t_r10_c50_11;
  wire [7:0] t_r10_c50_12;
  wire [7:0] t_r10_c51_0;
  wire [7:0] t_r10_c51_1;
  wire [7:0] t_r10_c51_2;
  wire [7:0] t_r10_c51_3;
  wire [7:0] t_r10_c51_4;
  wire [7:0] t_r10_c51_5;
  wire [7:0] t_r10_c51_6;
  wire [7:0] t_r10_c51_7;
  wire [7:0] t_r10_c51_8;
  wire [7:0] t_r10_c51_9;
  wire [7:0] t_r10_c51_10;
  wire [7:0] t_r10_c51_11;
  wire [7:0] t_r10_c51_12;
  wire [7:0] t_r10_c52_0;
  wire [7:0] t_r10_c52_1;
  wire [7:0] t_r10_c52_2;
  wire [7:0] t_r10_c52_3;
  wire [7:0] t_r10_c52_4;
  wire [7:0] t_r10_c52_5;
  wire [7:0] t_r10_c52_6;
  wire [7:0] t_r10_c52_7;
  wire [7:0] t_r10_c52_8;
  wire [7:0] t_r10_c52_9;
  wire [7:0] t_r10_c52_10;
  wire [7:0] t_r10_c52_11;
  wire [7:0] t_r10_c52_12;
  wire [7:0] t_r10_c53_0;
  wire [7:0] t_r10_c53_1;
  wire [7:0] t_r10_c53_2;
  wire [7:0] t_r10_c53_3;
  wire [7:0] t_r10_c53_4;
  wire [7:0] t_r10_c53_5;
  wire [7:0] t_r10_c53_6;
  wire [7:0] t_r10_c53_7;
  wire [7:0] t_r10_c53_8;
  wire [7:0] t_r10_c53_9;
  wire [7:0] t_r10_c53_10;
  wire [7:0] t_r10_c53_11;
  wire [7:0] t_r10_c53_12;
  wire [7:0] t_r10_c54_0;
  wire [7:0] t_r10_c54_1;
  wire [7:0] t_r10_c54_2;
  wire [7:0] t_r10_c54_3;
  wire [7:0] t_r10_c54_4;
  wire [7:0] t_r10_c54_5;
  wire [7:0] t_r10_c54_6;
  wire [7:0] t_r10_c54_7;
  wire [7:0] t_r10_c54_8;
  wire [7:0] t_r10_c54_9;
  wire [7:0] t_r10_c54_10;
  wire [7:0] t_r10_c54_11;
  wire [7:0] t_r10_c54_12;
  wire [7:0] t_r10_c55_0;
  wire [7:0] t_r10_c55_1;
  wire [7:0] t_r10_c55_2;
  wire [7:0] t_r10_c55_3;
  wire [7:0] t_r10_c55_4;
  wire [7:0] t_r10_c55_5;
  wire [7:0] t_r10_c55_6;
  wire [7:0] t_r10_c55_7;
  wire [7:0] t_r10_c55_8;
  wire [7:0] t_r10_c55_9;
  wire [7:0] t_r10_c55_10;
  wire [7:0] t_r10_c55_11;
  wire [7:0] t_r10_c55_12;
  wire [7:0] t_r10_c56_0;
  wire [7:0] t_r10_c56_1;
  wire [7:0] t_r10_c56_2;
  wire [7:0] t_r10_c56_3;
  wire [7:0] t_r10_c56_4;
  wire [7:0] t_r10_c56_5;
  wire [7:0] t_r10_c56_6;
  wire [7:0] t_r10_c56_7;
  wire [7:0] t_r10_c56_8;
  wire [7:0] t_r10_c56_9;
  wire [7:0] t_r10_c56_10;
  wire [7:0] t_r10_c56_11;
  wire [7:0] t_r10_c56_12;
  wire [7:0] t_r10_c57_0;
  wire [7:0] t_r10_c57_1;
  wire [7:0] t_r10_c57_2;
  wire [7:0] t_r10_c57_3;
  wire [7:0] t_r10_c57_4;
  wire [7:0] t_r10_c57_5;
  wire [7:0] t_r10_c57_6;
  wire [7:0] t_r10_c57_7;
  wire [7:0] t_r10_c57_8;
  wire [7:0] t_r10_c57_9;
  wire [7:0] t_r10_c57_10;
  wire [7:0] t_r10_c57_11;
  wire [7:0] t_r10_c57_12;
  wire [7:0] t_r10_c58_0;
  wire [7:0] t_r10_c58_1;
  wire [7:0] t_r10_c58_2;
  wire [7:0] t_r10_c58_3;
  wire [7:0] t_r10_c58_4;
  wire [7:0] t_r10_c58_5;
  wire [7:0] t_r10_c58_6;
  wire [7:0] t_r10_c58_7;
  wire [7:0] t_r10_c58_8;
  wire [7:0] t_r10_c58_9;
  wire [7:0] t_r10_c58_10;
  wire [7:0] t_r10_c58_11;
  wire [7:0] t_r10_c58_12;
  wire [7:0] t_r10_c59_0;
  wire [7:0] t_r10_c59_1;
  wire [7:0] t_r10_c59_2;
  wire [7:0] t_r10_c59_3;
  wire [7:0] t_r10_c59_4;
  wire [7:0] t_r10_c59_5;
  wire [7:0] t_r10_c59_6;
  wire [7:0] t_r10_c59_7;
  wire [7:0] t_r10_c59_8;
  wire [7:0] t_r10_c59_9;
  wire [7:0] t_r10_c59_10;
  wire [7:0] t_r10_c59_11;
  wire [7:0] t_r10_c59_12;
  wire [7:0] t_r10_c60_0;
  wire [7:0] t_r10_c60_1;
  wire [7:0] t_r10_c60_2;
  wire [7:0] t_r10_c60_3;
  wire [7:0] t_r10_c60_4;
  wire [7:0] t_r10_c60_5;
  wire [7:0] t_r10_c60_6;
  wire [7:0] t_r10_c60_7;
  wire [7:0] t_r10_c60_8;
  wire [7:0] t_r10_c60_9;
  wire [7:0] t_r10_c60_10;
  wire [7:0] t_r10_c60_11;
  wire [7:0] t_r10_c60_12;
  wire [7:0] t_r10_c61_0;
  wire [7:0] t_r10_c61_1;
  wire [7:0] t_r10_c61_2;
  wire [7:0] t_r10_c61_3;
  wire [7:0] t_r10_c61_4;
  wire [7:0] t_r10_c61_5;
  wire [7:0] t_r10_c61_6;
  wire [7:0] t_r10_c61_7;
  wire [7:0] t_r10_c61_8;
  wire [7:0] t_r10_c61_9;
  wire [7:0] t_r10_c61_10;
  wire [7:0] t_r10_c61_11;
  wire [7:0] t_r10_c61_12;
  wire [7:0] t_r10_c62_0;
  wire [7:0] t_r10_c62_1;
  wire [7:0] t_r10_c62_2;
  wire [7:0] t_r10_c62_3;
  wire [7:0] t_r10_c62_4;
  wire [7:0] t_r10_c62_5;
  wire [7:0] t_r10_c62_6;
  wire [7:0] t_r10_c62_7;
  wire [7:0] t_r10_c62_8;
  wire [7:0] t_r10_c62_9;
  wire [7:0] t_r10_c62_10;
  wire [7:0] t_r10_c62_11;
  wire [7:0] t_r10_c62_12;
  wire [7:0] t_r10_c63_0;
  wire [7:0] t_r10_c63_1;
  wire [7:0] t_r10_c63_2;
  wire [7:0] t_r10_c63_3;
  wire [7:0] t_r10_c63_4;
  wire [7:0] t_r10_c63_5;
  wire [7:0] t_r10_c63_6;
  wire [7:0] t_r10_c63_7;
  wire [7:0] t_r10_c63_8;
  wire [7:0] t_r10_c63_9;
  wire [7:0] t_r10_c63_10;
  wire [7:0] t_r10_c63_11;
  wire [7:0] t_r10_c63_12;
  wire [7:0] t_r10_c64_0;
  wire [7:0] t_r10_c64_1;
  wire [7:0] t_r10_c64_2;
  wire [7:0] t_r10_c64_3;
  wire [7:0] t_r10_c64_4;
  wire [7:0] t_r10_c64_5;
  wire [7:0] t_r10_c64_6;
  wire [7:0] t_r10_c64_7;
  wire [7:0] t_r10_c64_8;
  wire [7:0] t_r10_c64_9;
  wire [7:0] t_r10_c64_10;
  wire [7:0] t_r10_c64_11;
  wire [7:0] t_r10_c64_12;
  wire [7:0] t_r10_c65_0;
  wire [7:0] t_r10_c65_1;
  wire [7:0] t_r10_c65_2;
  wire [7:0] t_r10_c65_3;
  wire [7:0] t_r10_c65_4;
  wire [7:0] t_r10_c65_5;
  wire [7:0] t_r10_c65_6;
  wire [7:0] t_r10_c65_7;
  wire [7:0] t_r10_c65_8;
  wire [7:0] t_r10_c65_9;
  wire [7:0] t_r10_c65_10;
  wire [7:0] t_r10_c65_11;
  wire [7:0] t_r10_c65_12;
  wire [7:0] t_r11_c0_0;
  wire [7:0] t_r11_c0_1;
  wire [7:0] t_r11_c0_2;
  wire [7:0] t_r11_c0_3;
  wire [7:0] t_r11_c0_4;
  wire [7:0] t_r11_c0_5;
  wire [7:0] t_r11_c0_6;
  wire [7:0] t_r11_c0_7;
  wire [7:0] t_r11_c0_8;
  wire [7:0] t_r11_c0_9;
  wire [7:0] t_r11_c0_10;
  wire [7:0] t_r11_c0_11;
  wire [7:0] t_r11_c0_12;
  wire [7:0] t_r11_c1_0;
  wire [7:0] t_r11_c1_1;
  wire [7:0] t_r11_c1_2;
  wire [7:0] t_r11_c1_3;
  wire [7:0] t_r11_c1_4;
  wire [7:0] t_r11_c1_5;
  wire [7:0] t_r11_c1_6;
  wire [7:0] t_r11_c1_7;
  wire [7:0] t_r11_c1_8;
  wire [7:0] t_r11_c1_9;
  wire [7:0] t_r11_c1_10;
  wire [7:0] t_r11_c1_11;
  wire [7:0] t_r11_c1_12;
  wire [7:0] t_r11_c2_0;
  wire [7:0] t_r11_c2_1;
  wire [7:0] t_r11_c2_2;
  wire [7:0] t_r11_c2_3;
  wire [7:0] t_r11_c2_4;
  wire [7:0] t_r11_c2_5;
  wire [7:0] t_r11_c2_6;
  wire [7:0] t_r11_c2_7;
  wire [7:0] t_r11_c2_8;
  wire [7:0] t_r11_c2_9;
  wire [7:0] t_r11_c2_10;
  wire [7:0] t_r11_c2_11;
  wire [7:0] t_r11_c2_12;
  wire [7:0] t_r11_c3_0;
  wire [7:0] t_r11_c3_1;
  wire [7:0] t_r11_c3_2;
  wire [7:0] t_r11_c3_3;
  wire [7:0] t_r11_c3_4;
  wire [7:0] t_r11_c3_5;
  wire [7:0] t_r11_c3_6;
  wire [7:0] t_r11_c3_7;
  wire [7:0] t_r11_c3_8;
  wire [7:0] t_r11_c3_9;
  wire [7:0] t_r11_c3_10;
  wire [7:0] t_r11_c3_11;
  wire [7:0] t_r11_c3_12;
  wire [7:0] t_r11_c4_0;
  wire [7:0] t_r11_c4_1;
  wire [7:0] t_r11_c4_2;
  wire [7:0] t_r11_c4_3;
  wire [7:0] t_r11_c4_4;
  wire [7:0] t_r11_c4_5;
  wire [7:0] t_r11_c4_6;
  wire [7:0] t_r11_c4_7;
  wire [7:0] t_r11_c4_8;
  wire [7:0] t_r11_c4_9;
  wire [7:0] t_r11_c4_10;
  wire [7:0] t_r11_c4_11;
  wire [7:0] t_r11_c4_12;
  wire [7:0] t_r11_c5_0;
  wire [7:0] t_r11_c5_1;
  wire [7:0] t_r11_c5_2;
  wire [7:0] t_r11_c5_3;
  wire [7:0] t_r11_c5_4;
  wire [7:0] t_r11_c5_5;
  wire [7:0] t_r11_c5_6;
  wire [7:0] t_r11_c5_7;
  wire [7:0] t_r11_c5_8;
  wire [7:0] t_r11_c5_9;
  wire [7:0] t_r11_c5_10;
  wire [7:0] t_r11_c5_11;
  wire [7:0] t_r11_c5_12;
  wire [7:0] t_r11_c6_0;
  wire [7:0] t_r11_c6_1;
  wire [7:0] t_r11_c6_2;
  wire [7:0] t_r11_c6_3;
  wire [7:0] t_r11_c6_4;
  wire [7:0] t_r11_c6_5;
  wire [7:0] t_r11_c6_6;
  wire [7:0] t_r11_c6_7;
  wire [7:0] t_r11_c6_8;
  wire [7:0] t_r11_c6_9;
  wire [7:0] t_r11_c6_10;
  wire [7:0] t_r11_c6_11;
  wire [7:0] t_r11_c6_12;
  wire [7:0] t_r11_c7_0;
  wire [7:0] t_r11_c7_1;
  wire [7:0] t_r11_c7_2;
  wire [7:0] t_r11_c7_3;
  wire [7:0] t_r11_c7_4;
  wire [7:0] t_r11_c7_5;
  wire [7:0] t_r11_c7_6;
  wire [7:0] t_r11_c7_7;
  wire [7:0] t_r11_c7_8;
  wire [7:0] t_r11_c7_9;
  wire [7:0] t_r11_c7_10;
  wire [7:0] t_r11_c7_11;
  wire [7:0] t_r11_c7_12;
  wire [7:0] t_r11_c8_0;
  wire [7:0] t_r11_c8_1;
  wire [7:0] t_r11_c8_2;
  wire [7:0] t_r11_c8_3;
  wire [7:0] t_r11_c8_4;
  wire [7:0] t_r11_c8_5;
  wire [7:0] t_r11_c8_6;
  wire [7:0] t_r11_c8_7;
  wire [7:0] t_r11_c8_8;
  wire [7:0] t_r11_c8_9;
  wire [7:0] t_r11_c8_10;
  wire [7:0] t_r11_c8_11;
  wire [7:0] t_r11_c8_12;
  wire [7:0] t_r11_c9_0;
  wire [7:0] t_r11_c9_1;
  wire [7:0] t_r11_c9_2;
  wire [7:0] t_r11_c9_3;
  wire [7:0] t_r11_c9_4;
  wire [7:0] t_r11_c9_5;
  wire [7:0] t_r11_c9_6;
  wire [7:0] t_r11_c9_7;
  wire [7:0] t_r11_c9_8;
  wire [7:0] t_r11_c9_9;
  wire [7:0] t_r11_c9_10;
  wire [7:0] t_r11_c9_11;
  wire [7:0] t_r11_c9_12;
  wire [7:0] t_r11_c10_0;
  wire [7:0] t_r11_c10_1;
  wire [7:0] t_r11_c10_2;
  wire [7:0] t_r11_c10_3;
  wire [7:0] t_r11_c10_4;
  wire [7:0] t_r11_c10_5;
  wire [7:0] t_r11_c10_6;
  wire [7:0] t_r11_c10_7;
  wire [7:0] t_r11_c10_8;
  wire [7:0] t_r11_c10_9;
  wire [7:0] t_r11_c10_10;
  wire [7:0] t_r11_c10_11;
  wire [7:0] t_r11_c10_12;
  wire [7:0] t_r11_c11_0;
  wire [7:0] t_r11_c11_1;
  wire [7:0] t_r11_c11_2;
  wire [7:0] t_r11_c11_3;
  wire [7:0] t_r11_c11_4;
  wire [7:0] t_r11_c11_5;
  wire [7:0] t_r11_c11_6;
  wire [7:0] t_r11_c11_7;
  wire [7:0] t_r11_c11_8;
  wire [7:0] t_r11_c11_9;
  wire [7:0] t_r11_c11_10;
  wire [7:0] t_r11_c11_11;
  wire [7:0] t_r11_c11_12;
  wire [7:0] t_r11_c12_0;
  wire [7:0] t_r11_c12_1;
  wire [7:0] t_r11_c12_2;
  wire [7:0] t_r11_c12_3;
  wire [7:0] t_r11_c12_4;
  wire [7:0] t_r11_c12_5;
  wire [7:0] t_r11_c12_6;
  wire [7:0] t_r11_c12_7;
  wire [7:0] t_r11_c12_8;
  wire [7:0] t_r11_c12_9;
  wire [7:0] t_r11_c12_10;
  wire [7:0] t_r11_c12_11;
  wire [7:0] t_r11_c12_12;
  wire [7:0] t_r11_c13_0;
  wire [7:0] t_r11_c13_1;
  wire [7:0] t_r11_c13_2;
  wire [7:0] t_r11_c13_3;
  wire [7:0] t_r11_c13_4;
  wire [7:0] t_r11_c13_5;
  wire [7:0] t_r11_c13_6;
  wire [7:0] t_r11_c13_7;
  wire [7:0] t_r11_c13_8;
  wire [7:0] t_r11_c13_9;
  wire [7:0] t_r11_c13_10;
  wire [7:0] t_r11_c13_11;
  wire [7:0] t_r11_c13_12;
  wire [7:0] t_r11_c14_0;
  wire [7:0] t_r11_c14_1;
  wire [7:0] t_r11_c14_2;
  wire [7:0] t_r11_c14_3;
  wire [7:0] t_r11_c14_4;
  wire [7:0] t_r11_c14_5;
  wire [7:0] t_r11_c14_6;
  wire [7:0] t_r11_c14_7;
  wire [7:0] t_r11_c14_8;
  wire [7:0] t_r11_c14_9;
  wire [7:0] t_r11_c14_10;
  wire [7:0] t_r11_c14_11;
  wire [7:0] t_r11_c14_12;
  wire [7:0] t_r11_c15_0;
  wire [7:0] t_r11_c15_1;
  wire [7:0] t_r11_c15_2;
  wire [7:0] t_r11_c15_3;
  wire [7:0] t_r11_c15_4;
  wire [7:0] t_r11_c15_5;
  wire [7:0] t_r11_c15_6;
  wire [7:0] t_r11_c15_7;
  wire [7:0] t_r11_c15_8;
  wire [7:0] t_r11_c15_9;
  wire [7:0] t_r11_c15_10;
  wire [7:0] t_r11_c15_11;
  wire [7:0] t_r11_c15_12;
  wire [7:0] t_r11_c16_0;
  wire [7:0] t_r11_c16_1;
  wire [7:0] t_r11_c16_2;
  wire [7:0] t_r11_c16_3;
  wire [7:0] t_r11_c16_4;
  wire [7:0] t_r11_c16_5;
  wire [7:0] t_r11_c16_6;
  wire [7:0] t_r11_c16_7;
  wire [7:0] t_r11_c16_8;
  wire [7:0] t_r11_c16_9;
  wire [7:0] t_r11_c16_10;
  wire [7:0] t_r11_c16_11;
  wire [7:0] t_r11_c16_12;
  wire [7:0] t_r11_c17_0;
  wire [7:0] t_r11_c17_1;
  wire [7:0] t_r11_c17_2;
  wire [7:0] t_r11_c17_3;
  wire [7:0] t_r11_c17_4;
  wire [7:0] t_r11_c17_5;
  wire [7:0] t_r11_c17_6;
  wire [7:0] t_r11_c17_7;
  wire [7:0] t_r11_c17_8;
  wire [7:0] t_r11_c17_9;
  wire [7:0] t_r11_c17_10;
  wire [7:0] t_r11_c17_11;
  wire [7:0] t_r11_c17_12;
  wire [7:0] t_r11_c18_0;
  wire [7:0] t_r11_c18_1;
  wire [7:0] t_r11_c18_2;
  wire [7:0] t_r11_c18_3;
  wire [7:0] t_r11_c18_4;
  wire [7:0] t_r11_c18_5;
  wire [7:0] t_r11_c18_6;
  wire [7:0] t_r11_c18_7;
  wire [7:0] t_r11_c18_8;
  wire [7:0] t_r11_c18_9;
  wire [7:0] t_r11_c18_10;
  wire [7:0] t_r11_c18_11;
  wire [7:0] t_r11_c18_12;
  wire [7:0] t_r11_c19_0;
  wire [7:0] t_r11_c19_1;
  wire [7:0] t_r11_c19_2;
  wire [7:0] t_r11_c19_3;
  wire [7:0] t_r11_c19_4;
  wire [7:0] t_r11_c19_5;
  wire [7:0] t_r11_c19_6;
  wire [7:0] t_r11_c19_7;
  wire [7:0] t_r11_c19_8;
  wire [7:0] t_r11_c19_9;
  wire [7:0] t_r11_c19_10;
  wire [7:0] t_r11_c19_11;
  wire [7:0] t_r11_c19_12;
  wire [7:0] t_r11_c20_0;
  wire [7:0] t_r11_c20_1;
  wire [7:0] t_r11_c20_2;
  wire [7:0] t_r11_c20_3;
  wire [7:0] t_r11_c20_4;
  wire [7:0] t_r11_c20_5;
  wire [7:0] t_r11_c20_6;
  wire [7:0] t_r11_c20_7;
  wire [7:0] t_r11_c20_8;
  wire [7:0] t_r11_c20_9;
  wire [7:0] t_r11_c20_10;
  wire [7:0] t_r11_c20_11;
  wire [7:0] t_r11_c20_12;
  wire [7:0] t_r11_c21_0;
  wire [7:0] t_r11_c21_1;
  wire [7:0] t_r11_c21_2;
  wire [7:0] t_r11_c21_3;
  wire [7:0] t_r11_c21_4;
  wire [7:0] t_r11_c21_5;
  wire [7:0] t_r11_c21_6;
  wire [7:0] t_r11_c21_7;
  wire [7:0] t_r11_c21_8;
  wire [7:0] t_r11_c21_9;
  wire [7:0] t_r11_c21_10;
  wire [7:0] t_r11_c21_11;
  wire [7:0] t_r11_c21_12;
  wire [7:0] t_r11_c22_0;
  wire [7:0] t_r11_c22_1;
  wire [7:0] t_r11_c22_2;
  wire [7:0] t_r11_c22_3;
  wire [7:0] t_r11_c22_4;
  wire [7:0] t_r11_c22_5;
  wire [7:0] t_r11_c22_6;
  wire [7:0] t_r11_c22_7;
  wire [7:0] t_r11_c22_8;
  wire [7:0] t_r11_c22_9;
  wire [7:0] t_r11_c22_10;
  wire [7:0] t_r11_c22_11;
  wire [7:0] t_r11_c22_12;
  wire [7:0] t_r11_c23_0;
  wire [7:0] t_r11_c23_1;
  wire [7:0] t_r11_c23_2;
  wire [7:0] t_r11_c23_3;
  wire [7:0] t_r11_c23_4;
  wire [7:0] t_r11_c23_5;
  wire [7:0] t_r11_c23_6;
  wire [7:0] t_r11_c23_7;
  wire [7:0] t_r11_c23_8;
  wire [7:0] t_r11_c23_9;
  wire [7:0] t_r11_c23_10;
  wire [7:0] t_r11_c23_11;
  wire [7:0] t_r11_c23_12;
  wire [7:0] t_r11_c24_0;
  wire [7:0] t_r11_c24_1;
  wire [7:0] t_r11_c24_2;
  wire [7:0] t_r11_c24_3;
  wire [7:0] t_r11_c24_4;
  wire [7:0] t_r11_c24_5;
  wire [7:0] t_r11_c24_6;
  wire [7:0] t_r11_c24_7;
  wire [7:0] t_r11_c24_8;
  wire [7:0] t_r11_c24_9;
  wire [7:0] t_r11_c24_10;
  wire [7:0] t_r11_c24_11;
  wire [7:0] t_r11_c24_12;
  wire [7:0] t_r11_c25_0;
  wire [7:0] t_r11_c25_1;
  wire [7:0] t_r11_c25_2;
  wire [7:0] t_r11_c25_3;
  wire [7:0] t_r11_c25_4;
  wire [7:0] t_r11_c25_5;
  wire [7:0] t_r11_c25_6;
  wire [7:0] t_r11_c25_7;
  wire [7:0] t_r11_c25_8;
  wire [7:0] t_r11_c25_9;
  wire [7:0] t_r11_c25_10;
  wire [7:0] t_r11_c25_11;
  wire [7:0] t_r11_c25_12;
  wire [7:0] t_r11_c26_0;
  wire [7:0] t_r11_c26_1;
  wire [7:0] t_r11_c26_2;
  wire [7:0] t_r11_c26_3;
  wire [7:0] t_r11_c26_4;
  wire [7:0] t_r11_c26_5;
  wire [7:0] t_r11_c26_6;
  wire [7:0] t_r11_c26_7;
  wire [7:0] t_r11_c26_8;
  wire [7:0] t_r11_c26_9;
  wire [7:0] t_r11_c26_10;
  wire [7:0] t_r11_c26_11;
  wire [7:0] t_r11_c26_12;
  wire [7:0] t_r11_c27_0;
  wire [7:0] t_r11_c27_1;
  wire [7:0] t_r11_c27_2;
  wire [7:0] t_r11_c27_3;
  wire [7:0] t_r11_c27_4;
  wire [7:0] t_r11_c27_5;
  wire [7:0] t_r11_c27_6;
  wire [7:0] t_r11_c27_7;
  wire [7:0] t_r11_c27_8;
  wire [7:0] t_r11_c27_9;
  wire [7:0] t_r11_c27_10;
  wire [7:0] t_r11_c27_11;
  wire [7:0] t_r11_c27_12;
  wire [7:0] t_r11_c28_0;
  wire [7:0] t_r11_c28_1;
  wire [7:0] t_r11_c28_2;
  wire [7:0] t_r11_c28_3;
  wire [7:0] t_r11_c28_4;
  wire [7:0] t_r11_c28_5;
  wire [7:0] t_r11_c28_6;
  wire [7:0] t_r11_c28_7;
  wire [7:0] t_r11_c28_8;
  wire [7:0] t_r11_c28_9;
  wire [7:0] t_r11_c28_10;
  wire [7:0] t_r11_c28_11;
  wire [7:0] t_r11_c28_12;
  wire [7:0] t_r11_c29_0;
  wire [7:0] t_r11_c29_1;
  wire [7:0] t_r11_c29_2;
  wire [7:0] t_r11_c29_3;
  wire [7:0] t_r11_c29_4;
  wire [7:0] t_r11_c29_5;
  wire [7:0] t_r11_c29_6;
  wire [7:0] t_r11_c29_7;
  wire [7:0] t_r11_c29_8;
  wire [7:0] t_r11_c29_9;
  wire [7:0] t_r11_c29_10;
  wire [7:0] t_r11_c29_11;
  wire [7:0] t_r11_c29_12;
  wire [7:0] t_r11_c30_0;
  wire [7:0] t_r11_c30_1;
  wire [7:0] t_r11_c30_2;
  wire [7:0] t_r11_c30_3;
  wire [7:0] t_r11_c30_4;
  wire [7:0] t_r11_c30_5;
  wire [7:0] t_r11_c30_6;
  wire [7:0] t_r11_c30_7;
  wire [7:0] t_r11_c30_8;
  wire [7:0] t_r11_c30_9;
  wire [7:0] t_r11_c30_10;
  wire [7:0] t_r11_c30_11;
  wire [7:0] t_r11_c30_12;
  wire [7:0] t_r11_c31_0;
  wire [7:0] t_r11_c31_1;
  wire [7:0] t_r11_c31_2;
  wire [7:0] t_r11_c31_3;
  wire [7:0] t_r11_c31_4;
  wire [7:0] t_r11_c31_5;
  wire [7:0] t_r11_c31_6;
  wire [7:0] t_r11_c31_7;
  wire [7:0] t_r11_c31_8;
  wire [7:0] t_r11_c31_9;
  wire [7:0] t_r11_c31_10;
  wire [7:0] t_r11_c31_11;
  wire [7:0] t_r11_c31_12;
  wire [7:0] t_r11_c32_0;
  wire [7:0] t_r11_c32_1;
  wire [7:0] t_r11_c32_2;
  wire [7:0] t_r11_c32_3;
  wire [7:0] t_r11_c32_4;
  wire [7:0] t_r11_c32_5;
  wire [7:0] t_r11_c32_6;
  wire [7:0] t_r11_c32_7;
  wire [7:0] t_r11_c32_8;
  wire [7:0] t_r11_c32_9;
  wire [7:0] t_r11_c32_10;
  wire [7:0] t_r11_c32_11;
  wire [7:0] t_r11_c32_12;
  wire [7:0] t_r11_c33_0;
  wire [7:0] t_r11_c33_1;
  wire [7:0] t_r11_c33_2;
  wire [7:0] t_r11_c33_3;
  wire [7:0] t_r11_c33_4;
  wire [7:0] t_r11_c33_5;
  wire [7:0] t_r11_c33_6;
  wire [7:0] t_r11_c33_7;
  wire [7:0] t_r11_c33_8;
  wire [7:0] t_r11_c33_9;
  wire [7:0] t_r11_c33_10;
  wire [7:0] t_r11_c33_11;
  wire [7:0] t_r11_c33_12;
  wire [7:0] t_r11_c34_0;
  wire [7:0] t_r11_c34_1;
  wire [7:0] t_r11_c34_2;
  wire [7:0] t_r11_c34_3;
  wire [7:0] t_r11_c34_4;
  wire [7:0] t_r11_c34_5;
  wire [7:0] t_r11_c34_6;
  wire [7:0] t_r11_c34_7;
  wire [7:0] t_r11_c34_8;
  wire [7:0] t_r11_c34_9;
  wire [7:0] t_r11_c34_10;
  wire [7:0] t_r11_c34_11;
  wire [7:0] t_r11_c34_12;
  wire [7:0] t_r11_c35_0;
  wire [7:0] t_r11_c35_1;
  wire [7:0] t_r11_c35_2;
  wire [7:0] t_r11_c35_3;
  wire [7:0] t_r11_c35_4;
  wire [7:0] t_r11_c35_5;
  wire [7:0] t_r11_c35_6;
  wire [7:0] t_r11_c35_7;
  wire [7:0] t_r11_c35_8;
  wire [7:0] t_r11_c35_9;
  wire [7:0] t_r11_c35_10;
  wire [7:0] t_r11_c35_11;
  wire [7:0] t_r11_c35_12;
  wire [7:0] t_r11_c36_0;
  wire [7:0] t_r11_c36_1;
  wire [7:0] t_r11_c36_2;
  wire [7:0] t_r11_c36_3;
  wire [7:0] t_r11_c36_4;
  wire [7:0] t_r11_c36_5;
  wire [7:0] t_r11_c36_6;
  wire [7:0] t_r11_c36_7;
  wire [7:0] t_r11_c36_8;
  wire [7:0] t_r11_c36_9;
  wire [7:0] t_r11_c36_10;
  wire [7:0] t_r11_c36_11;
  wire [7:0] t_r11_c36_12;
  wire [7:0] t_r11_c37_0;
  wire [7:0] t_r11_c37_1;
  wire [7:0] t_r11_c37_2;
  wire [7:0] t_r11_c37_3;
  wire [7:0] t_r11_c37_4;
  wire [7:0] t_r11_c37_5;
  wire [7:0] t_r11_c37_6;
  wire [7:0] t_r11_c37_7;
  wire [7:0] t_r11_c37_8;
  wire [7:0] t_r11_c37_9;
  wire [7:0] t_r11_c37_10;
  wire [7:0] t_r11_c37_11;
  wire [7:0] t_r11_c37_12;
  wire [7:0] t_r11_c38_0;
  wire [7:0] t_r11_c38_1;
  wire [7:0] t_r11_c38_2;
  wire [7:0] t_r11_c38_3;
  wire [7:0] t_r11_c38_4;
  wire [7:0] t_r11_c38_5;
  wire [7:0] t_r11_c38_6;
  wire [7:0] t_r11_c38_7;
  wire [7:0] t_r11_c38_8;
  wire [7:0] t_r11_c38_9;
  wire [7:0] t_r11_c38_10;
  wire [7:0] t_r11_c38_11;
  wire [7:0] t_r11_c38_12;
  wire [7:0] t_r11_c39_0;
  wire [7:0] t_r11_c39_1;
  wire [7:0] t_r11_c39_2;
  wire [7:0] t_r11_c39_3;
  wire [7:0] t_r11_c39_4;
  wire [7:0] t_r11_c39_5;
  wire [7:0] t_r11_c39_6;
  wire [7:0] t_r11_c39_7;
  wire [7:0] t_r11_c39_8;
  wire [7:0] t_r11_c39_9;
  wire [7:0] t_r11_c39_10;
  wire [7:0] t_r11_c39_11;
  wire [7:0] t_r11_c39_12;
  wire [7:0] t_r11_c40_0;
  wire [7:0] t_r11_c40_1;
  wire [7:0] t_r11_c40_2;
  wire [7:0] t_r11_c40_3;
  wire [7:0] t_r11_c40_4;
  wire [7:0] t_r11_c40_5;
  wire [7:0] t_r11_c40_6;
  wire [7:0] t_r11_c40_7;
  wire [7:0] t_r11_c40_8;
  wire [7:0] t_r11_c40_9;
  wire [7:0] t_r11_c40_10;
  wire [7:0] t_r11_c40_11;
  wire [7:0] t_r11_c40_12;
  wire [7:0] t_r11_c41_0;
  wire [7:0] t_r11_c41_1;
  wire [7:0] t_r11_c41_2;
  wire [7:0] t_r11_c41_3;
  wire [7:0] t_r11_c41_4;
  wire [7:0] t_r11_c41_5;
  wire [7:0] t_r11_c41_6;
  wire [7:0] t_r11_c41_7;
  wire [7:0] t_r11_c41_8;
  wire [7:0] t_r11_c41_9;
  wire [7:0] t_r11_c41_10;
  wire [7:0] t_r11_c41_11;
  wire [7:0] t_r11_c41_12;
  wire [7:0] t_r11_c42_0;
  wire [7:0] t_r11_c42_1;
  wire [7:0] t_r11_c42_2;
  wire [7:0] t_r11_c42_3;
  wire [7:0] t_r11_c42_4;
  wire [7:0] t_r11_c42_5;
  wire [7:0] t_r11_c42_6;
  wire [7:0] t_r11_c42_7;
  wire [7:0] t_r11_c42_8;
  wire [7:0] t_r11_c42_9;
  wire [7:0] t_r11_c42_10;
  wire [7:0] t_r11_c42_11;
  wire [7:0] t_r11_c42_12;
  wire [7:0] t_r11_c43_0;
  wire [7:0] t_r11_c43_1;
  wire [7:0] t_r11_c43_2;
  wire [7:0] t_r11_c43_3;
  wire [7:0] t_r11_c43_4;
  wire [7:0] t_r11_c43_5;
  wire [7:0] t_r11_c43_6;
  wire [7:0] t_r11_c43_7;
  wire [7:0] t_r11_c43_8;
  wire [7:0] t_r11_c43_9;
  wire [7:0] t_r11_c43_10;
  wire [7:0] t_r11_c43_11;
  wire [7:0] t_r11_c43_12;
  wire [7:0] t_r11_c44_0;
  wire [7:0] t_r11_c44_1;
  wire [7:0] t_r11_c44_2;
  wire [7:0] t_r11_c44_3;
  wire [7:0] t_r11_c44_4;
  wire [7:0] t_r11_c44_5;
  wire [7:0] t_r11_c44_6;
  wire [7:0] t_r11_c44_7;
  wire [7:0] t_r11_c44_8;
  wire [7:0] t_r11_c44_9;
  wire [7:0] t_r11_c44_10;
  wire [7:0] t_r11_c44_11;
  wire [7:0] t_r11_c44_12;
  wire [7:0] t_r11_c45_0;
  wire [7:0] t_r11_c45_1;
  wire [7:0] t_r11_c45_2;
  wire [7:0] t_r11_c45_3;
  wire [7:0] t_r11_c45_4;
  wire [7:0] t_r11_c45_5;
  wire [7:0] t_r11_c45_6;
  wire [7:0] t_r11_c45_7;
  wire [7:0] t_r11_c45_8;
  wire [7:0] t_r11_c45_9;
  wire [7:0] t_r11_c45_10;
  wire [7:0] t_r11_c45_11;
  wire [7:0] t_r11_c45_12;
  wire [7:0] t_r11_c46_0;
  wire [7:0] t_r11_c46_1;
  wire [7:0] t_r11_c46_2;
  wire [7:0] t_r11_c46_3;
  wire [7:0] t_r11_c46_4;
  wire [7:0] t_r11_c46_5;
  wire [7:0] t_r11_c46_6;
  wire [7:0] t_r11_c46_7;
  wire [7:0] t_r11_c46_8;
  wire [7:0] t_r11_c46_9;
  wire [7:0] t_r11_c46_10;
  wire [7:0] t_r11_c46_11;
  wire [7:0] t_r11_c46_12;
  wire [7:0] t_r11_c47_0;
  wire [7:0] t_r11_c47_1;
  wire [7:0] t_r11_c47_2;
  wire [7:0] t_r11_c47_3;
  wire [7:0] t_r11_c47_4;
  wire [7:0] t_r11_c47_5;
  wire [7:0] t_r11_c47_6;
  wire [7:0] t_r11_c47_7;
  wire [7:0] t_r11_c47_8;
  wire [7:0] t_r11_c47_9;
  wire [7:0] t_r11_c47_10;
  wire [7:0] t_r11_c47_11;
  wire [7:0] t_r11_c47_12;
  wire [7:0] t_r11_c48_0;
  wire [7:0] t_r11_c48_1;
  wire [7:0] t_r11_c48_2;
  wire [7:0] t_r11_c48_3;
  wire [7:0] t_r11_c48_4;
  wire [7:0] t_r11_c48_5;
  wire [7:0] t_r11_c48_6;
  wire [7:0] t_r11_c48_7;
  wire [7:0] t_r11_c48_8;
  wire [7:0] t_r11_c48_9;
  wire [7:0] t_r11_c48_10;
  wire [7:0] t_r11_c48_11;
  wire [7:0] t_r11_c48_12;
  wire [7:0] t_r11_c49_0;
  wire [7:0] t_r11_c49_1;
  wire [7:0] t_r11_c49_2;
  wire [7:0] t_r11_c49_3;
  wire [7:0] t_r11_c49_4;
  wire [7:0] t_r11_c49_5;
  wire [7:0] t_r11_c49_6;
  wire [7:0] t_r11_c49_7;
  wire [7:0] t_r11_c49_8;
  wire [7:0] t_r11_c49_9;
  wire [7:0] t_r11_c49_10;
  wire [7:0] t_r11_c49_11;
  wire [7:0] t_r11_c49_12;
  wire [7:0] t_r11_c50_0;
  wire [7:0] t_r11_c50_1;
  wire [7:0] t_r11_c50_2;
  wire [7:0] t_r11_c50_3;
  wire [7:0] t_r11_c50_4;
  wire [7:0] t_r11_c50_5;
  wire [7:0] t_r11_c50_6;
  wire [7:0] t_r11_c50_7;
  wire [7:0] t_r11_c50_8;
  wire [7:0] t_r11_c50_9;
  wire [7:0] t_r11_c50_10;
  wire [7:0] t_r11_c50_11;
  wire [7:0] t_r11_c50_12;
  wire [7:0] t_r11_c51_0;
  wire [7:0] t_r11_c51_1;
  wire [7:0] t_r11_c51_2;
  wire [7:0] t_r11_c51_3;
  wire [7:0] t_r11_c51_4;
  wire [7:0] t_r11_c51_5;
  wire [7:0] t_r11_c51_6;
  wire [7:0] t_r11_c51_7;
  wire [7:0] t_r11_c51_8;
  wire [7:0] t_r11_c51_9;
  wire [7:0] t_r11_c51_10;
  wire [7:0] t_r11_c51_11;
  wire [7:0] t_r11_c51_12;
  wire [7:0] t_r11_c52_0;
  wire [7:0] t_r11_c52_1;
  wire [7:0] t_r11_c52_2;
  wire [7:0] t_r11_c52_3;
  wire [7:0] t_r11_c52_4;
  wire [7:0] t_r11_c52_5;
  wire [7:0] t_r11_c52_6;
  wire [7:0] t_r11_c52_7;
  wire [7:0] t_r11_c52_8;
  wire [7:0] t_r11_c52_9;
  wire [7:0] t_r11_c52_10;
  wire [7:0] t_r11_c52_11;
  wire [7:0] t_r11_c52_12;
  wire [7:0] t_r11_c53_0;
  wire [7:0] t_r11_c53_1;
  wire [7:0] t_r11_c53_2;
  wire [7:0] t_r11_c53_3;
  wire [7:0] t_r11_c53_4;
  wire [7:0] t_r11_c53_5;
  wire [7:0] t_r11_c53_6;
  wire [7:0] t_r11_c53_7;
  wire [7:0] t_r11_c53_8;
  wire [7:0] t_r11_c53_9;
  wire [7:0] t_r11_c53_10;
  wire [7:0] t_r11_c53_11;
  wire [7:0] t_r11_c53_12;
  wire [7:0] t_r11_c54_0;
  wire [7:0] t_r11_c54_1;
  wire [7:0] t_r11_c54_2;
  wire [7:0] t_r11_c54_3;
  wire [7:0] t_r11_c54_4;
  wire [7:0] t_r11_c54_5;
  wire [7:0] t_r11_c54_6;
  wire [7:0] t_r11_c54_7;
  wire [7:0] t_r11_c54_8;
  wire [7:0] t_r11_c54_9;
  wire [7:0] t_r11_c54_10;
  wire [7:0] t_r11_c54_11;
  wire [7:0] t_r11_c54_12;
  wire [7:0] t_r11_c55_0;
  wire [7:0] t_r11_c55_1;
  wire [7:0] t_r11_c55_2;
  wire [7:0] t_r11_c55_3;
  wire [7:0] t_r11_c55_4;
  wire [7:0] t_r11_c55_5;
  wire [7:0] t_r11_c55_6;
  wire [7:0] t_r11_c55_7;
  wire [7:0] t_r11_c55_8;
  wire [7:0] t_r11_c55_9;
  wire [7:0] t_r11_c55_10;
  wire [7:0] t_r11_c55_11;
  wire [7:0] t_r11_c55_12;
  wire [7:0] t_r11_c56_0;
  wire [7:0] t_r11_c56_1;
  wire [7:0] t_r11_c56_2;
  wire [7:0] t_r11_c56_3;
  wire [7:0] t_r11_c56_4;
  wire [7:0] t_r11_c56_5;
  wire [7:0] t_r11_c56_6;
  wire [7:0] t_r11_c56_7;
  wire [7:0] t_r11_c56_8;
  wire [7:0] t_r11_c56_9;
  wire [7:0] t_r11_c56_10;
  wire [7:0] t_r11_c56_11;
  wire [7:0] t_r11_c56_12;
  wire [7:0] t_r11_c57_0;
  wire [7:0] t_r11_c57_1;
  wire [7:0] t_r11_c57_2;
  wire [7:0] t_r11_c57_3;
  wire [7:0] t_r11_c57_4;
  wire [7:0] t_r11_c57_5;
  wire [7:0] t_r11_c57_6;
  wire [7:0] t_r11_c57_7;
  wire [7:0] t_r11_c57_8;
  wire [7:0] t_r11_c57_9;
  wire [7:0] t_r11_c57_10;
  wire [7:0] t_r11_c57_11;
  wire [7:0] t_r11_c57_12;
  wire [7:0] t_r11_c58_0;
  wire [7:0] t_r11_c58_1;
  wire [7:0] t_r11_c58_2;
  wire [7:0] t_r11_c58_3;
  wire [7:0] t_r11_c58_4;
  wire [7:0] t_r11_c58_5;
  wire [7:0] t_r11_c58_6;
  wire [7:0] t_r11_c58_7;
  wire [7:0] t_r11_c58_8;
  wire [7:0] t_r11_c58_9;
  wire [7:0] t_r11_c58_10;
  wire [7:0] t_r11_c58_11;
  wire [7:0] t_r11_c58_12;
  wire [7:0] t_r11_c59_0;
  wire [7:0] t_r11_c59_1;
  wire [7:0] t_r11_c59_2;
  wire [7:0] t_r11_c59_3;
  wire [7:0] t_r11_c59_4;
  wire [7:0] t_r11_c59_5;
  wire [7:0] t_r11_c59_6;
  wire [7:0] t_r11_c59_7;
  wire [7:0] t_r11_c59_8;
  wire [7:0] t_r11_c59_9;
  wire [7:0] t_r11_c59_10;
  wire [7:0] t_r11_c59_11;
  wire [7:0] t_r11_c59_12;
  wire [7:0] t_r11_c60_0;
  wire [7:0] t_r11_c60_1;
  wire [7:0] t_r11_c60_2;
  wire [7:0] t_r11_c60_3;
  wire [7:0] t_r11_c60_4;
  wire [7:0] t_r11_c60_5;
  wire [7:0] t_r11_c60_6;
  wire [7:0] t_r11_c60_7;
  wire [7:0] t_r11_c60_8;
  wire [7:0] t_r11_c60_9;
  wire [7:0] t_r11_c60_10;
  wire [7:0] t_r11_c60_11;
  wire [7:0] t_r11_c60_12;
  wire [7:0] t_r11_c61_0;
  wire [7:0] t_r11_c61_1;
  wire [7:0] t_r11_c61_2;
  wire [7:0] t_r11_c61_3;
  wire [7:0] t_r11_c61_4;
  wire [7:0] t_r11_c61_5;
  wire [7:0] t_r11_c61_6;
  wire [7:0] t_r11_c61_7;
  wire [7:0] t_r11_c61_8;
  wire [7:0] t_r11_c61_9;
  wire [7:0] t_r11_c61_10;
  wire [7:0] t_r11_c61_11;
  wire [7:0] t_r11_c61_12;
  wire [7:0] t_r11_c62_0;
  wire [7:0] t_r11_c62_1;
  wire [7:0] t_r11_c62_2;
  wire [7:0] t_r11_c62_3;
  wire [7:0] t_r11_c62_4;
  wire [7:0] t_r11_c62_5;
  wire [7:0] t_r11_c62_6;
  wire [7:0] t_r11_c62_7;
  wire [7:0] t_r11_c62_8;
  wire [7:0] t_r11_c62_9;
  wire [7:0] t_r11_c62_10;
  wire [7:0] t_r11_c62_11;
  wire [7:0] t_r11_c62_12;
  wire [7:0] t_r11_c63_0;
  wire [7:0] t_r11_c63_1;
  wire [7:0] t_r11_c63_2;
  wire [7:0] t_r11_c63_3;
  wire [7:0] t_r11_c63_4;
  wire [7:0] t_r11_c63_5;
  wire [7:0] t_r11_c63_6;
  wire [7:0] t_r11_c63_7;
  wire [7:0] t_r11_c63_8;
  wire [7:0] t_r11_c63_9;
  wire [7:0] t_r11_c63_10;
  wire [7:0] t_r11_c63_11;
  wire [7:0] t_r11_c63_12;
  wire [7:0] t_r11_c64_0;
  wire [7:0] t_r11_c64_1;
  wire [7:0] t_r11_c64_2;
  wire [7:0] t_r11_c64_3;
  wire [7:0] t_r11_c64_4;
  wire [7:0] t_r11_c64_5;
  wire [7:0] t_r11_c64_6;
  wire [7:0] t_r11_c64_7;
  wire [7:0] t_r11_c64_8;
  wire [7:0] t_r11_c64_9;
  wire [7:0] t_r11_c64_10;
  wire [7:0] t_r11_c64_11;
  wire [7:0] t_r11_c64_12;
  wire [7:0] t_r11_c65_0;
  wire [7:0] t_r11_c65_1;
  wire [7:0] t_r11_c65_2;
  wire [7:0] t_r11_c65_3;
  wire [7:0] t_r11_c65_4;
  wire [7:0] t_r11_c65_5;
  wire [7:0] t_r11_c65_6;
  wire [7:0] t_r11_c65_7;
  wire [7:0] t_r11_c65_8;
  wire [7:0] t_r11_c65_9;
  wire [7:0] t_r11_c65_10;
  wire [7:0] t_r11_c65_11;
  wire [7:0] t_r11_c65_12;
  wire [7:0] t_r12_c0_0;
  wire [7:0] t_r12_c0_1;
  wire [7:0] t_r12_c0_2;
  wire [7:0] t_r12_c0_3;
  wire [7:0] t_r12_c0_4;
  wire [7:0] t_r12_c0_5;
  wire [7:0] t_r12_c0_6;
  wire [7:0] t_r12_c0_7;
  wire [7:0] t_r12_c0_8;
  wire [7:0] t_r12_c0_9;
  wire [7:0] t_r12_c0_10;
  wire [7:0] t_r12_c0_11;
  wire [7:0] t_r12_c0_12;
  wire [7:0] t_r12_c1_0;
  wire [7:0] t_r12_c1_1;
  wire [7:0] t_r12_c1_2;
  wire [7:0] t_r12_c1_3;
  wire [7:0] t_r12_c1_4;
  wire [7:0] t_r12_c1_5;
  wire [7:0] t_r12_c1_6;
  wire [7:0] t_r12_c1_7;
  wire [7:0] t_r12_c1_8;
  wire [7:0] t_r12_c1_9;
  wire [7:0] t_r12_c1_10;
  wire [7:0] t_r12_c1_11;
  wire [7:0] t_r12_c1_12;
  wire [7:0] t_r12_c2_0;
  wire [7:0] t_r12_c2_1;
  wire [7:0] t_r12_c2_2;
  wire [7:0] t_r12_c2_3;
  wire [7:0] t_r12_c2_4;
  wire [7:0] t_r12_c2_5;
  wire [7:0] t_r12_c2_6;
  wire [7:0] t_r12_c2_7;
  wire [7:0] t_r12_c2_8;
  wire [7:0] t_r12_c2_9;
  wire [7:0] t_r12_c2_10;
  wire [7:0] t_r12_c2_11;
  wire [7:0] t_r12_c2_12;
  wire [7:0] t_r12_c3_0;
  wire [7:0] t_r12_c3_1;
  wire [7:0] t_r12_c3_2;
  wire [7:0] t_r12_c3_3;
  wire [7:0] t_r12_c3_4;
  wire [7:0] t_r12_c3_5;
  wire [7:0] t_r12_c3_6;
  wire [7:0] t_r12_c3_7;
  wire [7:0] t_r12_c3_8;
  wire [7:0] t_r12_c3_9;
  wire [7:0] t_r12_c3_10;
  wire [7:0] t_r12_c3_11;
  wire [7:0] t_r12_c3_12;
  wire [7:0] t_r12_c4_0;
  wire [7:0] t_r12_c4_1;
  wire [7:0] t_r12_c4_2;
  wire [7:0] t_r12_c4_3;
  wire [7:0] t_r12_c4_4;
  wire [7:0] t_r12_c4_5;
  wire [7:0] t_r12_c4_6;
  wire [7:0] t_r12_c4_7;
  wire [7:0] t_r12_c4_8;
  wire [7:0] t_r12_c4_9;
  wire [7:0] t_r12_c4_10;
  wire [7:0] t_r12_c4_11;
  wire [7:0] t_r12_c4_12;
  wire [7:0] t_r12_c5_0;
  wire [7:0] t_r12_c5_1;
  wire [7:0] t_r12_c5_2;
  wire [7:0] t_r12_c5_3;
  wire [7:0] t_r12_c5_4;
  wire [7:0] t_r12_c5_5;
  wire [7:0] t_r12_c5_6;
  wire [7:0] t_r12_c5_7;
  wire [7:0] t_r12_c5_8;
  wire [7:0] t_r12_c5_9;
  wire [7:0] t_r12_c5_10;
  wire [7:0] t_r12_c5_11;
  wire [7:0] t_r12_c5_12;
  wire [7:0] t_r12_c6_0;
  wire [7:0] t_r12_c6_1;
  wire [7:0] t_r12_c6_2;
  wire [7:0] t_r12_c6_3;
  wire [7:0] t_r12_c6_4;
  wire [7:0] t_r12_c6_5;
  wire [7:0] t_r12_c6_6;
  wire [7:0] t_r12_c6_7;
  wire [7:0] t_r12_c6_8;
  wire [7:0] t_r12_c6_9;
  wire [7:0] t_r12_c6_10;
  wire [7:0] t_r12_c6_11;
  wire [7:0] t_r12_c6_12;
  wire [7:0] t_r12_c7_0;
  wire [7:0] t_r12_c7_1;
  wire [7:0] t_r12_c7_2;
  wire [7:0] t_r12_c7_3;
  wire [7:0] t_r12_c7_4;
  wire [7:0] t_r12_c7_5;
  wire [7:0] t_r12_c7_6;
  wire [7:0] t_r12_c7_7;
  wire [7:0] t_r12_c7_8;
  wire [7:0] t_r12_c7_9;
  wire [7:0] t_r12_c7_10;
  wire [7:0] t_r12_c7_11;
  wire [7:0] t_r12_c7_12;
  wire [7:0] t_r12_c8_0;
  wire [7:0] t_r12_c8_1;
  wire [7:0] t_r12_c8_2;
  wire [7:0] t_r12_c8_3;
  wire [7:0] t_r12_c8_4;
  wire [7:0] t_r12_c8_5;
  wire [7:0] t_r12_c8_6;
  wire [7:0] t_r12_c8_7;
  wire [7:0] t_r12_c8_8;
  wire [7:0] t_r12_c8_9;
  wire [7:0] t_r12_c8_10;
  wire [7:0] t_r12_c8_11;
  wire [7:0] t_r12_c8_12;
  wire [7:0] t_r12_c9_0;
  wire [7:0] t_r12_c9_1;
  wire [7:0] t_r12_c9_2;
  wire [7:0] t_r12_c9_3;
  wire [7:0] t_r12_c9_4;
  wire [7:0] t_r12_c9_5;
  wire [7:0] t_r12_c9_6;
  wire [7:0] t_r12_c9_7;
  wire [7:0] t_r12_c9_8;
  wire [7:0] t_r12_c9_9;
  wire [7:0] t_r12_c9_10;
  wire [7:0] t_r12_c9_11;
  wire [7:0] t_r12_c9_12;
  wire [7:0] t_r12_c10_0;
  wire [7:0] t_r12_c10_1;
  wire [7:0] t_r12_c10_2;
  wire [7:0] t_r12_c10_3;
  wire [7:0] t_r12_c10_4;
  wire [7:0] t_r12_c10_5;
  wire [7:0] t_r12_c10_6;
  wire [7:0] t_r12_c10_7;
  wire [7:0] t_r12_c10_8;
  wire [7:0] t_r12_c10_9;
  wire [7:0] t_r12_c10_10;
  wire [7:0] t_r12_c10_11;
  wire [7:0] t_r12_c10_12;
  wire [7:0] t_r12_c11_0;
  wire [7:0] t_r12_c11_1;
  wire [7:0] t_r12_c11_2;
  wire [7:0] t_r12_c11_3;
  wire [7:0] t_r12_c11_4;
  wire [7:0] t_r12_c11_5;
  wire [7:0] t_r12_c11_6;
  wire [7:0] t_r12_c11_7;
  wire [7:0] t_r12_c11_8;
  wire [7:0] t_r12_c11_9;
  wire [7:0] t_r12_c11_10;
  wire [7:0] t_r12_c11_11;
  wire [7:0] t_r12_c11_12;
  wire [7:0] t_r12_c12_0;
  wire [7:0] t_r12_c12_1;
  wire [7:0] t_r12_c12_2;
  wire [7:0] t_r12_c12_3;
  wire [7:0] t_r12_c12_4;
  wire [7:0] t_r12_c12_5;
  wire [7:0] t_r12_c12_6;
  wire [7:0] t_r12_c12_7;
  wire [7:0] t_r12_c12_8;
  wire [7:0] t_r12_c12_9;
  wire [7:0] t_r12_c12_10;
  wire [7:0] t_r12_c12_11;
  wire [7:0] t_r12_c12_12;
  wire [7:0] t_r12_c13_0;
  wire [7:0] t_r12_c13_1;
  wire [7:0] t_r12_c13_2;
  wire [7:0] t_r12_c13_3;
  wire [7:0] t_r12_c13_4;
  wire [7:0] t_r12_c13_5;
  wire [7:0] t_r12_c13_6;
  wire [7:0] t_r12_c13_7;
  wire [7:0] t_r12_c13_8;
  wire [7:0] t_r12_c13_9;
  wire [7:0] t_r12_c13_10;
  wire [7:0] t_r12_c13_11;
  wire [7:0] t_r12_c13_12;
  wire [7:0] t_r12_c14_0;
  wire [7:0] t_r12_c14_1;
  wire [7:0] t_r12_c14_2;
  wire [7:0] t_r12_c14_3;
  wire [7:0] t_r12_c14_4;
  wire [7:0] t_r12_c14_5;
  wire [7:0] t_r12_c14_6;
  wire [7:0] t_r12_c14_7;
  wire [7:0] t_r12_c14_8;
  wire [7:0] t_r12_c14_9;
  wire [7:0] t_r12_c14_10;
  wire [7:0] t_r12_c14_11;
  wire [7:0] t_r12_c14_12;
  wire [7:0] t_r12_c15_0;
  wire [7:0] t_r12_c15_1;
  wire [7:0] t_r12_c15_2;
  wire [7:0] t_r12_c15_3;
  wire [7:0] t_r12_c15_4;
  wire [7:0] t_r12_c15_5;
  wire [7:0] t_r12_c15_6;
  wire [7:0] t_r12_c15_7;
  wire [7:0] t_r12_c15_8;
  wire [7:0] t_r12_c15_9;
  wire [7:0] t_r12_c15_10;
  wire [7:0] t_r12_c15_11;
  wire [7:0] t_r12_c15_12;
  wire [7:0] t_r12_c16_0;
  wire [7:0] t_r12_c16_1;
  wire [7:0] t_r12_c16_2;
  wire [7:0] t_r12_c16_3;
  wire [7:0] t_r12_c16_4;
  wire [7:0] t_r12_c16_5;
  wire [7:0] t_r12_c16_6;
  wire [7:0] t_r12_c16_7;
  wire [7:0] t_r12_c16_8;
  wire [7:0] t_r12_c16_9;
  wire [7:0] t_r12_c16_10;
  wire [7:0] t_r12_c16_11;
  wire [7:0] t_r12_c16_12;
  wire [7:0] t_r12_c17_0;
  wire [7:0] t_r12_c17_1;
  wire [7:0] t_r12_c17_2;
  wire [7:0] t_r12_c17_3;
  wire [7:0] t_r12_c17_4;
  wire [7:0] t_r12_c17_5;
  wire [7:0] t_r12_c17_6;
  wire [7:0] t_r12_c17_7;
  wire [7:0] t_r12_c17_8;
  wire [7:0] t_r12_c17_9;
  wire [7:0] t_r12_c17_10;
  wire [7:0] t_r12_c17_11;
  wire [7:0] t_r12_c17_12;
  wire [7:0] t_r12_c18_0;
  wire [7:0] t_r12_c18_1;
  wire [7:0] t_r12_c18_2;
  wire [7:0] t_r12_c18_3;
  wire [7:0] t_r12_c18_4;
  wire [7:0] t_r12_c18_5;
  wire [7:0] t_r12_c18_6;
  wire [7:0] t_r12_c18_7;
  wire [7:0] t_r12_c18_8;
  wire [7:0] t_r12_c18_9;
  wire [7:0] t_r12_c18_10;
  wire [7:0] t_r12_c18_11;
  wire [7:0] t_r12_c18_12;
  wire [7:0] t_r12_c19_0;
  wire [7:0] t_r12_c19_1;
  wire [7:0] t_r12_c19_2;
  wire [7:0] t_r12_c19_3;
  wire [7:0] t_r12_c19_4;
  wire [7:0] t_r12_c19_5;
  wire [7:0] t_r12_c19_6;
  wire [7:0] t_r12_c19_7;
  wire [7:0] t_r12_c19_8;
  wire [7:0] t_r12_c19_9;
  wire [7:0] t_r12_c19_10;
  wire [7:0] t_r12_c19_11;
  wire [7:0] t_r12_c19_12;
  wire [7:0] t_r12_c20_0;
  wire [7:0] t_r12_c20_1;
  wire [7:0] t_r12_c20_2;
  wire [7:0] t_r12_c20_3;
  wire [7:0] t_r12_c20_4;
  wire [7:0] t_r12_c20_5;
  wire [7:0] t_r12_c20_6;
  wire [7:0] t_r12_c20_7;
  wire [7:0] t_r12_c20_8;
  wire [7:0] t_r12_c20_9;
  wire [7:0] t_r12_c20_10;
  wire [7:0] t_r12_c20_11;
  wire [7:0] t_r12_c20_12;
  wire [7:0] t_r12_c21_0;
  wire [7:0] t_r12_c21_1;
  wire [7:0] t_r12_c21_2;
  wire [7:0] t_r12_c21_3;
  wire [7:0] t_r12_c21_4;
  wire [7:0] t_r12_c21_5;
  wire [7:0] t_r12_c21_6;
  wire [7:0] t_r12_c21_7;
  wire [7:0] t_r12_c21_8;
  wire [7:0] t_r12_c21_9;
  wire [7:0] t_r12_c21_10;
  wire [7:0] t_r12_c21_11;
  wire [7:0] t_r12_c21_12;
  wire [7:0] t_r12_c22_0;
  wire [7:0] t_r12_c22_1;
  wire [7:0] t_r12_c22_2;
  wire [7:0] t_r12_c22_3;
  wire [7:0] t_r12_c22_4;
  wire [7:0] t_r12_c22_5;
  wire [7:0] t_r12_c22_6;
  wire [7:0] t_r12_c22_7;
  wire [7:0] t_r12_c22_8;
  wire [7:0] t_r12_c22_9;
  wire [7:0] t_r12_c22_10;
  wire [7:0] t_r12_c22_11;
  wire [7:0] t_r12_c22_12;
  wire [7:0] t_r12_c23_0;
  wire [7:0] t_r12_c23_1;
  wire [7:0] t_r12_c23_2;
  wire [7:0] t_r12_c23_3;
  wire [7:0] t_r12_c23_4;
  wire [7:0] t_r12_c23_5;
  wire [7:0] t_r12_c23_6;
  wire [7:0] t_r12_c23_7;
  wire [7:0] t_r12_c23_8;
  wire [7:0] t_r12_c23_9;
  wire [7:0] t_r12_c23_10;
  wire [7:0] t_r12_c23_11;
  wire [7:0] t_r12_c23_12;
  wire [7:0] t_r12_c24_0;
  wire [7:0] t_r12_c24_1;
  wire [7:0] t_r12_c24_2;
  wire [7:0] t_r12_c24_3;
  wire [7:0] t_r12_c24_4;
  wire [7:0] t_r12_c24_5;
  wire [7:0] t_r12_c24_6;
  wire [7:0] t_r12_c24_7;
  wire [7:0] t_r12_c24_8;
  wire [7:0] t_r12_c24_9;
  wire [7:0] t_r12_c24_10;
  wire [7:0] t_r12_c24_11;
  wire [7:0] t_r12_c24_12;
  wire [7:0] t_r12_c25_0;
  wire [7:0] t_r12_c25_1;
  wire [7:0] t_r12_c25_2;
  wire [7:0] t_r12_c25_3;
  wire [7:0] t_r12_c25_4;
  wire [7:0] t_r12_c25_5;
  wire [7:0] t_r12_c25_6;
  wire [7:0] t_r12_c25_7;
  wire [7:0] t_r12_c25_8;
  wire [7:0] t_r12_c25_9;
  wire [7:0] t_r12_c25_10;
  wire [7:0] t_r12_c25_11;
  wire [7:0] t_r12_c25_12;
  wire [7:0] t_r12_c26_0;
  wire [7:0] t_r12_c26_1;
  wire [7:0] t_r12_c26_2;
  wire [7:0] t_r12_c26_3;
  wire [7:0] t_r12_c26_4;
  wire [7:0] t_r12_c26_5;
  wire [7:0] t_r12_c26_6;
  wire [7:0] t_r12_c26_7;
  wire [7:0] t_r12_c26_8;
  wire [7:0] t_r12_c26_9;
  wire [7:0] t_r12_c26_10;
  wire [7:0] t_r12_c26_11;
  wire [7:0] t_r12_c26_12;
  wire [7:0] t_r12_c27_0;
  wire [7:0] t_r12_c27_1;
  wire [7:0] t_r12_c27_2;
  wire [7:0] t_r12_c27_3;
  wire [7:0] t_r12_c27_4;
  wire [7:0] t_r12_c27_5;
  wire [7:0] t_r12_c27_6;
  wire [7:0] t_r12_c27_7;
  wire [7:0] t_r12_c27_8;
  wire [7:0] t_r12_c27_9;
  wire [7:0] t_r12_c27_10;
  wire [7:0] t_r12_c27_11;
  wire [7:0] t_r12_c27_12;
  wire [7:0] t_r12_c28_0;
  wire [7:0] t_r12_c28_1;
  wire [7:0] t_r12_c28_2;
  wire [7:0] t_r12_c28_3;
  wire [7:0] t_r12_c28_4;
  wire [7:0] t_r12_c28_5;
  wire [7:0] t_r12_c28_6;
  wire [7:0] t_r12_c28_7;
  wire [7:0] t_r12_c28_8;
  wire [7:0] t_r12_c28_9;
  wire [7:0] t_r12_c28_10;
  wire [7:0] t_r12_c28_11;
  wire [7:0] t_r12_c28_12;
  wire [7:0] t_r12_c29_0;
  wire [7:0] t_r12_c29_1;
  wire [7:0] t_r12_c29_2;
  wire [7:0] t_r12_c29_3;
  wire [7:0] t_r12_c29_4;
  wire [7:0] t_r12_c29_5;
  wire [7:0] t_r12_c29_6;
  wire [7:0] t_r12_c29_7;
  wire [7:0] t_r12_c29_8;
  wire [7:0] t_r12_c29_9;
  wire [7:0] t_r12_c29_10;
  wire [7:0] t_r12_c29_11;
  wire [7:0] t_r12_c29_12;
  wire [7:0] t_r12_c30_0;
  wire [7:0] t_r12_c30_1;
  wire [7:0] t_r12_c30_2;
  wire [7:0] t_r12_c30_3;
  wire [7:0] t_r12_c30_4;
  wire [7:0] t_r12_c30_5;
  wire [7:0] t_r12_c30_6;
  wire [7:0] t_r12_c30_7;
  wire [7:0] t_r12_c30_8;
  wire [7:0] t_r12_c30_9;
  wire [7:0] t_r12_c30_10;
  wire [7:0] t_r12_c30_11;
  wire [7:0] t_r12_c30_12;
  wire [7:0] t_r12_c31_0;
  wire [7:0] t_r12_c31_1;
  wire [7:0] t_r12_c31_2;
  wire [7:0] t_r12_c31_3;
  wire [7:0] t_r12_c31_4;
  wire [7:0] t_r12_c31_5;
  wire [7:0] t_r12_c31_6;
  wire [7:0] t_r12_c31_7;
  wire [7:0] t_r12_c31_8;
  wire [7:0] t_r12_c31_9;
  wire [7:0] t_r12_c31_10;
  wire [7:0] t_r12_c31_11;
  wire [7:0] t_r12_c31_12;
  wire [7:0] t_r12_c32_0;
  wire [7:0] t_r12_c32_1;
  wire [7:0] t_r12_c32_2;
  wire [7:0] t_r12_c32_3;
  wire [7:0] t_r12_c32_4;
  wire [7:0] t_r12_c32_5;
  wire [7:0] t_r12_c32_6;
  wire [7:0] t_r12_c32_7;
  wire [7:0] t_r12_c32_8;
  wire [7:0] t_r12_c32_9;
  wire [7:0] t_r12_c32_10;
  wire [7:0] t_r12_c32_11;
  wire [7:0] t_r12_c32_12;
  wire [7:0] t_r12_c33_0;
  wire [7:0] t_r12_c33_1;
  wire [7:0] t_r12_c33_2;
  wire [7:0] t_r12_c33_3;
  wire [7:0] t_r12_c33_4;
  wire [7:0] t_r12_c33_5;
  wire [7:0] t_r12_c33_6;
  wire [7:0] t_r12_c33_7;
  wire [7:0] t_r12_c33_8;
  wire [7:0] t_r12_c33_9;
  wire [7:0] t_r12_c33_10;
  wire [7:0] t_r12_c33_11;
  wire [7:0] t_r12_c33_12;
  wire [7:0] t_r12_c34_0;
  wire [7:0] t_r12_c34_1;
  wire [7:0] t_r12_c34_2;
  wire [7:0] t_r12_c34_3;
  wire [7:0] t_r12_c34_4;
  wire [7:0] t_r12_c34_5;
  wire [7:0] t_r12_c34_6;
  wire [7:0] t_r12_c34_7;
  wire [7:0] t_r12_c34_8;
  wire [7:0] t_r12_c34_9;
  wire [7:0] t_r12_c34_10;
  wire [7:0] t_r12_c34_11;
  wire [7:0] t_r12_c34_12;
  wire [7:0] t_r12_c35_0;
  wire [7:0] t_r12_c35_1;
  wire [7:0] t_r12_c35_2;
  wire [7:0] t_r12_c35_3;
  wire [7:0] t_r12_c35_4;
  wire [7:0] t_r12_c35_5;
  wire [7:0] t_r12_c35_6;
  wire [7:0] t_r12_c35_7;
  wire [7:0] t_r12_c35_8;
  wire [7:0] t_r12_c35_9;
  wire [7:0] t_r12_c35_10;
  wire [7:0] t_r12_c35_11;
  wire [7:0] t_r12_c35_12;
  wire [7:0] t_r12_c36_0;
  wire [7:0] t_r12_c36_1;
  wire [7:0] t_r12_c36_2;
  wire [7:0] t_r12_c36_3;
  wire [7:0] t_r12_c36_4;
  wire [7:0] t_r12_c36_5;
  wire [7:0] t_r12_c36_6;
  wire [7:0] t_r12_c36_7;
  wire [7:0] t_r12_c36_8;
  wire [7:0] t_r12_c36_9;
  wire [7:0] t_r12_c36_10;
  wire [7:0] t_r12_c36_11;
  wire [7:0] t_r12_c36_12;
  wire [7:0] t_r12_c37_0;
  wire [7:0] t_r12_c37_1;
  wire [7:0] t_r12_c37_2;
  wire [7:0] t_r12_c37_3;
  wire [7:0] t_r12_c37_4;
  wire [7:0] t_r12_c37_5;
  wire [7:0] t_r12_c37_6;
  wire [7:0] t_r12_c37_7;
  wire [7:0] t_r12_c37_8;
  wire [7:0] t_r12_c37_9;
  wire [7:0] t_r12_c37_10;
  wire [7:0] t_r12_c37_11;
  wire [7:0] t_r12_c37_12;
  wire [7:0] t_r12_c38_0;
  wire [7:0] t_r12_c38_1;
  wire [7:0] t_r12_c38_2;
  wire [7:0] t_r12_c38_3;
  wire [7:0] t_r12_c38_4;
  wire [7:0] t_r12_c38_5;
  wire [7:0] t_r12_c38_6;
  wire [7:0] t_r12_c38_7;
  wire [7:0] t_r12_c38_8;
  wire [7:0] t_r12_c38_9;
  wire [7:0] t_r12_c38_10;
  wire [7:0] t_r12_c38_11;
  wire [7:0] t_r12_c38_12;
  wire [7:0] t_r12_c39_0;
  wire [7:0] t_r12_c39_1;
  wire [7:0] t_r12_c39_2;
  wire [7:0] t_r12_c39_3;
  wire [7:0] t_r12_c39_4;
  wire [7:0] t_r12_c39_5;
  wire [7:0] t_r12_c39_6;
  wire [7:0] t_r12_c39_7;
  wire [7:0] t_r12_c39_8;
  wire [7:0] t_r12_c39_9;
  wire [7:0] t_r12_c39_10;
  wire [7:0] t_r12_c39_11;
  wire [7:0] t_r12_c39_12;
  wire [7:0] t_r12_c40_0;
  wire [7:0] t_r12_c40_1;
  wire [7:0] t_r12_c40_2;
  wire [7:0] t_r12_c40_3;
  wire [7:0] t_r12_c40_4;
  wire [7:0] t_r12_c40_5;
  wire [7:0] t_r12_c40_6;
  wire [7:0] t_r12_c40_7;
  wire [7:0] t_r12_c40_8;
  wire [7:0] t_r12_c40_9;
  wire [7:0] t_r12_c40_10;
  wire [7:0] t_r12_c40_11;
  wire [7:0] t_r12_c40_12;
  wire [7:0] t_r12_c41_0;
  wire [7:0] t_r12_c41_1;
  wire [7:0] t_r12_c41_2;
  wire [7:0] t_r12_c41_3;
  wire [7:0] t_r12_c41_4;
  wire [7:0] t_r12_c41_5;
  wire [7:0] t_r12_c41_6;
  wire [7:0] t_r12_c41_7;
  wire [7:0] t_r12_c41_8;
  wire [7:0] t_r12_c41_9;
  wire [7:0] t_r12_c41_10;
  wire [7:0] t_r12_c41_11;
  wire [7:0] t_r12_c41_12;
  wire [7:0] t_r12_c42_0;
  wire [7:0] t_r12_c42_1;
  wire [7:0] t_r12_c42_2;
  wire [7:0] t_r12_c42_3;
  wire [7:0] t_r12_c42_4;
  wire [7:0] t_r12_c42_5;
  wire [7:0] t_r12_c42_6;
  wire [7:0] t_r12_c42_7;
  wire [7:0] t_r12_c42_8;
  wire [7:0] t_r12_c42_9;
  wire [7:0] t_r12_c42_10;
  wire [7:0] t_r12_c42_11;
  wire [7:0] t_r12_c42_12;
  wire [7:0] t_r12_c43_0;
  wire [7:0] t_r12_c43_1;
  wire [7:0] t_r12_c43_2;
  wire [7:0] t_r12_c43_3;
  wire [7:0] t_r12_c43_4;
  wire [7:0] t_r12_c43_5;
  wire [7:0] t_r12_c43_6;
  wire [7:0] t_r12_c43_7;
  wire [7:0] t_r12_c43_8;
  wire [7:0] t_r12_c43_9;
  wire [7:0] t_r12_c43_10;
  wire [7:0] t_r12_c43_11;
  wire [7:0] t_r12_c43_12;
  wire [7:0] t_r12_c44_0;
  wire [7:0] t_r12_c44_1;
  wire [7:0] t_r12_c44_2;
  wire [7:0] t_r12_c44_3;
  wire [7:0] t_r12_c44_4;
  wire [7:0] t_r12_c44_5;
  wire [7:0] t_r12_c44_6;
  wire [7:0] t_r12_c44_7;
  wire [7:0] t_r12_c44_8;
  wire [7:0] t_r12_c44_9;
  wire [7:0] t_r12_c44_10;
  wire [7:0] t_r12_c44_11;
  wire [7:0] t_r12_c44_12;
  wire [7:0] t_r12_c45_0;
  wire [7:0] t_r12_c45_1;
  wire [7:0] t_r12_c45_2;
  wire [7:0] t_r12_c45_3;
  wire [7:0] t_r12_c45_4;
  wire [7:0] t_r12_c45_5;
  wire [7:0] t_r12_c45_6;
  wire [7:0] t_r12_c45_7;
  wire [7:0] t_r12_c45_8;
  wire [7:0] t_r12_c45_9;
  wire [7:0] t_r12_c45_10;
  wire [7:0] t_r12_c45_11;
  wire [7:0] t_r12_c45_12;
  wire [7:0] t_r12_c46_0;
  wire [7:0] t_r12_c46_1;
  wire [7:0] t_r12_c46_2;
  wire [7:0] t_r12_c46_3;
  wire [7:0] t_r12_c46_4;
  wire [7:0] t_r12_c46_5;
  wire [7:0] t_r12_c46_6;
  wire [7:0] t_r12_c46_7;
  wire [7:0] t_r12_c46_8;
  wire [7:0] t_r12_c46_9;
  wire [7:0] t_r12_c46_10;
  wire [7:0] t_r12_c46_11;
  wire [7:0] t_r12_c46_12;
  wire [7:0] t_r12_c47_0;
  wire [7:0] t_r12_c47_1;
  wire [7:0] t_r12_c47_2;
  wire [7:0] t_r12_c47_3;
  wire [7:0] t_r12_c47_4;
  wire [7:0] t_r12_c47_5;
  wire [7:0] t_r12_c47_6;
  wire [7:0] t_r12_c47_7;
  wire [7:0] t_r12_c47_8;
  wire [7:0] t_r12_c47_9;
  wire [7:0] t_r12_c47_10;
  wire [7:0] t_r12_c47_11;
  wire [7:0] t_r12_c47_12;
  wire [7:0] t_r12_c48_0;
  wire [7:0] t_r12_c48_1;
  wire [7:0] t_r12_c48_2;
  wire [7:0] t_r12_c48_3;
  wire [7:0] t_r12_c48_4;
  wire [7:0] t_r12_c48_5;
  wire [7:0] t_r12_c48_6;
  wire [7:0] t_r12_c48_7;
  wire [7:0] t_r12_c48_8;
  wire [7:0] t_r12_c48_9;
  wire [7:0] t_r12_c48_10;
  wire [7:0] t_r12_c48_11;
  wire [7:0] t_r12_c48_12;
  wire [7:0] t_r12_c49_0;
  wire [7:0] t_r12_c49_1;
  wire [7:0] t_r12_c49_2;
  wire [7:0] t_r12_c49_3;
  wire [7:0] t_r12_c49_4;
  wire [7:0] t_r12_c49_5;
  wire [7:0] t_r12_c49_6;
  wire [7:0] t_r12_c49_7;
  wire [7:0] t_r12_c49_8;
  wire [7:0] t_r12_c49_9;
  wire [7:0] t_r12_c49_10;
  wire [7:0] t_r12_c49_11;
  wire [7:0] t_r12_c49_12;
  wire [7:0] t_r12_c50_0;
  wire [7:0] t_r12_c50_1;
  wire [7:0] t_r12_c50_2;
  wire [7:0] t_r12_c50_3;
  wire [7:0] t_r12_c50_4;
  wire [7:0] t_r12_c50_5;
  wire [7:0] t_r12_c50_6;
  wire [7:0] t_r12_c50_7;
  wire [7:0] t_r12_c50_8;
  wire [7:0] t_r12_c50_9;
  wire [7:0] t_r12_c50_10;
  wire [7:0] t_r12_c50_11;
  wire [7:0] t_r12_c50_12;
  wire [7:0] t_r12_c51_0;
  wire [7:0] t_r12_c51_1;
  wire [7:0] t_r12_c51_2;
  wire [7:0] t_r12_c51_3;
  wire [7:0] t_r12_c51_4;
  wire [7:0] t_r12_c51_5;
  wire [7:0] t_r12_c51_6;
  wire [7:0] t_r12_c51_7;
  wire [7:0] t_r12_c51_8;
  wire [7:0] t_r12_c51_9;
  wire [7:0] t_r12_c51_10;
  wire [7:0] t_r12_c51_11;
  wire [7:0] t_r12_c51_12;
  wire [7:0] t_r12_c52_0;
  wire [7:0] t_r12_c52_1;
  wire [7:0] t_r12_c52_2;
  wire [7:0] t_r12_c52_3;
  wire [7:0] t_r12_c52_4;
  wire [7:0] t_r12_c52_5;
  wire [7:0] t_r12_c52_6;
  wire [7:0] t_r12_c52_7;
  wire [7:0] t_r12_c52_8;
  wire [7:0] t_r12_c52_9;
  wire [7:0] t_r12_c52_10;
  wire [7:0] t_r12_c52_11;
  wire [7:0] t_r12_c52_12;
  wire [7:0] t_r12_c53_0;
  wire [7:0] t_r12_c53_1;
  wire [7:0] t_r12_c53_2;
  wire [7:0] t_r12_c53_3;
  wire [7:0] t_r12_c53_4;
  wire [7:0] t_r12_c53_5;
  wire [7:0] t_r12_c53_6;
  wire [7:0] t_r12_c53_7;
  wire [7:0] t_r12_c53_8;
  wire [7:0] t_r12_c53_9;
  wire [7:0] t_r12_c53_10;
  wire [7:0] t_r12_c53_11;
  wire [7:0] t_r12_c53_12;
  wire [7:0] t_r12_c54_0;
  wire [7:0] t_r12_c54_1;
  wire [7:0] t_r12_c54_2;
  wire [7:0] t_r12_c54_3;
  wire [7:0] t_r12_c54_4;
  wire [7:0] t_r12_c54_5;
  wire [7:0] t_r12_c54_6;
  wire [7:0] t_r12_c54_7;
  wire [7:0] t_r12_c54_8;
  wire [7:0] t_r12_c54_9;
  wire [7:0] t_r12_c54_10;
  wire [7:0] t_r12_c54_11;
  wire [7:0] t_r12_c54_12;
  wire [7:0] t_r12_c55_0;
  wire [7:0] t_r12_c55_1;
  wire [7:0] t_r12_c55_2;
  wire [7:0] t_r12_c55_3;
  wire [7:0] t_r12_c55_4;
  wire [7:0] t_r12_c55_5;
  wire [7:0] t_r12_c55_6;
  wire [7:0] t_r12_c55_7;
  wire [7:0] t_r12_c55_8;
  wire [7:0] t_r12_c55_9;
  wire [7:0] t_r12_c55_10;
  wire [7:0] t_r12_c55_11;
  wire [7:0] t_r12_c55_12;
  wire [7:0] t_r12_c56_0;
  wire [7:0] t_r12_c56_1;
  wire [7:0] t_r12_c56_2;
  wire [7:0] t_r12_c56_3;
  wire [7:0] t_r12_c56_4;
  wire [7:0] t_r12_c56_5;
  wire [7:0] t_r12_c56_6;
  wire [7:0] t_r12_c56_7;
  wire [7:0] t_r12_c56_8;
  wire [7:0] t_r12_c56_9;
  wire [7:0] t_r12_c56_10;
  wire [7:0] t_r12_c56_11;
  wire [7:0] t_r12_c56_12;
  wire [7:0] t_r12_c57_0;
  wire [7:0] t_r12_c57_1;
  wire [7:0] t_r12_c57_2;
  wire [7:0] t_r12_c57_3;
  wire [7:0] t_r12_c57_4;
  wire [7:0] t_r12_c57_5;
  wire [7:0] t_r12_c57_6;
  wire [7:0] t_r12_c57_7;
  wire [7:0] t_r12_c57_8;
  wire [7:0] t_r12_c57_9;
  wire [7:0] t_r12_c57_10;
  wire [7:0] t_r12_c57_11;
  wire [7:0] t_r12_c57_12;
  wire [7:0] t_r12_c58_0;
  wire [7:0] t_r12_c58_1;
  wire [7:0] t_r12_c58_2;
  wire [7:0] t_r12_c58_3;
  wire [7:0] t_r12_c58_4;
  wire [7:0] t_r12_c58_5;
  wire [7:0] t_r12_c58_6;
  wire [7:0] t_r12_c58_7;
  wire [7:0] t_r12_c58_8;
  wire [7:0] t_r12_c58_9;
  wire [7:0] t_r12_c58_10;
  wire [7:0] t_r12_c58_11;
  wire [7:0] t_r12_c58_12;
  wire [7:0] t_r12_c59_0;
  wire [7:0] t_r12_c59_1;
  wire [7:0] t_r12_c59_2;
  wire [7:0] t_r12_c59_3;
  wire [7:0] t_r12_c59_4;
  wire [7:0] t_r12_c59_5;
  wire [7:0] t_r12_c59_6;
  wire [7:0] t_r12_c59_7;
  wire [7:0] t_r12_c59_8;
  wire [7:0] t_r12_c59_9;
  wire [7:0] t_r12_c59_10;
  wire [7:0] t_r12_c59_11;
  wire [7:0] t_r12_c59_12;
  wire [7:0] t_r12_c60_0;
  wire [7:0] t_r12_c60_1;
  wire [7:0] t_r12_c60_2;
  wire [7:0] t_r12_c60_3;
  wire [7:0] t_r12_c60_4;
  wire [7:0] t_r12_c60_5;
  wire [7:0] t_r12_c60_6;
  wire [7:0] t_r12_c60_7;
  wire [7:0] t_r12_c60_8;
  wire [7:0] t_r12_c60_9;
  wire [7:0] t_r12_c60_10;
  wire [7:0] t_r12_c60_11;
  wire [7:0] t_r12_c60_12;
  wire [7:0] t_r12_c61_0;
  wire [7:0] t_r12_c61_1;
  wire [7:0] t_r12_c61_2;
  wire [7:0] t_r12_c61_3;
  wire [7:0] t_r12_c61_4;
  wire [7:0] t_r12_c61_5;
  wire [7:0] t_r12_c61_6;
  wire [7:0] t_r12_c61_7;
  wire [7:0] t_r12_c61_8;
  wire [7:0] t_r12_c61_9;
  wire [7:0] t_r12_c61_10;
  wire [7:0] t_r12_c61_11;
  wire [7:0] t_r12_c61_12;
  wire [7:0] t_r12_c62_0;
  wire [7:0] t_r12_c62_1;
  wire [7:0] t_r12_c62_2;
  wire [7:0] t_r12_c62_3;
  wire [7:0] t_r12_c62_4;
  wire [7:0] t_r12_c62_5;
  wire [7:0] t_r12_c62_6;
  wire [7:0] t_r12_c62_7;
  wire [7:0] t_r12_c62_8;
  wire [7:0] t_r12_c62_9;
  wire [7:0] t_r12_c62_10;
  wire [7:0] t_r12_c62_11;
  wire [7:0] t_r12_c62_12;
  wire [7:0] t_r12_c63_0;
  wire [7:0] t_r12_c63_1;
  wire [7:0] t_r12_c63_2;
  wire [7:0] t_r12_c63_3;
  wire [7:0] t_r12_c63_4;
  wire [7:0] t_r12_c63_5;
  wire [7:0] t_r12_c63_6;
  wire [7:0] t_r12_c63_7;
  wire [7:0] t_r12_c63_8;
  wire [7:0] t_r12_c63_9;
  wire [7:0] t_r12_c63_10;
  wire [7:0] t_r12_c63_11;
  wire [7:0] t_r12_c63_12;
  wire [7:0] t_r12_c64_0;
  wire [7:0] t_r12_c64_1;
  wire [7:0] t_r12_c64_2;
  wire [7:0] t_r12_c64_3;
  wire [7:0] t_r12_c64_4;
  wire [7:0] t_r12_c64_5;
  wire [7:0] t_r12_c64_6;
  wire [7:0] t_r12_c64_7;
  wire [7:0] t_r12_c64_8;
  wire [7:0] t_r12_c64_9;
  wire [7:0] t_r12_c64_10;
  wire [7:0] t_r12_c64_11;
  wire [7:0] t_r12_c64_12;
  wire [7:0] t_r12_c65_0;
  wire [7:0] t_r12_c65_1;
  wire [7:0] t_r12_c65_2;
  wire [7:0] t_r12_c65_3;
  wire [7:0] t_r12_c65_4;
  wire [7:0] t_r12_c65_5;
  wire [7:0] t_r12_c65_6;
  wire [7:0] t_r12_c65_7;
  wire [7:0] t_r12_c65_8;
  wire [7:0] t_r12_c65_9;
  wire [7:0] t_r12_c65_10;
  wire [7:0] t_r12_c65_11;
  wire [7:0] t_r12_c65_12;
  wire [7:0] t_r13_c0_0;
  wire [7:0] t_r13_c0_1;
  wire [7:0] t_r13_c0_2;
  wire [7:0] t_r13_c0_3;
  wire [7:0] t_r13_c0_4;
  wire [7:0] t_r13_c0_5;
  wire [7:0] t_r13_c0_6;
  wire [7:0] t_r13_c0_7;
  wire [7:0] t_r13_c0_8;
  wire [7:0] t_r13_c0_9;
  wire [7:0] t_r13_c0_10;
  wire [7:0] t_r13_c0_11;
  wire [7:0] t_r13_c0_12;
  wire [7:0] t_r13_c1_0;
  wire [7:0] t_r13_c1_1;
  wire [7:0] t_r13_c1_2;
  wire [7:0] t_r13_c1_3;
  wire [7:0] t_r13_c1_4;
  wire [7:0] t_r13_c1_5;
  wire [7:0] t_r13_c1_6;
  wire [7:0] t_r13_c1_7;
  wire [7:0] t_r13_c1_8;
  wire [7:0] t_r13_c1_9;
  wire [7:0] t_r13_c1_10;
  wire [7:0] t_r13_c1_11;
  wire [7:0] t_r13_c1_12;
  wire [7:0] t_r13_c2_0;
  wire [7:0] t_r13_c2_1;
  wire [7:0] t_r13_c2_2;
  wire [7:0] t_r13_c2_3;
  wire [7:0] t_r13_c2_4;
  wire [7:0] t_r13_c2_5;
  wire [7:0] t_r13_c2_6;
  wire [7:0] t_r13_c2_7;
  wire [7:0] t_r13_c2_8;
  wire [7:0] t_r13_c2_9;
  wire [7:0] t_r13_c2_10;
  wire [7:0] t_r13_c2_11;
  wire [7:0] t_r13_c2_12;
  wire [7:0] t_r13_c3_0;
  wire [7:0] t_r13_c3_1;
  wire [7:0] t_r13_c3_2;
  wire [7:0] t_r13_c3_3;
  wire [7:0] t_r13_c3_4;
  wire [7:0] t_r13_c3_5;
  wire [7:0] t_r13_c3_6;
  wire [7:0] t_r13_c3_7;
  wire [7:0] t_r13_c3_8;
  wire [7:0] t_r13_c3_9;
  wire [7:0] t_r13_c3_10;
  wire [7:0] t_r13_c3_11;
  wire [7:0] t_r13_c3_12;
  wire [7:0] t_r13_c4_0;
  wire [7:0] t_r13_c4_1;
  wire [7:0] t_r13_c4_2;
  wire [7:0] t_r13_c4_3;
  wire [7:0] t_r13_c4_4;
  wire [7:0] t_r13_c4_5;
  wire [7:0] t_r13_c4_6;
  wire [7:0] t_r13_c4_7;
  wire [7:0] t_r13_c4_8;
  wire [7:0] t_r13_c4_9;
  wire [7:0] t_r13_c4_10;
  wire [7:0] t_r13_c4_11;
  wire [7:0] t_r13_c4_12;
  wire [7:0] t_r13_c5_0;
  wire [7:0] t_r13_c5_1;
  wire [7:0] t_r13_c5_2;
  wire [7:0] t_r13_c5_3;
  wire [7:0] t_r13_c5_4;
  wire [7:0] t_r13_c5_5;
  wire [7:0] t_r13_c5_6;
  wire [7:0] t_r13_c5_7;
  wire [7:0] t_r13_c5_8;
  wire [7:0] t_r13_c5_9;
  wire [7:0] t_r13_c5_10;
  wire [7:0] t_r13_c5_11;
  wire [7:0] t_r13_c5_12;
  wire [7:0] t_r13_c6_0;
  wire [7:0] t_r13_c6_1;
  wire [7:0] t_r13_c6_2;
  wire [7:0] t_r13_c6_3;
  wire [7:0] t_r13_c6_4;
  wire [7:0] t_r13_c6_5;
  wire [7:0] t_r13_c6_6;
  wire [7:0] t_r13_c6_7;
  wire [7:0] t_r13_c6_8;
  wire [7:0] t_r13_c6_9;
  wire [7:0] t_r13_c6_10;
  wire [7:0] t_r13_c6_11;
  wire [7:0] t_r13_c6_12;
  wire [7:0] t_r13_c7_0;
  wire [7:0] t_r13_c7_1;
  wire [7:0] t_r13_c7_2;
  wire [7:0] t_r13_c7_3;
  wire [7:0] t_r13_c7_4;
  wire [7:0] t_r13_c7_5;
  wire [7:0] t_r13_c7_6;
  wire [7:0] t_r13_c7_7;
  wire [7:0] t_r13_c7_8;
  wire [7:0] t_r13_c7_9;
  wire [7:0] t_r13_c7_10;
  wire [7:0] t_r13_c7_11;
  wire [7:0] t_r13_c7_12;
  wire [7:0] t_r13_c8_0;
  wire [7:0] t_r13_c8_1;
  wire [7:0] t_r13_c8_2;
  wire [7:0] t_r13_c8_3;
  wire [7:0] t_r13_c8_4;
  wire [7:0] t_r13_c8_5;
  wire [7:0] t_r13_c8_6;
  wire [7:0] t_r13_c8_7;
  wire [7:0] t_r13_c8_8;
  wire [7:0] t_r13_c8_9;
  wire [7:0] t_r13_c8_10;
  wire [7:0] t_r13_c8_11;
  wire [7:0] t_r13_c8_12;
  wire [7:0] t_r13_c9_0;
  wire [7:0] t_r13_c9_1;
  wire [7:0] t_r13_c9_2;
  wire [7:0] t_r13_c9_3;
  wire [7:0] t_r13_c9_4;
  wire [7:0] t_r13_c9_5;
  wire [7:0] t_r13_c9_6;
  wire [7:0] t_r13_c9_7;
  wire [7:0] t_r13_c9_8;
  wire [7:0] t_r13_c9_9;
  wire [7:0] t_r13_c9_10;
  wire [7:0] t_r13_c9_11;
  wire [7:0] t_r13_c9_12;
  wire [7:0] t_r13_c10_0;
  wire [7:0] t_r13_c10_1;
  wire [7:0] t_r13_c10_2;
  wire [7:0] t_r13_c10_3;
  wire [7:0] t_r13_c10_4;
  wire [7:0] t_r13_c10_5;
  wire [7:0] t_r13_c10_6;
  wire [7:0] t_r13_c10_7;
  wire [7:0] t_r13_c10_8;
  wire [7:0] t_r13_c10_9;
  wire [7:0] t_r13_c10_10;
  wire [7:0] t_r13_c10_11;
  wire [7:0] t_r13_c10_12;
  wire [7:0] t_r13_c11_0;
  wire [7:0] t_r13_c11_1;
  wire [7:0] t_r13_c11_2;
  wire [7:0] t_r13_c11_3;
  wire [7:0] t_r13_c11_4;
  wire [7:0] t_r13_c11_5;
  wire [7:0] t_r13_c11_6;
  wire [7:0] t_r13_c11_7;
  wire [7:0] t_r13_c11_8;
  wire [7:0] t_r13_c11_9;
  wire [7:0] t_r13_c11_10;
  wire [7:0] t_r13_c11_11;
  wire [7:0] t_r13_c11_12;
  wire [7:0] t_r13_c12_0;
  wire [7:0] t_r13_c12_1;
  wire [7:0] t_r13_c12_2;
  wire [7:0] t_r13_c12_3;
  wire [7:0] t_r13_c12_4;
  wire [7:0] t_r13_c12_5;
  wire [7:0] t_r13_c12_6;
  wire [7:0] t_r13_c12_7;
  wire [7:0] t_r13_c12_8;
  wire [7:0] t_r13_c12_9;
  wire [7:0] t_r13_c12_10;
  wire [7:0] t_r13_c12_11;
  wire [7:0] t_r13_c12_12;
  wire [7:0] t_r13_c13_0;
  wire [7:0] t_r13_c13_1;
  wire [7:0] t_r13_c13_2;
  wire [7:0] t_r13_c13_3;
  wire [7:0] t_r13_c13_4;
  wire [7:0] t_r13_c13_5;
  wire [7:0] t_r13_c13_6;
  wire [7:0] t_r13_c13_7;
  wire [7:0] t_r13_c13_8;
  wire [7:0] t_r13_c13_9;
  wire [7:0] t_r13_c13_10;
  wire [7:0] t_r13_c13_11;
  wire [7:0] t_r13_c13_12;
  wire [7:0] t_r13_c14_0;
  wire [7:0] t_r13_c14_1;
  wire [7:0] t_r13_c14_2;
  wire [7:0] t_r13_c14_3;
  wire [7:0] t_r13_c14_4;
  wire [7:0] t_r13_c14_5;
  wire [7:0] t_r13_c14_6;
  wire [7:0] t_r13_c14_7;
  wire [7:0] t_r13_c14_8;
  wire [7:0] t_r13_c14_9;
  wire [7:0] t_r13_c14_10;
  wire [7:0] t_r13_c14_11;
  wire [7:0] t_r13_c14_12;
  wire [7:0] t_r13_c15_0;
  wire [7:0] t_r13_c15_1;
  wire [7:0] t_r13_c15_2;
  wire [7:0] t_r13_c15_3;
  wire [7:0] t_r13_c15_4;
  wire [7:0] t_r13_c15_5;
  wire [7:0] t_r13_c15_6;
  wire [7:0] t_r13_c15_7;
  wire [7:0] t_r13_c15_8;
  wire [7:0] t_r13_c15_9;
  wire [7:0] t_r13_c15_10;
  wire [7:0] t_r13_c15_11;
  wire [7:0] t_r13_c15_12;
  wire [7:0] t_r13_c16_0;
  wire [7:0] t_r13_c16_1;
  wire [7:0] t_r13_c16_2;
  wire [7:0] t_r13_c16_3;
  wire [7:0] t_r13_c16_4;
  wire [7:0] t_r13_c16_5;
  wire [7:0] t_r13_c16_6;
  wire [7:0] t_r13_c16_7;
  wire [7:0] t_r13_c16_8;
  wire [7:0] t_r13_c16_9;
  wire [7:0] t_r13_c16_10;
  wire [7:0] t_r13_c16_11;
  wire [7:0] t_r13_c16_12;
  wire [7:0] t_r13_c17_0;
  wire [7:0] t_r13_c17_1;
  wire [7:0] t_r13_c17_2;
  wire [7:0] t_r13_c17_3;
  wire [7:0] t_r13_c17_4;
  wire [7:0] t_r13_c17_5;
  wire [7:0] t_r13_c17_6;
  wire [7:0] t_r13_c17_7;
  wire [7:0] t_r13_c17_8;
  wire [7:0] t_r13_c17_9;
  wire [7:0] t_r13_c17_10;
  wire [7:0] t_r13_c17_11;
  wire [7:0] t_r13_c17_12;
  wire [7:0] t_r13_c18_0;
  wire [7:0] t_r13_c18_1;
  wire [7:0] t_r13_c18_2;
  wire [7:0] t_r13_c18_3;
  wire [7:0] t_r13_c18_4;
  wire [7:0] t_r13_c18_5;
  wire [7:0] t_r13_c18_6;
  wire [7:0] t_r13_c18_7;
  wire [7:0] t_r13_c18_8;
  wire [7:0] t_r13_c18_9;
  wire [7:0] t_r13_c18_10;
  wire [7:0] t_r13_c18_11;
  wire [7:0] t_r13_c18_12;
  wire [7:0] t_r13_c19_0;
  wire [7:0] t_r13_c19_1;
  wire [7:0] t_r13_c19_2;
  wire [7:0] t_r13_c19_3;
  wire [7:0] t_r13_c19_4;
  wire [7:0] t_r13_c19_5;
  wire [7:0] t_r13_c19_6;
  wire [7:0] t_r13_c19_7;
  wire [7:0] t_r13_c19_8;
  wire [7:0] t_r13_c19_9;
  wire [7:0] t_r13_c19_10;
  wire [7:0] t_r13_c19_11;
  wire [7:0] t_r13_c19_12;
  wire [7:0] t_r13_c20_0;
  wire [7:0] t_r13_c20_1;
  wire [7:0] t_r13_c20_2;
  wire [7:0] t_r13_c20_3;
  wire [7:0] t_r13_c20_4;
  wire [7:0] t_r13_c20_5;
  wire [7:0] t_r13_c20_6;
  wire [7:0] t_r13_c20_7;
  wire [7:0] t_r13_c20_8;
  wire [7:0] t_r13_c20_9;
  wire [7:0] t_r13_c20_10;
  wire [7:0] t_r13_c20_11;
  wire [7:0] t_r13_c20_12;
  wire [7:0] t_r13_c21_0;
  wire [7:0] t_r13_c21_1;
  wire [7:0] t_r13_c21_2;
  wire [7:0] t_r13_c21_3;
  wire [7:0] t_r13_c21_4;
  wire [7:0] t_r13_c21_5;
  wire [7:0] t_r13_c21_6;
  wire [7:0] t_r13_c21_7;
  wire [7:0] t_r13_c21_8;
  wire [7:0] t_r13_c21_9;
  wire [7:0] t_r13_c21_10;
  wire [7:0] t_r13_c21_11;
  wire [7:0] t_r13_c21_12;
  wire [7:0] t_r13_c22_0;
  wire [7:0] t_r13_c22_1;
  wire [7:0] t_r13_c22_2;
  wire [7:0] t_r13_c22_3;
  wire [7:0] t_r13_c22_4;
  wire [7:0] t_r13_c22_5;
  wire [7:0] t_r13_c22_6;
  wire [7:0] t_r13_c22_7;
  wire [7:0] t_r13_c22_8;
  wire [7:0] t_r13_c22_9;
  wire [7:0] t_r13_c22_10;
  wire [7:0] t_r13_c22_11;
  wire [7:0] t_r13_c22_12;
  wire [7:0] t_r13_c23_0;
  wire [7:0] t_r13_c23_1;
  wire [7:0] t_r13_c23_2;
  wire [7:0] t_r13_c23_3;
  wire [7:0] t_r13_c23_4;
  wire [7:0] t_r13_c23_5;
  wire [7:0] t_r13_c23_6;
  wire [7:0] t_r13_c23_7;
  wire [7:0] t_r13_c23_8;
  wire [7:0] t_r13_c23_9;
  wire [7:0] t_r13_c23_10;
  wire [7:0] t_r13_c23_11;
  wire [7:0] t_r13_c23_12;
  wire [7:0] t_r13_c24_0;
  wire [7:0] t_r13_c24_1;
  wire [7:0] t_r13_c24_2;
  wire [7:0] t_r13_c24_3;
  wire [7:0] t_r13_c24_4;
  wire [7:0] t_r13_c24_5;
  wire [7:0] t_r13_c24_6;
  wire [7:0] t_r13_c24_7;
  wire [7:0] t_r13_c24_8;
  wire [7:0] t_r13_c24_9;
  wire [7:0] t_r13_c24_10;
  wire [7:0] t_r13_c24_11;
  wire [7:0] t_r13_c24_12;
  wire [7:0] t_r13_c25_0;
  wire [7:0] t_r13_c25_1;
  wire [7:0] t_r13_c25_2;
  wire [7:0] t_r13_c25_3;
  wire [7:0] t_r13_c25_4;
  wire [7:0] t_r13_c25_5;
  wire [7:0] t_r13_c25_6;
  wire [7:0] t_r13_c25_7;
  wire [7:0] t_r13_c25_8;
  wire [7:0] t_r13_c25_9;
  wire [7:0] t_r13_c25_10;
  wire [7:0] t_r13_c25_11;
  wire [7:0] t_r13_c25_12;
  wire [7:0] t_r13_c26_0;
  wire [7:0] t_r13_c26_1;
  wire [7:0] t_r13_c26_2;
  wire [7:0] t_r13_c26_3;
  wire [7:0] t_r13_c26_4;
  wire [7:0] t_r13_c26_5;
  wire [7:0] t_r13_c26_6;
  wire [7:0] t_r13_c26_7;
  wire [7:0] t_r13_c26_8;
  wire [7:0] t_r13_c26_9;
  wire [7:0] t_r13_c26_10;
  wire [7:0] t_r13_c26_11;
  wire [7:0] t_r13_c26_12;
  wire [7:0] t_r13_c27_0;
  wire [7:0] t_r13_c27_1;
  wire [7:0] t_r13_c27_2;
  wire [7:0] t_r13_c27_3;
  wire [7:0] t_r13_c27_4;
  wire [7:0] t_r13_c27_5;
  wire [7:0] t_r13_c27_6;
  wire [7:0] t_r13_c27_7;
  wire [7:0] t_r13_c27_8;
  wire [7:0] t_r13_c27_9;
  wire [7:0] t_r13_c27_10;
  wire [7:0] t_r13_c27_11;
  wire [7:0] t_r13_c27_12;
  wire [7:0] t_r13_c28_0;
  wire [7:0] t_r13_c28_1;
  wire [7:0] t_r13_c28_2;
  wire [7:0] t_r13_c28_3;
  wire [7:0] t_r13_c28_4;
  wire [7:0] t_r13_c28_5;
  wire [7:0] t_r13_c28_6;
  wire [7:0] t_r13_c28_7;
  wire [7:0] t_r13_c28_8;
  wire [7:0] t_r13_c28_9;
  wire [7:0] t_r13_c28_10;
  wire [7:0] t_r13_c28_11;
  wire [7:0] t_r13_c28_12;
  wire [7:0] t_r13_c29_0;
  wire [7:0] t_r13_c29_1;
  wire [7:0] t_r13_c29_2;
  wire [7:0] t_r13_c29_3;
  wire [7:0] t_r13_c29_4;
  wire [7:0] t_r13_c29_5;
  wire [7:0] t_r13_c29_6;
  wire [7:0] t_r13_c29_7;
  wire [7:0] t_r13_c29_8;
  wire [7:0] t_r13_c29_9;
  wire [7:0] t_r13_c29_10;
  wire [7:0] t_r13_c29_11;
  wire [7:0] t_r13_c29_12;
  wire [7:0] t_r13_c30_0;
  wire [7:0] t_r13_c30_1;
  wire [7:0] t_r13_c30_2;
  wire [7:0] t_r13_c30_3;
  wire [7:0] t_r13_c30_4;
  wire [7:0] t_r13_c30_5;
  wire [7:0] t_r13_c30_6;
  wire [7:0] t_r13_c30_7;
  wire [7:0] t_r13_c30_8;
  wire [7:0] t_r13_c30_9;
  wire [7:0] t_r13_c30_10;
  wire [7:0] t_r13_c30_11;
  wire [7:0] t_r13_c30_12;
  wire [7:0] t_r13_c31_0;
  wire [7:0] t_r13_c31_1;
  wire [7:0] t_r13_c31_2;
  wire [7:0] t_r13_c31_3;
  wire [7:0] t_r13_c31_4;
  wire [7:0] t_r13_c31_5;
  wire [7:0] t_r13_c31_6;
  wire [7:0] t_r13_c31_7;
  wire [7:0] t_r13_c31_8;
  wire [7:0] t_r13_c31_9;
  wire [7:0] t_r13_c31_10;
  wire [7:0] t_r13_c31_11;
  wire [7:0] t_r13_c31_12;
  wire [7:0] t_r13_c32_0;
  wire [7:0] t_r13_c32_1;
  wire [7:0] t_r13_c32_2;
  wire [7:0] t_r13_c32_3;
  wire [7:0] t_r13_c32_4;
  wire [7:0] t_r13_c32_5;
  wire [7:0] t_r13_c32_6;
  wire [7:0] t_r13_c32_7;
  wire [7:0] t_r13_c32_8;
  wire [7:0] t_r13_c32_9;
  wire [7:0] t_r13_c32_10;
  wire [7:0] t_r13_c32_11;
  wire [7:0] t_r13_c32_12;
  wire [7:0] t_r13_c33_0;
  wire [7:0] t_r13_c33_1;
  wire [7:0] t_r13_c33_2;
  wire [7:0] t_r13_c33_3;
  wire [7:0] t_r13_c33_4;
  wire [7:0] t_r13_c33_5;
  wire [7:0] t_r13_c33_6;
  wire [7:0] t_r13_c33_7;
  wire [7:0] t_r13_c33_8;
  wire [7:0] t_r13_c33_9;
  wire [7:0] t_r13_c33_10;
  wire [7:0] t_r13_c33_11;
  wire [7:0] t_r13_c33_12;
  wire [7:0] t_r13_c34_0;
  wire [7:0] t_r13_c34_1;
  wire [7:0] t_r13_c34_2;
  wire [7:0] t_r13_c34_3;
  wire [7:0] t_r13_c34_4;
  wire [7:0] t_r13_c34_5;
  wire [7:0] t_r13_c34_6;
  wire [7:0] t_r13_c34_7;
  wire [7:0] t_r13_c34_8;
  wire [7:0] t_r13_c34_9;
  wire [7:0] t_r13_c34_10;
  wire [7:0] t_r13_c34_11;
  wire [7:0] t_r13_c34_12;
  wire [7:0] t_r13_c35_0;
  wire [7:0] t_r13_c35_1;
  wire [7:0] t_r13_c35_2;
  wire [7:0] t_r13_c35_3;
  wire [7:0] t_r13_c35_4;
  wire [7:0] t_r13_c35_5;
  wire [7:0] t_r13_c35_6;
  wire [7:0] t_r13_c35_7;
  wire [7:0] t_r13_c35_8;
  wire [7:0] t_r13_c35_9;
  wire [7:0] t_r13_c35_10;
  wire [7:0] t_r13_c35_11;
  wire [7:0] t_r13_c35_12;
  wire [7:0] t_r13_c36_0;
  wire [7:0] t_r13_c36_1;
  wire [7:0] t_r13_c36_2;
  wire [7:0] t_r13_c36_3;
  wire [7:0] t_r13_c36_4;
  wire [7:0] t_r13_c36_5;
  wire [7:0] t_r13_c36_6;
  wire [7:0] t_r13_c36_7;
  wire [7:0] t_r13_c36_8;
  wire [7:0] t_r13_c36_9;
  wire [7:0] t_r13_c36_10;
  wire [7:0] t_r13_c36_11;
  wire [7:0] t_r13_c36_12;
  wire [7:0] t_r13_c37_0;
  wire [7:0] t_r13_c37_1;
  wire [7:0] t_r13_c37_2;
  wire [7:0] t_r13_c37_3;
  wire [7:0] t_r13_c37_4;
  wire [7:0] t_r13_c37_5;
  wire [7:0] t_r13_c37_6;
  wire [7:0] t_r13_c37_7;
  wire [7:0] t_r13_c37_8;
  wire [7:0] t_r13_c37_9;
  wire [7:0] t_r13_c37_10;
  wire [7:0] t_r13_c37_11;
  wire [7:0] t_r13_c37_12;
  wire [7:0] t_r13_c38_0;
  wire [7:0] t_r13_c38_1;
  wire [7:0] t_r13_c38_2;
  wire [7:0] t_r13_c38_3;
  wire [7:0] t_r13_c38_4;
  wire [7:0] t_r13_c38_5;
  wire [7:0] t_r13_c38_6;
  wire [7:0] t_r13_c38_7;
  wire [7:0] t_r13_c38_8;
  wire [7:0] t_r13_c38_9;
  wire [7:0] t_r13_c38_10;
  wire [7:0] t_r13_c38_11;
  wire [7:0] t_r13_c38_12;
  wire [7:0] t_r13_c39_0;
  wire [7:0] t_r13_c39_1;
  wire [7:0] t_r13_c39_2;
  wire [7:0] t_r13_c39_3;
  wire [7:0] t_r13_c39_4;
  wire [7:0] t_r13_c39_5;
  wire [7:0] t_r13_c39_6;
  wire [7:0] t_r13_c39_7;
  wire [7:0] t_r13_c39_8;
  wire [7:0] t_r13_c39_9;
  wire [7:0] t_r13_c39_10;
  wire [7:0] t_r13_c39_11;
  wire [7:0] t_r13_c39_12;
  wire [7:0] t_r13_c40_0;
  wire [7:0] t_r13_c40_1;
  wire [7:0] t_r13_c40_2;
  wire [7:0] t_r13_c40_3;
  wire [7:0] t_r13_c40_4;
  wire [7:0] t_r13_c40_5;
  wire [7:0] t_r13_c40_6;
  wire [7:0] t_r13_c40_7;
  wire [7:0] t_r13_c40_8;
  wire [7:0] t_r13_c40_9;
  wire [7:0] t_r13_c40_10;
  wire [7:0] t_r13_c40_11;
  wire [7:0] t_r13_c40_12;
  wire [7:0] t_r13_c41_0;
  wire [7:0] t_r13_c41_1;
  wire [7:0] t_r13_c41_2;
  wire [7:0] t_r13_c41_3;
  wire [7:0] t_r13_c41_4;
  wire [7:0] t_r13_c41_5;
  wire [7:0] t_r13_c41_6;
  wire [7:0] t_r13_c41_7;
  wire [7:0] t_r13_c41_8;
  wire [7:0] t_r13_c41_9;
  wire [7:0] t_r13_c41_10;
  wire [7:0] t_r13_c41_11;
  wire [7:0] t_r13_c41_12;
  wire [7:0] t_r13_c42_0;
  wire [7:0] t_r13_c42_1;
  wire [7:0] t_r13_c42_2;
  wire [7:0] t_r13_c42_3;
  wire [7:0] t_r13_c42_4;
  wire [7:0] t_r13_c42_5;
  wire [7:0] t_r13_c42_6;
  wire [7:0] t_r13_c42_7;
  wire [7:0] t_r13_c42_8;
  wire [7:0] t_r13_c42_9;
  wire [7:0] t_r13_c42_10;
  wire [7:0] t_r13_c42_11;
  wire [7:0] t_r13_c42_12;
  wire [7:0] t_r13_c43_0;
  wire [7:0] t_r13_c43_1;
  wire [7:0] t_r13_c43_2;
  wire [7:0] t_r13_c43_3;
  wire [7:0] t_r13_c43_4;
  wire [7:0] t_r13_c43_5;
  wire [7:0] t_r13_c43_6;
  wire [7:0] t_r13_c43_7;
  wire [7:0] t_r13_c43_8;
  wire [7:0] t_r13_c43_9;
  wire [7:0] t_r13_c43_10;
  wire [7:0] t_r13_c43_11;
  wire [7:0] t_r13_c43_12;
  wire [7:0] t_r13_c44_0;
  wire [7:0] t_r13_c44_1;
  wire [7:0] t_r13_c44_2;
  wire [7:0] t_r13_c44_3;
  wire [7:0] t_r13_c44_4;
  wire [7:0] t_r13_c44_5;
  wire [7:0] t_r13_c44_6;
  wire [7:0] t_r13_c44_7;
  wire [7:0] t_r13_c44_8;
  wire [7:0] t_r13_c44_9;
  wire [7:0] t_r13_c44_10;
  wire [7:0] t_r13_c44_11;
  wire [7:0] t_r13_c44_12;
  wire [7:0] t_r13_c45_0;
  wire [7:0] t_r13_c45_1;
  wire [7:0] t_r13_c45_2;
  wire [7:0] t_r13_c45_3;
  wire [7:0] t_r13_c45_4;
  wire [7:0] t_r13_c45_5;
  wire [7:0] t_r13_c45_6;
  wire [7:0] t_r13_c45_7;
  wire [7:0] t_r13_c45_8;
  wire [7:0] t_r13_c45_9;
  wire [7:0] t_r13_c45_10;
  wire [7:0] t_r13_c45_11;
  wire [7:0] t_r13_c45_12;
  wire [7:0] t_r13_c46_0;
  wire [7:0] t_r13_c46_1;
  wire [7:0] t_r13_c46_2;
  wire [7:0] t_r13_c46_3;
  wire [7:0] t_r13_c46_4;
  wire [7:0] t_r13_c46_5;
  wire [7:0] t_r13_c46_6;
  wire [7:0] t_r13_c46_7;
  wire [7:0] t_r13_c46_8;
  wire [7:0] t_r13_c46_9;
  wire [7:0] t_r13_c46_10;
  wire [7:0] t_r13_c46_11;
  wire [7:0] t_r13_c46_12;
  wire [7:0] t_r13_c47_0;
  wire [7:0] t_r13_c47_1;
  wire [7:0] t_r13_c47_2;
  wire [7:0] t_r13_c47_3;
  wire [7:0] t_r13_c47_4;
  wire [7:0] t_r13_c47_5;
  wire [7:0] t_r13_c47_6;
  wire [7:0] t_r13_c47_7;
  wire [7:0] t_r13_c47_8;
  wire [7:0] t_r13_c47_9;
  wire [7:0] t_r13_c47_10;
  wire [7:0] t_r13_c47_11;
  wire [7:0] t_r13_c47_12;
  wire [7:0] t_r13_c48_0;
  wire [7:0] t_r13_c48_1;
  wire [7:0] t_r13_c48_2;
  wire [7:0] t_r13_c48_3;
  wire [7:0] t_r13_c48_4;
  wire [7:0] t_r13_c48_5;
  wire [7:0] t_r13_c48_6;
  wire [7:0] t_r13_c48_7;
  wire [7:0] t_r13_c48_8;
  wire [7:0] t_r13_c48_9;
  wire [7:0] t_r13_c48_10;
  wire [7:0] t_r13_c48_11;
  wire [7:0] t_r13_c48_12;
  wire [7:0] t_r13_c49_0;
  wire [7:0] t_r13_c49_1;
  wire [7:0] t_r13_c49_2;
  wire [7:0] t_r13_c49_3;
  wire [7:0] t_r13_c49_4;
  wire [7:0] t_r13_c49_5;
  wire [7:0] t_r13_c49_6;
  wire [7:0] t_r13_c49_7;
  wire [7:0] t_r13_c49_8;
  wire [7:0] t_r13_c49_9;
  wire [7:0] t_r13_c49_10;
  wire [7:0] t_r13_c49_11;
  wire [7:0] t_r13_c49_12;
  wire [7:0] t_r13_c50_0;
  wire [7:0] t_r13_c50_1;
  wire [7:0] t_r13_c50_2;
  wire [7:0] t_r13_c50_3;
  wire [7:0] t_r13_c50_4;
  wire [7:0] t_r13_c50_5;
  wire [7:0] t_r13_c50_6;
  wire [7:0] t_r13_c50_7;
  wire [7:0] t_r13_c50_8;
  wire [7:0] t_r13_c50_9;
  wire [7:0] t_r13_c50_10;
  wire [7:0] t_r13_c50_11;
  wire [7:0] t_r13_c50_12;
  wire [7:0] t_r13_c51_0;
  wire [7:0] t_r13_c51_1;
  wire [7:0] t_r13_c51_2;
  wire [7:0] t_r13_c51_3;
  wire [7:0] t_r13_c51_4;
  wire [7:0] t_r13_c51_5;
  wire [7:0] t_r13_c51_6;
  wire [7:0] t_r13_c51_7;
  wire [7:0] t_r13_c51_8;
  wire [7:0] t_r13_c51_9;
  wire [7:0] t_r13_c51_10;
  wire [7:0] t_r13_c51_11;
  wire [7:0] t_r13_c51_12;
  wire [7:0] t_r13_c52_0;
  wire [7:0] t_r13_c52_1;
  wire [7:0] t_r13_c52_2;
  wire [7:0] t_r13_c52_3;
  wire [7:0] t_r13_c52_4;
  wire [7:0] t_r13_c52_5;
  wire [7:0] t_r13_c52_6;
  wire [7:0] t_r13_c52_7;
  wire [7:0] t_r13_c52_8;
  wire [7:0] t_r13_c52_9;
  wire [7:0] t_r13_c52_10;
  wire [7:0] t_r13_c52_11;
  wire [7:0] t_r13_c52_12;
  wire [7:0] t_r13_c53_0;
  wire [7:0] t_r13_c53_1;
  wire [7:0] t_r13_c53_2;
  wire [7:0] t_r13_c53_3;
  wire [7:0] t_r13_c53_4;
  wire [7:0] t_r13_c53_5;
  wire [7:0] t_r13_c53_6;
  wire [7:0] t_r13_c53_7;
  wire [7:0] t_r13_c53_8;
  wire [7:0] t_r13_c53_9;
  wire [7:0] t_r13_c53_10;
  wire [7:0] t_r13_c53_11;
  wire [7:0] t_r13_c53_12;
  wire [7:0] t_r13_c54_0;
  wire [7:0] t_r13_c54_1;
  wire [7:0] t_r13_c54_2;
  wire [7:0] t_r13_c54_3;
  wire [7:0] t_r13_c54_4;
  wire [7:0] t_r13_c54_5;
  wire [7:0] t_r13_c54_6;
  wire [7:0] t_r13_c54_7;
  wire [7:0] t_r13_c54_8;
  wire [7:0] t_r13_c54_9;
  wire [7:0] t_r13_c54_10;
  wire [7:0] t_r13_c54_11;
  wire [7:0] t_r13_c54_12;
  wire [7:0] t_r13_c55_0;
  wire [7:0] t_r13_c55_1;
  wire [7:0] t_r13_c55_2;
  wire [7:0] t_r13_c55_3;
  wire [7:0] t_r13_c55_4;
  wire [7:0] t_r13_c55_5;
  wire [7:0] t_r13_c55_6;
  wire [7:0] t_r13_c55_7;
  wire [7:0] t_r13_c55_8;
  wire [7:0] t_r13_c55_9;
  wire [7:0] t_r13_c55_10;
  wire [7:0] t_r13_c55_11;
  wire [7:0] t_r13_c55_12;
  wire [7:0] t_r13_c56_0;
  wire [7:0] t_r13_c56_1;
  wire [7:0] t_r13_c56_2;
  wire [7:0] t_r13_c56_3;
  wire [7:0] t_r13_c56_4;
  wire [7:0] t_r13_c56_5;
  wire [7:0] t_r13_c56_6;
  wire [7:0] t_r13_c56_7;
  wire [7:0] t_r13_c56_8;
  wire [7:0] t_r13_c56_9;
  wire [7:0] t_r13_c56_10;
  wire [7:0] t_r13_c56_11;
  wire [7:0] t_r13_c56_12;
  wire [7:0] t_r13_c57_0;
  wire [7:0] t_r13_c57_1;
  wire [7:0] t_r13_c57_2;
  wire [7:0] t_r13_c57_3;
  wire [7:0] t_r13_c57_4;
  wire [7:0] t_r13_c57_5;
  wire [7:0] t_r13_c57_6;
  wire [7:0] t_r13_c57_7;
  wire [7:0] t_r13_c57_8;
  wire [7:0] t_r13_c57_9;
  wire [7:0] t_r13_c57_10;
  wire [7:0] t_r13_c57_11;
  wire [7:0] t_r13_c57_12;
  wire [7:0] t_r13_c58_0;
  wire [7:0] t_r13_c58_1;
  wire [7:0] t_r13_c58_2;
  wire [7:0] t_r13_c58_3;
  wire [7:0] t_r13_c58_4;
  wire [7:0] t_r13_c58_5;
  wire [7:0] t_r13_c58_6;
  wire [7:0] t_r13_c58_7;
  wire [7:0] t_r13_c58_8;
  wire [7:0] t_r13_c58_9;
  wire [7:0] t_r13_c58_10;
  wire [7:0] t_r13_c58_11;
  wire [7:0] t_r13_c58_12;
  wire [7:0] t_r13_c59_0;
  wire [7:0] t_r13_c59_1;
  wire [7:0] t_r13_c59_2;
  wire [7:0] t_r13_c59_3;
  wire [7:0] t_r13_c59_4;
  wire [7:0] t_r13_c59_5;
  wire [7:0] t_r13_c59_6;
  wire [7:0] t_r13_c59_7;
  wire [7:0] t_r13_c59_8;
  wire [7:0] t_r13_c59_9;
  wire [7:0] t_r13_c59_10;
  wire [7:0] t_r13_c59_11;
  wire [7:0] t_r13_c59_12;
  wire [7:0] t_r13_c60_0;
  wire [7:0] t_r13_c60_1;
  wire [7:0] t_r13_c60_2;
  wire [7:0] t_r13_c60_3;
  wire [7:0] t_r13_c60_4;
  wire [7:0] t_r13_c60_5;
  wire [7:0] t_r13_c60_6;
  wire [7:0] t_r13_c60_7;
  wire [7:0] t_r13_c60_8;
  wire [7:0] t_r13_c60_9;
  wire [7:0] t_r13_c60_10;
  wire [7:0] t_r13_c60_11;
  wire [7:0] t_r13_c60_12;
  wire [7:0] t_r13_c61_0;
  wire [7:0] t_r13_c61_1;
  wire [7:0] t_r13_c61_2;
  wire [7:0] t_r13_c61_3;
  wire [7:0] t_r13_c61_4;
  wire [7:0] t_r13_c61_5;
  wire [7:0] t_r13_c61_6;
  wire [7:0] t_r13_c61_7;
  wire [7:0] t_r13_c61_8;
  wire [7:0] t_r13_c61_9;
  wire [7:0] t_r13_c61_10;
  wire [7:0] t_r13_c61_11;
  wire [7:0] t_r13_c61_12;
  wire [7:0] t_r13_c62_0;
  wire [7:0] t_r13_c62_1;
  wire [7:0] t_r13_c62_2;
  wire [7:0] t_r13_c62_3;
  wire [7:0] t_r13_c62_4;
  wire [7:0] t_r13_c62_5;
  wire [7:0] t_r13_c62_6;
  wire [7:0] t_r13_c62_7;
  wire [7:0] t_r13_c62_8;
  wire [7:0] t_r13_c62_9;
  wire [7:0] t_r13_c62_10;
  wire [7:0] t_r13_c62_11;
  wire [7:0] t_r13_c62_12;
  wire [7:0] t_r13_c63_0;
  wire [7:0] t_r13_c63_1;
  wire [7:0] t_r13_c63_2;
  wire [7:0] t_r13_c63_3;
  wire [7:0] t_r13_c63_4;
  wire [7:0] t_r13_c63_5;
  wire [7:0] t_r13_c63_6;
  wire [7:0] t_r13_c63_7;
  wire [7:0] t_r13_c63_8;
  wire [7:0] t_r13_c63_9;
  wire [7:0] t_r13_c63_10;
  wire [7:0] t_r13_c63_11;
  wire [7:0] t_r13_c63_12;
  wire [7:0] t_r13_c64_0;
  wire [7:0] t_r13_c64_1;
  wire [7:0] t_r13_c64_2;
  wire [7:0] t_r13_c64_3;
  wire [7:0] t_r13_c64_4;
  wire [7:0] t_r13_c64_5;
  wire [7:0] t_r13_c64_6;
  wire [7:0] t_r13_c64_7;
  wire [7:0] t_r13_c64_8;
  wire [7:0] t_r13_c64_9;
  wire [7:0] t_r13_c64_10;
  wire [7:0] t_r13_c64_11;
  wire [7:0] t_r13_c64_12;
  wire [7:0] t_r13_c65_0;
  wire [7:0] t_r13_c65_1;
  wire [7:0] t_r13_c65_2;
  wire [7:0] t_r13_c65_3;
  wire [7:0] t_r13_c65_4;
  wire [7:0] t_r13_c65_5;
  wire [7:0] t_r13_c65_6;
  wire [7:0] t_r13_c65_7;
  wire [7:0] t_r13_c65_8;
  wire [7:0] t_r13_c65_9;
  wire [7:0] t_r13_c65_10;
  wire [7:0] t_r13_c65_11;
  wire [7:0] t_r13_c65_12;
  wire [7:0] t_r14_c0_0;
  wire [7:0] t_r14_c0_1;
  wire [7:0] t_r14_c0_2;
  wire [7:0] t_r14_c0_3;
  wire [7:0] t_r14_c0_4;
  wire [7:0] t_r14_c0_5;
  wire [7:0] t_r14_c0_6;
  wire [7:0] t_r14_c0_7;
  wire [7:0] t_r14_c0_8;
  wire [7:0] t_r14_c0_9;
  wire [7:0] t_r14_c0_10;
  wire [7:0] t_r14_c0_11;
  wire [7:0] t_r14_c0_12;
  wire [7:0] t_r14_c1_0;
  wire [7:0] t_r14_c1_1;
  wire [7:0] t_r14_c1_2;
  wire [7:0] t_r14_c1_3;
  wire [7:0] t_r14_c1_4;
  wire [7:0] t_r14_c1_5;
  wire [7:0] t_r14_c1_6;
  wire [7:0] t_r14_c1_7;
  wire [7:0] t_r14_c1_8;
  wire [7:0] t_r14_c1_9;
  wire [7:0] t_r14_c1_10;
  wire [7:0] t_r14_c1_11;
  wire [7:0] t_r14_c1_12;
  wire [7:0] t_r14_c2_0;
  wire [7:0] t_r14_c2_1;
  wire [7:0] t_r14_c2_2;
  wire [7:0] t_r14_c2_3;
  wire [7:0] t_r14_c2_4;
  wire [7:0] t_r14_c2_5;
  wire [7:0] t_r14_c2_6;
  wire [7:0] t_r14_c2_7;
  wire [7:0] t_r14_c2_8;
  wire [7:0] t_r14_c2_9;
  wire [7:0] t_r14_c2_10;
  wire [7:0] t_r14_c2_11;
  wire [7:0] t_r14_c2_12;
  wire [7:0] t_r14_c3_0;
  wire [7:0] t_r14_c3_1;
  wire [7:0] t_r14_c3_2;
  wire [7:0] t_r14_c3_3;
  wire [7:0] t_r14_c3_4;
  wire [7:0] t_r14_c3_5;
  wire [7:0] t_r14_c3_6;
  wire [7:0] t_r14_c3_7;
  wire [7:0] t_r14_c3_8;
  wire [7:0] t_r14_c3_9;
  wire [7:0] t_r14_c3_10;
  wire [7:0] t_r14_c3_11;
  wire [7:0] t_r14_c3_12;
  wire [7:0] t_r14_c4_0;
  wire [7:0] t_r14_c4_1;
  wire [7:0] t_r14_c4_2;
  wire [7:0] t_r14_c4_3;
  wire [7:0] t_r14_c4_4;
  wire [7:0] t_r14_c4_5;
  wire [7:0] t_r14_c4_6;
  wire [7:0] t_r14_c4_7;
  wire [7:0] t_r14_c4_8;
  wire [7:0] t_r14_c4_9;
  wire [7:0] t_r14_c4_10;
  wire [7:0] t_r14_c4_11;
  wire [7:0] t_r14_c4_12;
  wire [7:0] t_r14_c5_0;
  wire [7:0] t_r14_c5_1;
  wire [7:0] t_r14_c5_2;
  wire [7:0] t_r14_c5_3;
  wire [7:0] t_r14_c5_4;
  wire [7:0] t_r14_c5_5;
  wire [7:0] t_r14_c5_6;
  wire [7:0] t_r14_c5_7;
  wire [7:0] t_r14_c5_8;
  wire [7:0] t_r14_c5_9;
  wire [7:0] t_r14_c5_10;
  wire [7:0] t_r14_c5_11;
  wire [7:0] t_r14_c5_12;
  wire [7:0] t_r14_c6_0;
  wire [7:0] t_r14_c6_1;
  wire [7:0] t_r14_c6_2;
  wire [7:0] t_r14_c6_3;
  wire [7:0] t_r14_c6_4;
  wire [7:0] t_r14_c6_5;
  wire [7:0] t_r14_c6_6;
  wire [7:0] t_r14_c6_7;
  wire [7:0] t_r14_c6_8;
  wire [7:0] t_r14_c6_9;
  wire [7:0] t_r14_c6_10;
  wire [7:0] t_r14_c6_11;
  wire [7:0] t_r14_c6_12;
  wire [7:0] t_r14_c7_0;
  wire [7:0] t_r14_c7_1;
  wire [7:0] t_r14_c7_2;
  wire [7:0] t_r14_c7_3;
  wire [7:0] t_r14_c7_4;
  wire [7:0] t_r14_c7_5;
  wire [7:0] t_r14_c7_6;
  wire [7:0] t_r14_c7_7;
  wire [7:0] t_r14_c7_8;
  wire [7:0] t_r14_c7_9;
  wire [7:0] t_r14_c7_10;
  wire [7:0] t_r14_c7_11;
  wire [7:0] t_r14_c7_12;
  wire [7:0] t_r14_c8_0;
  wire [7:0] t_r14_c8_1;
  wire [7:0] t_r14_c8_2;
  wire [7:0] t_r14_c8_3;
  wire [7:0] t_r14_c8_4;
  wire [7:0] t_r14_c8_5;
  wire [7:0] t_r14_c8_6;
  wire [7:0] t_r14_c8_7;
  wire [7:0] t_r14_c8_8;
  wire [7:0] t_r14_c8_9;
  wire [7:0] t_r14_c8_10;
  wire [7:0] t_r14_c8_11;
  wire [7:0] t_r14_c8_12;
  wire [7:0] t_r14_c9_0;
  wire [7:0] t_r14_c9_1;
  wire [7:0] t_r14_c9_2;
  wire [7:0] t_r14_c9_3;
  wire [7:0] t_r14_c9_4;
  wire [7:0] t_r14_c9_5;
  wire [7:0] t_r14_c9_6;
  wire [7:0] t_r14_c9_7;
  wire [7:0] t_r14_c9_8;
  wire [7:0] t_r14_c9_9;
  wire [7:0] t_r14_c9_10;
  wire [7:0] t_r14_c9_11;
  wire [7:0] t_r14_c9_12;
  wire [7:0] t_r14_c10_0;
  wire [7:0] t_r14_c10_1;
  wire [7:0] t_r14_c10_2;
  wire [7:0] t_r14_c10_3;
  wire [7:0] t_r14_c10_4;
  wire [7:0] t_r14_c10_5;
  wire [7:0] t_r14_c10_6;
  wire [7:0] t_r14_c10_7;
  wire [7:0] t_r14_c10_8;
  wire [7:0] t_r14_c10_9;
  wire [7:0] t_r14_c10_10;
  wire [7:0] t_r14_c10_11;
  wire [7:0] t_r14_c10_12;
  wire [7:0] t_r14_c11_0;
  wire [7:0] t_r14_c11_1;
  wire [7:0] t_r14_c11_2;
  wire [7:0] t_r14_c11_3;
  wire [7:0] t_r14_c11_4;
  wire [7:0] t_r14_c11_5;
  wire [7:0] t_r14_c11_6;
  wire [7:0] t_r14_c11_7;
  wire [7:0] t_r14_c11_8;
  wire [7:0] t_r14_c11_9;
  wire [7:0] t_r14_c11_10;
  wire [7:0] t_r14_c11_11;
  wire [7:0] t_r14_c11_12;
  wire [7:0] t_r14_c12_0;
  wire [7:0] t_r14_c12_1;
  wire [7:0] t_r14_c12_2;
  wire [7:0] t_r14_c12_3;
  wire [7:0] t_r14_c12_4;
  wire [7:0] t_r14_c12_5;
  wire [7:0] t_r14_c12_6;
  wire [7:0] t_r14_c12_7;
  wire [7:0] t_r14_c12_8;
  wire [7:0] t_r14_c12_9;
  wire [7:0] t_r14_c12_10;
  wire [7:0] t_r14_c12_11;
  wire [7:0] t_r14_c12_12;
  wire [7:0] t_r14_c13_0;
  wire [7:0] t_r14_c13_1;
  wire [7:0] t_r14_c13_2;
  wire [7:0] t_r14_c13_3;
  wire [7:0] t_r14_c13_4;
  wire [7:0] t_r14_c13_5;
  wire [7:0] t_r14_c13_6;
  wire [7:0] t_r14_c13_7;
  wire [7:0] t_r14_c13_8;
  wire [7:0] t_r14_c13_9;
  wire [7:0] t_r14_c13_10;
  wire [7:0] t_r14_c13_11;
  wire [7:0] t_r14_c13_12;
  wire [7:0] t_r14_c14_0;
  wire [7:0] t_r14_c14_1;
  wire [7:0] t_r14_c14_2;
  wire [7:0] t_r14_c14_3;
  wire [7:0] t_r14_c14_4;
  wire [7:0] t_r14_c14_5;
  wire [7:0] t_r14_c14_6;
  wire [7:0] t_r14_c14_7;
  wire [7:0] t_r14_c14_8;
  wire [7:0] t_r14_c14_9;
  wire [7:0] t_r14_c14_10;
  wire [7:0] t_r14_c14_11;
  wire [7:0] t_r14_c14_12;
  wire [7:0] t_r14_c15_0;
  wire [7:0] t_r14_c15_1;
  wire [7:0] t_r14_c15_2;
  wire [7:0] t_r14_c15_3;
  wire [7:0] t_r14_c15_4;
  wire [7:0] t_r14_c15_5;
  wire [7:0] t_r14_c15_6;
  wire [7:0] t_r14_c15_7;
  wire [7:0] t_r14_c15_8;
  wire [7:0] t_r14_c15_9;
  wire [7:0] t_r14_c15_10;
  wire [7:0] t_r14_c15_11;
  wire [7:0] t_r14_c15_12;
  wire [7:0] t_r14_c16_0;
  wire [7:0] t_r14_c16_1;
  wire [7:0] t_r14_c16_2;
  wire [7:0] t_r14_c16_3;
  wire [7:0] t_r14_c16_4;
  wire [7:0] t_r14_c16_5;
  wire [7:0] t_r14_c16_6;
  wire [7:0] t_r14_c16_7;
  wire [7:0] t_r14_c16_8;
  wire [7:0] t_r14_c16_9;
  wire [7:0] t_r14_c16_10;
  wire [7:0] t_r14_c16_11;
  wire [7:0] t_r14_c16_12;
  wire [7:0] t_r14_c17_0;
  wire [7:0] t_r14_c17_1;
  wire [7:0] t_r14_c17_2;
  wire [7:0] t_r14_c17_3;
  wire [7:0] t_r14_c17_4;
  wire [7:0] t_r14_c17_5;
  wire [7:0] t_r14_c17_6;
  wire [7:0] t_r14_c17_7;
  wire [7:0] t_r14_c17_8;
  wire [7:0] t_r14_c17_9;
  wire [7:0] t_r14_c17_10;
  wire [7:0] t_r14_c17_11;
  wire [7:0] t_r14_c17_12;
  wire [7:0] t_r14_c18_0;
  wire [7:0] t_r14_c18_1;
  wire [7:0] t_r14_c18_2;
  wire [7:0] t_r14_c18_3;
  wire [7:0] t_r14_c18_4;
  wire [7:0] t_r14_c18_5;
  wire [7:0] t_r14_c18_6;
  wire [7:0] t_r14_c18_7;
  wire [7:0] t_r14_c18_8;
  wire [7:0] t_r14_c18_9;
  wire [7:0] t_r14_c18_10;
  wire [7:0] t_r14_c18_11;
  wire [7:0] t_r14_c18_12;
  wire [7:0] t_r14_c19_0;
  wire [7:0] t_r14_c19_1;
  wire [7:0] t_r14_c19_2;
  wire [7:0] t_r14_c19_3;
  wire [7:0] t_r14_c19_4;
  wire [7:0] t_r14_c19_5;
  wire [7:0] t_r14_c19_6;
  wire [7:0] t_r14_c19_7;
  wire [7:0] t_r14_c19_8;
  wire [7:0] t_r14_c19_9;
  wire [7:0] t_r14_c19_10;
  wire [7:0] t_r14_c19_11;
  wire [7:0] t_r14_c19_12;
  wire [7:0] t_r14_c20_0;
  wire [7:0] t_r14_c20_1;
  wire [7:0] t_r14_c20_2;
  wire [7:0] t_r14_c20_3;
  wire [7:0] t_r14_c20_4;
  wire [7:0] t_r14_c20_5;
  wire [7:0] t_r14_c20_6;
  wire [7:0] t_r14_c20_7;
  wire [7:0] t_r14_c20_8;
  wire [7:0] t_r14_c20_9;
  wire [7:0] t_r14_c20_10;
  wire [7:0] t_r14_c20_11;
  wire [7:0] t_r14_c20_12;
  wire [7:0] t_r14_c21_0;
  wire [7:0] t_r14_c21_1;
  wire [7:0] t_r14_c21_2;
  wire [7:0] t_r14_c21_3;
  wire [7:0] t_r14_c21_4;
  wire [7:0] t_r14_c21_5;
  wire [7:0] t_r14_c21_6;
  wire [7:0] t_r14_c21_7;
  wire [7:0] t_r14_c21_8;
  wire [7:0] t_r14_c21_9;
  wire [7:0] t_r14_c21_10;
  wire [7:0] t_r14_c21_11;
  wire [7:0] t_r14_c21_12;
  wire [7:0] t_r14_c22_0;
  wire [7:0] t_r14_c22_1;
  wire [7:0] t_r14_c22_2;
  wire [7:0] t_r14_c22_3;
  wire [7:0] t_r14_c22_4;
  wire [7:0] t_r14_c22_5;
  wire [7:0] t_r14_c22_6;
  wire [7:0] t_r14_c22_7;
  wire [7:0] t_r14_c22_8;
  wire [7:0] t_r14_c22_9;
  wire [7:0] t_r14_c22_10;
  wire [7:0] t_r14_c22_11;
  wire [7:0] t_r14_c22_12;
  wire [7:0] t_r14_c23_0;
  wire [7:0] t_r14_c23_1;
  wire [7:0] t_r14_c23_2;
  wire [7:0] t_r14_c23_3;
  wire [7:0] t_r14_c23_4;
  wire [7:0] t_r14_c23_5;
  wire [7:0] t_r14_c23_6;
  wire [7:0] t_r14_c23_7;
  wire [7:0] t_r14_c23_8;
  wire [7:0] t_r14_c23_9;
  wire [7:0] t_r14_c23_10;
  wire [7:0] t_r14_c23_11;
  wire [7:0] t_r14_c23_12;
  wire [7:0] t_r14_c24_0;
  wire [7:0] t_r14_c24_1;
  wire [7:0] t_r14_c24_2;
  wire [7:0] t_r14_c24_3;
  wire [7:0] t_r14_c24_4;
  wire [7:0] t_r14_c24_5;
  wire [7:0] t_r14_c24_6;
  wire [7:0] t_r14_c24_7;
  wire [7:0] t_r14_c24_8;
  wire [7:0] t_r14_c24_9;
  wire [7:0] t_r14_c24_10;
  wire [7:0] t_r14_c24_11;
  wire [7:0] t_r14_c24_12;
  wire [7:0] t_r14_c25_0;
  wire [7:0] t_r14_c25_1;
  wire [7:0] t_r14_c25_2;
  wire [7:0] t_r14_c25_3;
  wire [7:0] t_r14_c25_4;
  wire [7:0] t_r14_c25_5;
  wire [7:0] t_r14_c25_6;
  wire [7:0] t_r14_c25_7;
  wire [7:0] t_r14_c25_8;
  wire [7:0] t_r14_c25_9;
  wire [7:0] t_r14_c25_10;
  wire [7:0] t_r14_c25_11;
  wire [7:0] t_r14_c25_12;
  wire [7:0] t_r14_c26_0;
  wire [7:0] t_r14_c26_1;
  wire [7:0] t_r14_c26_2;
  wire [7:0] t_r14_c26_3;
  wire [7:0] t_r14_c26_4;
  wire [7:0] t_r14_c26_5;
  wire [7:0] t_r14_c26_6;
  wire [7:0] t_r14_c26_7;
  wire [7:0] t_r14_c26_8;
  wire [7:0] t_r14_c26_9;
  wire [7:0] t_r14_c26_10;
  wire [7:0] t_r14_c26_11;
  wire [7:0] t_r14_c26_12;
  wire [7:0] t_r14_c27_0;
  wire [7:0] t_r14_c27_1;
  wire [7:0] t_r14_c27_2;
  wire [7:0] t_r14_c27_3;
  wire [7:0] t_r14_c27_4;
  wire [7:0] t_r14_c27_5;
  wire [7:0] t_r14_c27_6;
  wire [7:0] t_r14_c27_7;
  wire [7:0] t_r14_c27_8;
  wire [7:0] t_r14_c27_9;
  wire [7:0] t_r14_c27_10;
  wire [7:0] t_r14_c27_11;
  wire [7:0] t_r14_c27_12;
  wire [7:0] t_r14_c28_0;
  wire [7:0] t_r14_c28_1;
  wire [7:0] t_r14_c28_2;
  wire [7:0] t_r14_c28_3;
  wire [7:0] t_r14_c28_4;
  wire [7:0] t_r14_c28_5;
  wire [7:0] t_r14_c28_6;
  wire [7:0] t_r14_c28_7;
  wire [7:0] t_r14_c28_8;
  wire [7:0] t_r14_c28_9;
  wire [7:0] t_r14_c28_10;
  wire [7:0] t_r14_c28_11;
  wire [7:0] t_r14_c28_12;
  wire [7:0] t_r14_c29_0;
  wire [7:0] t_r14_c29_1;
  wire [7:0] t_r14_c29_2;
  wire [7:0] t_r14_c29_3;
  wire [7:0] t_r14_c29_4;
  wire [7:0] t_r14_c29_5;
  wire [7:0] t_r14_c29_6;
  wire [7:0] t_r14_c29_7;
  wire [7:0] t_r14_c29_8;
  wire [7:0] t_r14_c29_9;
  wire [7:0] t_r14_c29_10;
  wire [7:0] t_r14_c29_11;
  wire [7:0] t_r14_c29_12;
  wire [7:0] t_r14_c30_0;
  wire [7:0] t_r14_c30_1;
  wire [7:0] t_r14_c30_2;
  wire [7:0] t_r14_c30_3;
  wire [7:0] t_r14_c30_4;
  wire [7:0] t_r14_c30_5;
  wire [7:0] t_r14_c30_6;
  wire [7:0] t_r14_c30_7;
  wire [7:0] t_r14_c30_8;
  wire [7:0] t_r14_c30_9;
  wire [7:0] t_r14_c30_10;
  wire [7:0] t_r14_c30_11;
  wire [7:0] t_r14_c30_12;
  wire [7:0] t_r14_c31_0;
  wire [7:0] t_r14_c31_1;
  wire [7:0] t_r14_c31_2;
  wire [7:0] t_r14_c31_3;
  wire [7:0] t_r14_c31_4;
  wire [7:0] t_r14_c31_5;
  wire [7:0] t_r14_c31_6;
  wire [7:0] t_r14_c31_7;
  wire [7:0] t_r14_c31_8;
  wire [7:0] t_r14_c31_9;
  wire [7:0] t_r14_c31_10;
  wire [7:0] t_r14_c31_11;
  wire [7:0] t_r14_c31_12;
  wire [7:0] t_r14_c32_0;
  wire [7:0] t_r14_c32_1;
  wire [7:0] t_r14_c32_2;
  wire [7:0] t_r14_c32_3;
  wire [7:0] t_r14_c32_4;
  wire [7:0] t_r14_c32_5;
  wire [7:0] t_r14_c32_6;
  wire [7:0] t_r14_c32_7;
  wire [7:0] t_r14_c32_8;
  wire [7:0] t_r14_c32_9;
  wire [7:0] t_r14_c32_10;
  wire [7:0] t_r14_c32_11;
  wire [7:0] t_r14_c32_12;
  wire [7:0] t_r14_c33_0;
  wire [7:0] t_r14_c33_1;
  wire [7:0] t_r14_c33_2;
  wire [7:0] t_r14_c33_3;
  wire [7:0] t_r14_c33_4;
  wire [7:0] t_r14_c33_5;
  wire [7:0] t_r14_c33_6;
  wire [7:0] t_r14_c33_7;
  wire [7:0] t_r14_c33_8;
  wire [7:0] t_r14_c33_9;
  wire [7:0] t_r14_c33_10;
  wire [7:0] t_r14_c33_11;
  wire [7:0] t_r14_c33_12;
  wire [7:0] t_r14_c34_0;
  wire [7:0] t_r14_c34_1;
  wire [7:0] t_r14_c34_2;
  wire [7:0] t_r14_c34_3;
  wire [7:0] t_r14_c34_4;
  wire [7:0] t_r14_c34_5;
  wire [7:0] t_r14_c34_6;
  wire [7:0] t_r14_c34_7;
  wire [7:0] t_r14_c34_8;
  wire [7:0] t_r14_c34_9;
  wire [7:0] t_r14_c34_10;
  wire [7:0] t_r14_c34_11;
  wire [7:0] t_r14_c34_12;
  wire [7:0] t_r14_c35_0;
  wire [7:0] t_r14_c35_1;
  wire [7:0] t_r14_c35_2;
  wire [7:0] t_r14_c35_3;
  wire [7:0] t_r14_c35_4;
  wire [7:0] t_r14_c35_5;
  wire [7:0] t_r14_c35_6;
  wire [7:0] t_r14_c35_7;
  wire [7:0] t_r14_c35_8;
  wire [7:0] t_r14_c35_9;
  wire [7:0] t_r14_c35_10;
  wire [7:0] t_r14_c35_11;
  wire [7:0] t_r14_c35_12;
  wire [7:0] t_r14_c36_0;
  wire [7:0] t_r14_c36_1;
  wire [7:0] t_r14_c36_2;
  wire [7:0] t_r14_c36_3;
  wire [7:0] t_r14_c36_4;
  wire [7:0] t_r14_c36_5;
  wire [7:0] t_r14_c36_6;
  wire [7:0] t_r14_c36_7;
  wire [7:0] t_r14_c36_8;
  wire [7:0] t_r14_c36_9;
  wire [7:0] t_r14_c36_10;
  wire [7:0] t_r14_c36_11;
  wire [7:0] t_r14_c36_12;
  wire [7:0] t_r14_c37_0;
  wire [7:0] t_r14_c37_1;
  wire [7:0] t_r14_c37_2;
  wire [7:0] t_r14_c37_3;
  wire [7:0] t_r14_c37_4;
  wire [7:0] t_r14_c37_5;
  wire [7:0] t_r14_c37_6;
  wire [7:0] t_r14_c37_7;
  wire [7:0] t_r14_c37_8;
  wire [7:0] t_r14_c37_9;
  wire [7:0] t_r14_c37_10;
  wire [7:0] t_r14_c37_11;
  wire [7:0] t_r14_c37_12;
  wire [7:0] t_r14_c38_0;
  wire [7:0] t_r14_c38_1;
  wire [7:0] t_r14_c38_2;
  wire [7:0] t_r14_c38_3;
  wire [7:0] t_r14_c38_4;
  wire [7:0] t_r14_c38_5;
  wire [7:0] t_r14_c38_6;
  wire [7:0] t_r14_c38_7;
  wire [7:0] t_r14_c38_8;
  wire [7:0] t_r14_c38_9;
  wire [7:0] t_r14_c38_10;
  wire [7:0] t_r14_c38_11;
  wire [7:0] t_r14_c38_12;
  wire [7:0] t_r14_c39_0;
  wire [7:0] t_r14_c39_1;
  wire [7:0] t_r14_c39_2;
  wire [7:0] t_r14_c39_3;
  wire [7:0] t_r14_c39_4;
  wire [7:0] t_r14_c39_5;
  wire [7:0] t_r14_c39_6;
  wire [7:0] t_r14_c39_7;
  wire [7:0] t_r14_c39_8;
  wire [7:0] t_r14_c39_9;
  wire [7:0] t_r14_c39_10;
  wire [7:0] t_r14_c39_11;
  wire [7:0] t_r14_c39_12;
  wire [7:0] t_r14_c40_0;
  wire [7:0] t_r14_c40_1;
  wire [7:0] t_r14_c40_2;
  wire [7:0] t_r14_c40_3;
  wire [7:0] t_r14_c40_4;
  wire [7:0] t_r14_c40_5;
  wire [7:0] t_r14_c40_6;
  wire [7:0] t_r14_c40_7;
  wire [7:0] t_r14_c40_8;
  wire [7:0] t_r14_c40_9;
  wire [7:0] t_r14_c40_10;
  wire [7:0] t_r14_c40_11;
  wire [7:0] t_r14_c40_12;
  wire [7:0] t_r14_c41_0;
  wire [7:0] t_r14_c41_1;
  wire [7:0] t_r14_c41_2;
  wire [7:0] t_r14_c41_3;
  wire [7:0] t_r14_c41_4;
  wire [7:0] t_r14_c41_5;
  wire [7:0] t_r14_c41_6;
  wire [7:0] t_r14_c41_7;
  wire [7:0] t_r14_c41_8;
  wire [7:0] t_r14_c41_9;
  wire [7:0] t_r14_c41_10;
  wire [7:0] t_r14_c41_11;
  wire [7:0] t_r14_c41_12;
  wire [7:0] t_r14_c42_0;
  wire [7:0] t_r14_c42_1;
  wire [7:0] t_r14_c42_2;
  wire [7:0] t_r14_c42_3;
  wire [7:0] t_r14_c42_4;
  wire [7:0] t_r14_c42_5;
  wire [7:0] t_r14_c42_6;
  wire [7:0] t_r14_c42_7;
  wire [7:0] t_r14_c42_8;
  wire [7:0] t_r14_c42_9;
  wire [7:0] t_r14_c42_10;
  wire [7:0] t_r14_c42_11;
  wire [7:0] t_r14_c42_12;
  wire [7:0] t_r14_c43_0;
  wire [7:0] t_r14_c43_1;
  wire [7:0] t_r14_c43_2;
  wire [7:0] t_r14_c43_3;
  wire [7:0] t_r14_c43_4;
  wire [7:0] t_r14_c43_5;
  wire [7:0] t_r14_c43_6;
  wire [7:0] t_r14_c43_7;
  wire [7:0] t_r14_c43_8;
  wire [7:0] t_r14_c43_9;
  wire [7:0] t_r14_c43_10;
  wire [7:0] t_r14_c43_11;
  wire [7:0] t_r14_c43_12;
  wire [7:0] t_r14_c44_0;
  wire [7:0] t_r14_c44_1;
  wire [7:0] t_r14_c44_2;
  wire [7:0] t_r14_c44_3;
  wire [7:0] t_r14_c44_4;
  wire [7:0] t_r14_c44_5;
  wire [7:0] t_r14_c44_6;
  wire [7:0] t_r14_c44_7;
  wire [7:0] t_r14_c44_8;
  wire [7:0] t_r14_c44_9;
  wire [7:0] t_r14_c44_10;
  wire [7:0] t_r14_c44_11;
  wire [7:0] t_r14_c44_12;
  wire [7:0] t_r14_c45_0;
  wire [7:0] t_r14_c45_1;
  wire [7:0] t_r14_c45_2;
  wire [7:0] t_r14_c45_3;
  wire [7:0] t_r14_c45_4;
  wire [7:0] t_r14_c45_5;
  wire [7:0] t_r14_c45_6;
  wire [7:0] t_r14_c45_7;
  wire [7:0] t_r14_c45_8;
  wire [7:0] t_r14_c45_9;
  wire [7:0] t_r14_c45_10;
  wire [7:0] t_r14_c45_11;
  wire [7:0] t_r14_c45_12;
  wire [7:0] t_r14_c46_0;
  wire [7:0] t_r14_c46_1;
  wire [7:0] t_r14_c46_2;
  wire [7:0] t_r14_c46_3;
  wire [7:0] t_r14_c46_4;
  wire [7:0] t_r14_c46_5;
  wire [7:0] t_r14_c46_6;
  wire [7:0] t_r14_c46_7;
  wire [7:0] t_r14_c46_8;
  wire [7:0] t_r14_c46_9;
  wire [7:0] t_r14_c46_10;
  wire [7:0] t_r14_c46_11;
  wire [7:0] t_r14_c46_12;
  wire [7:0] t_r14_c47_0;
  wire [7:0] t_r14_c47_1;
  wire [7:0] t_r14_c47_2;
  wire [7:0] t_r14_c47_3;
  wire [7:0] t_r14_c47_4;
  wire [7:0] t_r14_c47_5;
  wire [7:0] t_r14_c47_6;
  wire [7:0] t_r14_c47_7;
  wire [7:0] t_r14_c47_8;
  wire [7:0] t_r14_c47_9;
  wire [7:0] t_r14_c47_10;
  wire [7:0] t_r14_c47_11;
  wire [7:0] t_r14_c47_12;
  wire [7:0] t_r14_c48_0;
  wire [7:0] t_r14_c48_1;
  wire [7:0] t_r14_c48_2;
  wire [7:0] t_r14_c48_3;
  wire [7:0] t_r14_c48_4;
  wire [7:0] t_r14_c48_5;
  wire [7:0] t_r14_c48_6;
  wire [7:0] t_r14_c48_7;
  wire [7:0] t_r14_c48_8;
  wire [7:0] t_r14_c48_9;
  wire [7:0] t_r14_c48_10;
  wire [7:0] t_r14_c48_11;
  wire [7:0] t_r14_c48_12;
  wire [7:0] t_r14_c49_0;
  wire [7:0] t_r14_c49_1;
  wire [7:0] t_r14_c49_2;
  wire [7:0] t_r14_c49_3;
  wire [7:0] t_r14_c49_4;
  wire [7:0] t_r14_c49_5;
  wire [7:0] t_r14_c49_6;
  wire [7:0] t_r14_c49_7;
  wire [7:0] t_r14_c49_8;
  wire [7:0] t_r14_c49_9;
  wire [7:0] t_r14_c49_10;
  wire [7:0] t_r14_c49_11;
  wire [7:0] t_r14_c49_12;
  wire [7:0] t_r14_c50_0;
  wire [7:0] t_r14_c50_1;
  wire [7:0] t_r14_c50_2;
  wire [7:0] t_r14_c50_3;
  wire [7:0] t_r14_c50_4;
  wire [7:0] t_r14_c50_5;
  wire [7:0] t_r14_c50_6;
  wire [7:0] t_r14_c50_7;
  wire [7:0] t_r14_c50_8;
  wire [7:0] t_r14_c50_9;
  wire [7:0] t_r14_c50_10;
  wire [7:0] t_r14_c50_11;
  wire [7:0] t_r14_c50_12;
  wire [7:0] t_r14_c51_0;
  wire [7:0] t_r14_c51_1;
  wire [7:0] t_r14_c51_2;
  wire [7:0] t_r14_c51_3;
  wire [7:0] t_r14_c51_4;
  wire [7:0] t_r14_c51_5;
  wire [7:0] t_r14_c51_6;
  wire [7:0] t_r14_c51_7;
  wire [7:0] t_r14_c51_8;
  wire [7:0] t_r14_c51_9;
  wire [7:0] t_r14_c51_10;
  wire [7:0] t_r14_c51_11;
  wire [7:0] t_r14_c51_12;
  wire [7:0] t_r14_c52_0;
  wire [7:0] t_r14_c52_1;
  wire [7:0] t_r14_c52_2;
  wire [7:0] t_r14_c52_3;
  wire [7:0] t_r14_c52_4;
  wire [7:0] t_r14_c52_5;
  wire [7:0] t_r14_c52_6;
  wire [7:0] t_r14_c52_7;
  wire [7:0] t_r14_c52_8;
  wire [7:0] t_r14_c52_9;
  wire [7:0] t_r14_c52_10;
  wire [7:0] t_r14_c52_11;
  wire [7:0] t_r14_c52_12;
  wire [7:0] t_r14_c53_0;
  wire [7:0] t_r14_c53_1;
  wire [7:0] t_r14_c53_2;
  wire [7:0] t_r14_c53_3;
  wire [7:0] t_r14_c53_4;
  wire [7:0] t_r14_c53_5;
  wire [7:0] t_r14_c53_6;
  wire [7:0] t_r14_c53_7;
  wire [7:0] t_r14_c53_8;
  wire [7:0] t_r14_c53_9;
  wire [7:0] t_r14_c53_10;
  wire [7:0] t_r14_c53_11;
  wire [7:0] t_r14_c53_12;
  wire [7:0] t_r14_c54_0;
  wire [7:0] t_r14_c54_1;
  wire [7:0] t_r14_c54_2;
  wire [7:0] t_r14_c54_3;
  wire [7:0] t_r14_c54_4;
  wire [7:0] t_r14_c54_5;
  wire [7:0] t_r14_c54_6;
  wire [7:0] t_r14_c54_7;
  wire [7:0] t_r14_c54_8;
  wire [7:0] t_r14_c54_9;
  wire [7:0] t_r14_c54_10;
  wire [7:0] t_r14_c54_11;
  wire [7:0] t_r14_c54_12;
  wire [7:0] t_r14_c55_0;
  wire [7:0] t_r14_c55_1;
  wire [7:0] t_r14_c55_2;
  wire [7:0] t_r14_c55_3;
  wire [7:0] t_r14_c55_4;
  wire [7:0] t_r14_c55_5;
  wire [7:0] t_r14_c55_6;
  wire [7:0] t_r14_c55_7;
  wire [7:0] t_r14_c55_8;
  wire [7:0] t_r14_c55_9;
  wire [7:0] t_r14_c55_10;
  wire [7:0] t_r14_c55_11;
  wire [7:0] t_r14_c55_12;
  wire [7:0] t_r14_c56_0;
  wire [7:0] t_r14_c56_1;
  wire [7:0] t_r14_c56_2;
  wire [7:0] t_r14_c56_3;
  wire [7:0] t_r14_c56_4;
  wire [7:0] t_r14_c56_5;
  wire [7:0] t_r14_c56_6;
  wire [7:0] t_r14_c56_7;
  wire [7:0] t_r14_c56_8;
  wire [7:0] t_r14_c56_9;
  wire [7:0] t_r14_c56_10;
  wire [7:0] t_r14_c56_11;
  wire [7:0] t_r14_c56_12;
  wire [7:0] t_r14_c57_0;
  wire [7:0] t_r14_c57_1;
  wire [7:0] t_r14_c57_2;
  wire [7:0] t_r14_c57_3;
  wire [7:0] t_r14_c57_4;
  wire [7:0] t_r14_c57_5;
  wire [7:0] t_r14_c57_6;
  wire [7:0] t_r14_c57_7;
  wire [7:0] t_r14_c57_8;
  wire [7:0] t_r14_c57_9;
  wire [7:0] t_r14_c57_10;
  wire [7:0] t_r14_c57_11;
  wire [7:0] t_r14_c57_12;
  wire [7:0] t_r14_c58_0;
  wire [7:0] t_r14_c58_1;
  wire [7:0] t_r14_c58_2;
  wire [7:0] t_r14_c58_3;
  wire [7:0] t_r14_c58_4;
  wire [7:0] t_r14_c58_5;
  wire [7:0] t_r14_c58_6;
  wire [7:0] t_r14_c58_7;
  wire [7:0] t_r14_c58_8;
  wire [7:0] t_r14_c58_9;
  wire [7:0] t_r14_c58_10;
  wire [7:0] t_r14_c58_11;
  wire [7:0] t_r14_c58_12;
  wire [7:0] t_r14_c59_0;
  wire [7:0] t_r14_c59_1;
  wire [7:0] t_r14_c59_2;
  wire [7:0] t_r14_c59_3;
  wire [7:0] t_r14_c59_4;
  wire [7:0] t_r14_c59_5;
  wire [7:0] t_r14_c59_6;
  wire [7:0] t_r14_c59_7;
  wire [7:0] t_r14_c59_8;
  wire [7:0] t_r14_c59_9;
  wire [7:0] t_r14_c59_10;
  wire [7:0] t_r14_c59_11;
  wire [7:0] t_r14_c59_12;
  wire [7:0] t_r14_c60_0;
  wire [7:0] t_r14_c60_1;
  wire [7:0] t_r14_c60_2;
  wire [7:0] t_r14_c60_3;
  wire [7:0] t_r14_c60_4;
  wire [7:0] t_r14_c60_5;
  wire [7:0] t_r14_c60_6;
  wire [7:0] t_r14_c60_7;
  wire [7:0] t_r14_c60_8;
  wire [7:0] t_r14_c60_9;
  wire [7:0] t_r14_c60_10;
  wire [7:0] t_r14_c60_11;
  wire [7:0] t_r14_c60_12;
  wire [7:0] t_r14_c61_0;
  wire [7:0] t_r14_c61_1;
  wire [7:0] t_r14_c61_2;
  wire [7:0] t_r14_c61_3;
  wire [7:0] t_r14_c61_4;
  wire [7:0] t_r14_c61_5;
  wire [7:0] t_r14_c61_6;
  wire [7:0] t_r14_c61_7;
  wire [7:0] t_r14_c61_8;
  wire [7:0] t_r14_c61_9;
  wire [7:0] t_r14_c61_10;
  wire [7:0] t_r14_c61_11;
  wire [7:0] t_r14_c61_12;
  wire [7:0] t_r14_c62_0;
  wire [7:0] t_r14_c62_1;
  wire [7:0] t_r14_c62_2;
  wire [7:0] t_r14_c62_3;
  wire [7:0] t_r14_c62_4;
  wire [7:0] t_r14_c62_5;
  wire [7:0] t_r14_c62_6;
  wire [7:0] t_r14_c62_7;
  wire [7:0] t_r14_c62_8;
  wire [7:0] t_r14_c62_9;
  wire [7:0] t_r14_c62_10;
  wire [7:0] t_r14_c62_11;
  wire [7:0] t_r14_c62_12;
  wire [7:0] t_r14_c63_0;
  wire [7:0] t_r14_c63_1;
  wire [7:0] t_r14_c63_2;
  wire [7:0] t_r14_c63_3;
  wire [7:0] t_r14_c63_4;
  wire [7:0] t_r14_c63_5;
  wire [7:0] t_r14_c63_6;
  wire [7:0] t_r14_c63_7;
  wire [7:0] t_r14_c63_8;
  wire [7:0] t_r14_c63_9;
  wire [7:0] t_r14_c63_10;
  wire [7:0] t_r14_c63_11;
  wire [7:0] t_r14_c63_12;
  wire [7:0] t_r14_c64_0;
  wire [7:0] t_r14_c64_1;
  wire [7:0] t_r14_c64_2;
  wire [7:0] t_r14_c64_3;
  wire [7:0] t_r14_c64_4;
  wire [7:0] t_r14_c64_5;
  wire [7:0] t_r14_c64_6;
  wire [7:0] t_r14_c64_7;
  wire [7:0] t_r14_c64_8;
  wire [7:0] t_r14_c64_9;
  wire [7:0] t_r14_c64_10;
  wire [7:0] t_r14_c64_11;
  wire [7:0] t_r14_c64_12;
  wire [7:0] t_r14_c65_0;
  wire [7:0] t_r14_c65_1;
  wire [7:0] t_r14_c65_2;
  wire [7:0] t_r14_c65_3;
  wire [7:0] t_r14_c65_4;
  wire [7:0] t_r14_c65_5;
  wire [7:0] t_r14_c65_6;
  wire [7:0] t_r14_c65_7;
  wire [7:0] t_r14_c65_8;
  wire [7:0] t_r14_c65_9;
  wire [7:0] t_r14_c65_10;
  wire [7:0] t_r14_c65_11;
  wire [7:0] t_r14_c65_12;
  wire [7:0] t_r15_c0_0;
  wire [7:0] t_r15_c0_1;
  wire [7:0] t_r15_c0_2;
  wire [7:0] t_r15_c0_3;
  wire [7:0] t_r15_c0_4;
  wire [7:0] t_r15_c0_5;
  wire [7:0] t_r15_c0_6;
  wire [7:0] t_r15_c0_7;
  wire [7:0] t_r15_c0_8;
  wire [7:0] t_r15_c0_9;
  wire [7:0] t_r15_c0_10;
  wire [7:0] t_r15_c0_11;
  wire [7:0] t_r15_c0_12;
  wire [7:0] t_r15_c1_0;
  wire [7:0] t_r15_c1_1;
  wire [7:0] t_r15_c1_2;
  wire [7:0] t_r15_c1_3;
  wire [7:0] t_r15_c1_4;
  wire [7:0] t_r15_c1_5;
  wire [7:0] t_r15_c1_6;
  wire [7:0] t_r15_c1_7;
  wire [7:0] t_r15_c1_8;
  wire [7:0] t_r15_c1_9;
  wire [7:0] t_r15_c1_10;
  wire [7:0] t_r15_c1_11;
  wire [7:0] t_r15_c1_12;
  wire [7:0] t_r15_c2_0;
  wire [7:0] t_r15_c2_1;
  wire [7:0] t_r15_c2_2;
  wire [7:0] t_r15_c2_3;
  wire [7:0] t_r15_c2_4;
  wire [7:0] t_r15_c2_5;
  wire [7:0] t_r15_c2_6;
  wire [7:0] t_r15_c2_7;
  wire [7:0] t_r15_c2_8;
  wire [7:0] t_r15_c2_9;
  wire [7:0] t_r15_c2_10;
  wire [7:0] t_r15_c2_11;
  wire [7:0] t_r15_c2_12;
  wire [7:0] t_r15_c3_0;
  wire [7:0] t_r15_c3_1;
  wire [7:0] t_r15_c3_2;
  wire [7:0] t_r15_c3_3;
  wire [7:0] t_r15_c3_4;
  wire [7:0] t_r15_c3_5;
  wire [7:0] t_r15_c3_6;
  wire [7:0] t_r15_c3_7;
  wire [7:0] t_r15_c3_8;
  wire [7:0] t_r15_c3_9;
  wire [7:0] t_r15_c3_10;
  wire [7:0] t_r15_c3_11;
  wire [7:0] t_r15_c3_12;
  wire [7:0] t_r15_c4_0;
  wire [7:0] t_r15_c4_1;
  wire [7:0] t_r15_c4_2;
  wire [7:0] t_r15_c4_3;
  wire [7:0] t_r15_c4_4;
  wire [7:0] t_r15_c4_5;
  wire [7:0] t_r15_c4_6;
  wire [7:0] t_r15_c4_7;
  wire [7:0] t_r15_c4_8;
  wire [7:0] t_r15_c4_9;
  wire [7:0] t_r15_c4_10;
  wire [7:0] t_r15_c4_11;
  wire [7:0] t_r15_c4_12;
  wire [7:0] t_r15_c5_0;
  wire [7:0] t_r15_c5_1;
  wire [7:0] t_r15_c5_2;
  wire [7:0] t_r15_c5_3;
  wire [7:0] t_r15_c5_4;
  wire [7:0] t_r15_c5_5;
  wire [7:0] t_r15_c5_6;
  wire [7:0] t_r15_c5_7;
  wire [7:0] t_r15_c5_8;
  wire [7:0] t_r15_c5_9;
  wire [7:0] t_r15_c5_10;
  wire [7:0] t_r15_c5_11;
  wire [7:0] t_r15_c5_12;
  wire [7:0] t_r15_c6_0;
  wire [7:0] t_r15_c6_1;
  wire [7:0] t_r15_c6_2;
  wire [7:0] t_r15_c6_3;
  wire [7:0] t_r15_c6_4;
  wire [7:0] t_r15_c6_5;
  wire [7:0] t_r15_c6_6;
  wire [7:0] t_r15_c6_7;
  wire [7:0] t_r15_c6_8;
  wire [7:0] t_r15_c6_9;
  wire [7:0] t_r15_c6_10;
  wire [7:0] t_r15_c6_11;
  wire [7:0] t_r15_c6_12;
  wire [7:0] t_r15_c7_0;
  wire [7:0] t_r15_c7_1;
  wire [7:0] t_r15_c7_2;
  wire [7:0] t_r15_c7_3;
  wire [7:0] t_r15_c7_4;
  wire [7:0] t_r15_c7_5;
  wire [7:0] t_r15_c7_6;
  wire [7:0] t_r15_c7_7;
  wire [7:0] t_r15_c7_8;
  wire [7:0] t_r15_c7_9;
  wire [7:0] t_r15_c7_10;
  wire [7:0] t_r15_c7_11;
  wire [7:0] t_r15_c7_12;
  wire [7:0] t_r15_c8_0;
  wire [7:0] t_r15_c8_1;
  wire [7:0] t_r15_c8_2;
  wire [7:0] t_r15_c8_3;
  wire [7:0] t_r15_c8_4;
  wire [7:0] t_r15_c8_5;
  wire [7:0] t_r15_c8_6;
  wire [7:0] t_r15_c8_7;
  wire [7:0] t_r15_c8_8;
  wire [7:0] t_r15_c8_9;
  wire [7:0] t_r15_c8_10;
  wire [7:0] t_r15_c8_11;
  wire [7:0] t_r15_c8_12;
  wire [7:0] t_r15_c9_0;
  wire [7:0] t_r15_c9_1;
  wire [7:0] t_r15_c9_2;
  wire [7:0] t_r15_c9_3;
  wire [7:0] t_r15_c9_4;
  wire [7:0] t_r15_c9_5;
  wire [7:0] t_r15_c9_6;
  wire [7:0] t_r15_c9_7;
  wire [7:0] t_r15_c9_8;
  wire [7:0] t_r15_c9_9;
  wire [7:0] t_r15_c9_10;
  wire [7:0] t_r15_c9_11;
  wire [7:0] t_r15_c9_12;
  wire [7:0] t_r15_c10_0;
  wire [7:0] t_r15_c10_1;
  wire [7:0] t_r15_c10_2;
  wire [7:0] t_r15_c10_3;
  wire [7:0] t_r15_c10_4;
  wire [7:0] t_r15_c10_5;
  wire [7:0] t_r15_c10_6;
  wire [7:0] t_r15_c10_7;
  wire [7:0] t_r15_c10_8;
  wire [7:0] t_r15_c10_9;
  wire [7:0] t_r15_c10_10;
  wire [7:0] t_r15_c10_11;
  wire [7:0] t_r15_c10_12;
  wire [7:0] t_r15_c11_0;
  wire [7:0] t_r15_c11_1;
  wire [7:0] t_r15_c11_2;
  wire [7:0] t_r15_c11_3;
  wire [7:0] t_r15_c11_4;
  wire [7:0] t_r15_c11_5;
  wire [7:0] t_r15_c11_6;
  wire [7:0] t_r15_c11_7;
  wire [7:0] t_r15_c11_8;
  wire [7:0] t_r15_c11_9;
  wire [7:0] t_r15_c11_10;
  wire [7:0] t_r15_c11_11;
  wire [7:0] t_r15_c11_12;
  wire [7:0] t_r15_c12_0;
  wire [7:0] t_r15_c12_1;
  wire [7:0] t_r15_c12_2;
  wire [7:0] t_r15_c12_3;
  wire [7:0] t_r15_c12_4;
  wire [7:0] t_r15_c12_5;
  wire [7:0] t_r15_c12_6;
  wire [7:0] t_r15_c12_7;
  wire [7:0] t_r15_c12_8;
  wire [7:0] t_r15_c12_9;
  wire [7:0] t_r15_c12_10;
  wire [7:0] t_r15_c12_11;
  wire [7:0] t_r15_c12_12;
  wire [7:0] t_r15_c13_0;
  wire [7:0] t_r15_c13_1;
  wire [7:0] t_r15_c13_2;
  wire [7:0] t_r15_c13_3;
  wire [7:0] t_r15_c13_4;
  wire [7:0] t_r15_c13_5;
  wire [7:0] t_r15_c13_6;
  wire [7:0] t_r15_c13_7;
  wire [7:0] t_r15_c13_8;
  wire [7:0] t_r15_c13_9;
  wire [7:0] t_r15_c13_10;
  wire [7:0] t_r15_c13_11;
  wire [7:0] t_r15_c13_12;
  wire [7:0] t_r15_c14_0;
  wire [7:0] t_r15_c14_1;
  wire [7:0] t_r15_c14_2;
  wire [7:0] t_r15_c14_3;
  wire [7:0] t_r15_c14_4;
  wire [7:0] t_r15_c14_5;
  wire [7:0] t_r15_c14_6;
  wire [7:0] t_r15_c14_7;
  wire [7:0] t_r15_c14_8;
  wire [7:0] t_r15_c14_9;
  wire [7:0] t_r15_c14_10;
  wire [7:0] t_r15_c14_11;
  wire [7:0] t_r15_c14_12;
  wire [7:0] t_r15_c15_0;
  wire [7:0] t_r15_c15_1;
  wire [7:0] t_r15_c15_2;
  wire [7:0] t_r15_c15_3;
  wire [7:0] t_r15_c15_4;
  wire [7:0] t_r15_c15_5;
  wire [7:0] t_r15_c15_6;
  wire [7:0] t_r15_c15_7;
  wire [7:0] t_r15_c15_8;
  wire [7:0] t_r15_c15_9;
  wire [7:0] t_r15_c15_10;
  wire [7:0] t_r15_c15_11;
  wire [7:0] t_r15_c15_12;
  wire [7:0] t_r15_c16_0;
  wire [7:0] t_r15_c16_1;
  wire [7:0] t_r15_c16_2;
  wire [7:0] t_r15_c16_3;
  wire [7:0] t_r15_c16_4;
  wire [7:0] t_r15_c16_5;
  wire [7:0] t_r15_c16_6;
  wire [7:0] t_r15_c16_7;
  wire [7:0] t_r15_c16_8;
  wire [7:0] t_r15_c16_9;
  wire [7:0] t_r15_c16_10;
  wire [7:0] t_r15_c16_11;
  wire [7:0] t_r15_c16_12;
  wire [7:0] t_r15_c17_0;
  wire [7:0] t_r15_c17_1;
  wire [7:0] t_r15_c17_2;
  wire [7:0] t_r15_c17_3;
  wire [7:0] t_r15_c17_4;
  wire [7:0] t_r15_c17_5;
  wire [7:0] t_r15_c17_6;
  wire [7:0] t_r15_c17_7;
  wire [7:0] t_r15_c17_8;
  wire [7:0] t_r15_c17_9;
  wire [7:0] t_r15_c17_10;
  wire [7:0] t_r15_c17_11;
  wire [7:0] t_r15_c17_12;
  wire [7:0] t_r15_c18_0;
  wire [7:0] t_r15_c18_1;
  wire [7:0] t_r15_c18_2;
  wire [7:0] t_r15_c18_3;
  wire [7:0] t_r15_c18_4;
  wire [7:0] t_r15_c18_5;
  wire [7:0] t_r15_c18_6;
  wire [7:0] t_r15_c18_7;
  wire [7:0] t_r15_c18_8;
  wire [7:0] t_r15_c18_9;
  wire [7:0] t_r15_c18_10;
  wire [7:0] t_r15_c18_11;
  wire [7:0] t_r15_c18_12;
  wire [7:0] t_r15_c19_0;
  wire [7:0] t_r15_c19_1;
  wire [7:0] t_r15_c19_2;
  wire [7:0] t_r15_c19_3;
  wire [7:0] t_r15_c19_4;
  wire [7:0] t_r15_c19_5;
  wire [7:0] t_r15_c19_6;
  wire [7:0] t_r15_c19_7;
  wire [7:0] t_r15_c19_8;
  wire [7:0] t_r15_c19_9;
  wire [7:0] t_r15_c19_10;
  wire [7:0] t_r15_c19_11;
  wire [7:0] t_r15_c19_12;
  wire [7:0] t_r15_c20_0;
  wire [7:0] t_r15_c20_1;
  wire [7:0] t_r15_c20_2;
  wire [7:0] t_r15_c20_3;
  wire [7:0] t_r15_c20_4;
  wire [7:0] t_r15_c20_5;
  wire [7:0] t_r15_c20_6;
  wire [7:0] t_r15_c20_7;
  wire [7:0] t_r15_c20_8;
  wire [7:0] t_r15_c20_9;
  wire [7:0] t_r15_c20_10;
  wire [7:0] t_r15_c20_11;
  wire [7:0] t_r15_c20_12;
  wire [7:0] t_r15_c21_0;
  wire [7:0] t_r15_c21_1;
  wire [7:0] t_r15_c21_2;
  wire [7:0] t_r15_c21_3;
  wire [7:0] t_r15_c21_4;
  wire [7:0] t_r15_c21_5;
  wire [7:0] t_r15_c21_6;
  wire [7:0] t_r15_c21_7;
  wire [7:0] t_r15_c21_8;
  wire [7:0] t_r15_c21_9;
  wire [7:0] t_r15_c21_10;
  wire [7:0] t_r15_c21_11;
  wire [7:0] t_r15_c21_12;
  wire [7:0] t_r15_c22_0;
  wire [7:0] t_r15_c22_1;
  wire [7:0] t_r15_c22_2;
  wire [7:0] t_r15_c22_3;
  wire [7:0] t_r15_c22_4;
  wire [7:0] t_r15_c22_5;
  wire [7:0] t_r15_c22_6;
  wire [7:0] t_r15_c22_7;
  wire [7:0] t_r15_c22_8;
  wire [7:0] t_r15_c22_9;
  wire [7:0] t_r15_c22_10;
  wire [7:0] t_r15_c22_11;
  wire [7:0] t_r15_c22_12;
  wire [7:0] t_r15_c23_0;
  wire [7:0] t_r15_c23_1;
  wire [7:0] t_r15_c23_2;
  wire [7:0] t_r15_c23_3;
  wire [7:0] t_r15_c23_4;
  wire [7:0] t_r15_c23_5;
  wire [7:0] t_r15_c23_6;
  wire [7:0] t_r15_c23_7;
  wire [7:0] t_r15_c23_8;
  wire [7:0] t_r15_c23_9;
  wire [7:0] t_r15_c23_10;
  wire [7:0] t_r15_c23_11;
  wire [7:0] t_r15_c23_12;
  wire [7:0] t_r15_c24_0;
  wire [7:0] t_r15_c24_1;
  wire [7:0] t_r15_c24_2;
  wire [7:0] t_r15_c24_3;
  wire [7:0] t_r15_c24_4;
  wire [7:0] t_r15_c24_5;
  wire [7:0] t_r15_c24_6;
  wire [7:0] t_r15_c24_7;
  wire [7:0] t_r15_c24_8;
  wire [7:0] t_r15_c24_9;
  wire [7:0] t_r15_c24_10;
  wire [7:0] t_r15_c24_11;
  wire [7:0] t_r15_c24_12;
  wire [7:0] t_r15_c25_0;
  wire [7:0] t_r15_c25_1;
  wire [7:0] t_r15_c25_2;
  wire [7:0] t_r15_c25_3;
  wire [7:0] t_r15_c25_4;
  wire [7:0] t_r15_c25_5;
  wire [7:0] t_r15_c25_6;
  wire [7:0] t_r15_c25_7;
  wire [7:0] t_r15_c25_8;
  wire [7:0] t_r15_c25_9;
  wire [7:0] t_r15_c25_10;
  wire [7:0] t_r15_c25_11;
  wire [7:0] t_r15_c25_12;
  wire [7:0] t_r15_c26_0;
  wire [7:0] t_r15_c26_1;
  wire [7:0] t_r15_c26_2;
  wire [7:0] t_r15_c26_3;
  wire [7:0] t_r15_c26_4;
  wire [7:0] t_r15_c26_5;
  wire [7:0] t_r15_c26_6;
  wire [7:0] t_r15_c26_7;
  wire [7:0] t_r15_c26_8;
  wire [7:0] t_r15_c26_9;
  wire [7:0] t_r15_c26_10;
  wire [7:0] t_r15_c26_11;
  wire [7:0] t_r15_c26_12;
  wire [7:0] t_r15_c27_0;
  wire [7:0] t_r15_c27_1;
  wire [7:0] t_r15_c27_2;
  wire [7:0] t_r15_c27_3;
  wire [7:0] t_r15_c27_4;
  wire [7:0] t_r15_c27_5;
  wire [7:0] t_r15_c27_6;
  wire [7:0] t_r15_c27_7;
  wire [7:0] t_r15_c27_8;
  wire [7:0] t_r15_c27_9;
  wire [7:0] t_r15_c27_10;
  wire [7:0] t_r15_c27_11;
  wire [7:0] t_r15_c27_12;
  wire [7:0] t_r15_c28_0;
  wire [7:0] t_r15_c28_1;
  wire [7:0] t_r15_c28_2;
  wire [7:0] t_r15_c28_3;
  wire [7:0] t_r15_c28_4;
  wire [7:0] t_r15_c28_5;
  wire [7:0] t_r15_c28_6;
  wire [7:0] t_r15_c28_7;
  wire [7:0] t_r15_c28_8;
  wire [7:0] t_r15_c28_9;
  wire [7:0] t_r15_c28_10;
  wire [7:0] t_r15_c28_11;
  wire [7:0] t_r15_c28_12;
  wire [7:0] t_r15_c29_0;
  wire [7:0] t_r15_c29_1;
  wire [7:0] t_r15_c29_2;
  wire [7:0] t_r15_c29_3;
  wire [7:0] t_r15_c29_4;
  wire [7:0] t_r15_c29_5;
  wire [7:0] t_r15_c29_6;
  wire [7:0] t_r15_c29_7;
  wire [7:0] t_r15_c29_8;
  wire [7:0] t_r15_c29_9;
  wire [7:0] t_r15_c29_10;
  wire [7:0] t_r15_c29_11;
  wire [7:0] t_r15_c29_12;
  wire [7:0] t_r15_c30_0;
  wire [7:0] t_r15_c30_1;
  wire [7:0] t_r15_c30_2;
  wire [7:0] t_r15_c30_3;
  wire [7:0] t_r15_c30_4;
  wire [7:0] t_r15_c30_5;
  wire [7:0] t_r15_c30_6;
  wire [7:0] t_r15_c30_7;
  wire [7:0] t_r15_c30_8;
  wire [7:0] t_r15_c30_9;
  wire [7:0] t_r15_c30_10;
  wire [7:0] t_r15_c30_11;
  wire [7:0] t_r15_c30_12;
  wire [7:0] t_r15_c31_0;
  wire [7:0] t_r15_c31_1;
  wire [7:0] t_r15_c31_2;
  wire [7:0] t_r15_c31_3;
  wire [7:0] t_r15_c31_4;
  wire [7:0] t_r15_c31_5;
  wire [7:0] t_r15_c31_6;
  wire [7:0] t_r15_c31_7;
  wire [7:0] t_r15_c31_8;
  wire [7:0] t_r15_c31_9;
  wire [7:0] t_r15_c31_10;
  wire [7:0] t_r15_c31_11;
  wire [7:0] t_r15_c31_12;
  wire [7:0] t_r15_c32_0;
  wire [7:0] t_r15_c32_1;
  wire [7:0] t_r15_c32_2;
  wire [7:0] t_r15_c32_3;
  wire [7:0] t_r15_c32_4;
  wire [7:0] t_r15_c32_5;
  wire [7:0] t_r15_c32_6;
  wire [7:0] t_r15_c32_7;
  wire [7:0] t_r15_c32_8;
  wire [7:0] t_r15_c32_9;
  wire [7:0] t_r15_c32_10;
  wire [7:0] t_r15_c32_11;
  wire [7:0] t_r15_c32_12;
  wire [7:0] t_r15_c33_0;
  wire [7:0] t_r15_c33_1;
  wire [7:0] t_r15_c33_2;
  wire [7:0] t_r15_c33_3;
  wire [7:0] t_r15_c33_4;
  wire [7:0] t_r15_c33_5;
  wire [7:0] t_r15_c33_6;
  wire [7:0] t_r15_c33_7;
  wire [7:0] t_r15_c33_8;
  wire [7:0] t_r15_c33_9;
  wire [7:0] t_r15_c33_10;
  wire [7:0] t_r15_c33_11;
  wire [7:0] t_r15_c33_12;
  wire [7:0] t_r15_c34_0;
  wire [7:0] t_r15_c34_1;
  wire [7:0] t_r15_c34_2;
  wire [7:0] t_r15_c34_3;
  wire [7:0] t_r15_c34_4;
  wire [7:0] t_r15_c34_5;
  wire [7:0] t_r15_c34_6;
  wire [7:0] t_r15_c34_7;
  wire [7:0] t_r15_c34_8;
  wire [7:0] t_r15_c34_9;
  wire [7:0] t_r15_c34_10;
  wire [7:0] t_r15_c34_11;
  wire [7:0] t_r15_c34_12;
  wire [7:0] t_r15_c35_0;
  wire [7:0] t_r15_c35_1;
  wire [7:0] t_r15_c35_2;
  wire [7:0] t_r15_c35_3;
  wire [7:0] t_r15_c35_4;
  wire [7:0] t_r15_c35_5;
  wire [7:0] t_r15_c35_6;
  wire [7:0] t_r15_c35_7;
  wire [7:0] t_r15_c35_8;
  wire [7:0] t_r15_c35_9;
  wire [7:0] t_r15_c35_10;
  wire [7:0] t_r15_c35_11;
  wire [7:0] t_r15_c35_12;
  wire [7:0] t_r15_c36_0;
  wire [7:0] t_r15_c36_1;
  wire [7:0] t_r15_c36_2;
  wire [7:0] t_r15_c36_3;
  wire [7:0] t_r15_c36_4;
  wire [7:0] t_r15_c36_5;
  wire [7:0] t_r15_c36_6;
  wire [7:0] t_r15_c36_7;
  wire [7:0] t_r15_c36_8;
  wire [7:0] t_r15_c36_9;
  wire [7:0] t_r15_c36_10;
  wire [7:0] t_r15_c36_11;
  wire [7:0] t_r15_c36_12;
  wire [7:0] t_r15_c37_0;
  wire [7:0] t_r15_c37_1;
  wire [7:0] t_r15_c37_2;
  wire [7:0] t_r15_c37_3;
  wire [7:0] t_r15_c37_4;
  wire [7:0] t_r15_c37_5;
  wire [7:0] t_r15_c37_6;
  wire [7:0] t_r15_c37_7;
  wire [7:0] t_r15_c37_8;
  wire [7:0] t_r15_c37_9;
  wire [7:0] t_r15_c37_10;
  wire [7:0] t_r15_c37_11;
  wire [7:0] t_r15_c37_12;
  wire [7:0] t_r15_c38_0;
  wire [7:0] t_r15_c38_1;
  wire [7:0] t_r15_c38_2;
  wire [7:0] t_r15_c38_3;
  wire [7:0] t_r15_c38_4;
  wire [7:0] t_r15_c38_5;
  wire [7:0] t_r15_c38_6;
  wire [7:0] t_r15_c38_7;
  wire [7:0] t_r15_c38_8;
  wire [7:0] t_r15_c38_9;
  wire [7:0] t_r15_c38_10;
  wire [7:0] t_r15_c38_11;
  wire [7:0] t_r15_c38_12;
  wire [7:0] t_r15_c39_0;
  wire [7:0] t_r15_c39_1;
  wire [7:0] t_r15_c39_2;
  wire [7:0] t_r15_c39_3;
  wire [7:0] t_r15_c39_4;
  wire [7:0] t_r15_c39_5;
  wire [7:0] t_r15_c39_6;
  wire [7:0] t_r15_c39_7;
  wire [7:0] t_r15_c39_8;
  wire [7:0] t_r15_c39_9;
  wire [7:0] t_r15_c39_10;
  wire [7:0] t_r15_c39_11;
  wire [7:0] t_r15_c39_12;
  wire [7:0] t_r15_c40_0;
  wire [7:0] t_r15_c40_1;
  wire [7:0] t_r15_c40_2;
  wire [7:0] t_r15_c40_3;
  wire [7:0] t_r15_c40_4;
  wire [7:0] t_r15_c40_5;
  wire [7:0] t_r15_c40_6;
  wire [7:0] t_r15_c40_7;
  wire [7:0] t_r15_c40_8;
  wire [7:0] t_r15_c40_9;
  wire [7:0] t_r15_c40_10;
  wire [7:0] t_r15_c40_11;
  wire [7:0] t_r15_c40_12;
  wire [7:0] t_r15_c41_0;
  wire [7:0] t_r15_c41_1;
  wire [7:0] t_r15_c41_2;
  wire [7:0] t_r15_c41_3;
  wire [7:0] t_r15_c41_4;
  wire [7:0] t_r15_c41_5;
  wire [7:0] t_r15_c41_6;
  wire [7:0] t_r15_c41_7;
  wire [7:0] t_r15_c41_8;
  wire [7:0] t_r15_c41_9;
  wire [7:0] t_r15_c41_10;
  wire [7:0] t_r15_c41_11;
  wire [7:0] t_r15_c41_12;
  wire [7:0] t_r15_c42_0;
  wire [7:0] t_r15_c42_1;
  wire [7:0] t_r15_c42_2;
  wire [7:0] t_r15_c42_3;
  wire [7:0] t_r15_c42_4;
  wire [7:0] t_r15_c42_5;
  wire [7:0] t_r15_c42_6;
  wire [7:0] t_r15_c42_7;
  wire [7:0] t_r15_c42_8;
  wire [7:0] t_r15_c42_9;
  wire [7:0] t_r15_c42_10;
  wire [7:0] t_r15_c42_11;
  wire [7:0] t_r15_c42_12;
  wire [7:0] t_r15_c43_0;
  wire [7:0] t_r15_c43_1;
  wire [7:0] t_r15_c43_2;
  wire [7:0] t_r15_c43_3;
  wire [7:0] t_r15_c43_4;
  wire [7:0] t_r15_c43_5;
  wire [7:0] t_r15_c43_6;
  wire [7:0] t_r15_c43_7;
  wire [7:0] t_r15_c43_8;
  wire [7:0] t_r15_c43_9;
  wire [7:0] t_r15_c43_10;
  wire [7:0] t_r15_c43_11;
  wire [7:0] t_r15_c43_12;
  wire [7:0] t_r15_c44_0;
  wire [7:0] t_r15_c44_1;
  wire [7:0] t_r15_c44_2;
  wire [7:0] t_r15_c44_3;
  wire [7:0] t_r15_c44_4;
  wire [7:0] t_r15_c44_5;
  wire [7:0] t_r15_c44_6;
  wire [7:0] t_r15_c44_7;
  wire [7:0] t_r15_c44_8;
  wire [7:0] t_r15_c44_9;
  wire [7:0] t_r15_c44_10;
  wire [7:0] t_r15_c44_11;
  wire [7:0] t_r15_c44_12;
  wire [7:0] t_r15_c45_0;
  wire [7:0] t_r15_c45_1;
  wire [7:0] t_r15_c45_2;
  wire [7:0] t_r15_c45_3;
  wire [7:0] t_r15_c45_4;
  wire [7:0] t_r15_c45_5;
  wire [7:0] t_r15_c45_6;
  wire [7:0] t_r15_c45_7;
  wire [7:0] t_r15_c45_8;
  wire [7:0] t_r15_c45_9;
  wire [7:0] t_r15_c45_10;
  wire [7:0] t_r15_c45_11;
  wire [7:0] t_r15_c45_12;
  wire [7:0] t_r15_c46_0;
  wire [7:0] t_r15_c46_1;
  wire [7:0] t_r15_c46_2;
  wire [7:0] t_r15_c46_3;
  wire [7:0] t_r15_c46_4;
  wire [7:0] t_r15_c46_5;
  wire [7:0] t_r15_c46_6;
  wire [7:0] t_r15_c46_7;
  wire [7:0] t_r15_c46_8;
  wire [7:0] t_r15_c46_9;
  wire [7:0] t_r15_c46_10;
  wire [7:0] t_r15_c46_11;
  wire [7:0] t_r15_c46_12;
  wire [7:0] t_r15_c47_0;
  wire [7:0] t_r15_c47_1;
  wire [7:0] t_r15_c47_2;
  wire [7:0] t_r15_c47_3;
  wire [7:0] t_r15_c47_4;
  wire [7:0] t_r15_c47_5;
  wire [7:0] t_r15_c47_6;
  wire [7:0] t_r15_c47_7;
  wire [7:0] t_r15_c47_8;
  wire [7:0] t_r15_c47_9;
  wire [7:0] t_r15_c47_10;
  wire [7:0] t_r15_c47_11;
  wire [7:0] t_r15_c47_12;
  wire [7:0] t_r15_c48_0;
  wire [7:0] t_r15_c48_1;
  wire [7:0] t_r15_c48_2;
  wire [7:0] t_r15_c48_3;
  wire [7:0] t_r15_c48_4;
  wire [7:0] t_r15_c48_5;
  wire [7:0] t_r15_c48_6;
  wire [7:0] t_r15_c48_7;
  wire [7:0] t_r15_c48_8;
  wire [7:0] t_r15_c48_9;
  wire [7:0] t_r15_c48_10;
  wire [7:0] t_r15_c48_11;
  wire [7:0] t_r15_c48_12;
  wire [7:0] t_r15_c49_0;
  wire [7:0] t_r15_c49_1;
  wire [7:0] t_r15_c49_2;
  wire [7:0] t_r15_c49_3;
  wire [7:0] t_r15_c49_4;
  wire [7:0] t_r15_c49_5;
  wire [7:0] t_r15_c49_6;
  wire [7:0] t_r15_c49_7;
  wire [7:0] t_r15_c49_8;
  wire [7:0] t_r15_c49_9;
  wire [7:0] t_r15_c49_10;
  wire [7:0] t_r15_c49_11;
  wire [7:0] t_r15_c49_12;
  wire [7:0] t_r15_c50_0;
  wire [7:0] t_r15_c50_1;
  wire [7:0] t_r15_c50_2;
  wire [7:0] t_r15_c50_3;
  wire [7:0] t_r15_c50_4;
  wire [7:0] t_r15_c50_5;
  wire [7:0] t_r15_c50_6;
  wire [7:0] t_r15_c50_7;
  wire [7:0] t_r15_c50_8;
  wire [7:0] t_r15_c50_9;
  wire [7:0] t_r15_c50_10;
  wire [7:0] t_r15_c50_11;
  wire [7:0] t_r15_c50_12;
  wire [7:0] t_r15_c51_0;
  wire [7:0] t_r15_c51_1;
  wire [7:0] t_r15_c51_2;
  wire [7:0] t_r15_c51_3;
  wire [7:0] t_r15_c51_4;
  wire [7:0] t_r15_c51_5;
  wire [7:0] t_r15_c51_6;
  wire [7:0] t_r15_c51_7;
  wire [7:0] t_r15_c51_8;
  wire [7:0] t_r15_c51_9;
  wire [7:0] t_r15_c51_10;
  wire [7:0] t_r15_c51_11;
  wire [7:0] t_r15_c51_12;
  wire [7:0] t_r15_c52_0;
  wire [7:0] t_r15_c52_1;
  wire [7:0] t_r15_c52_2;
  wire [7:0] t_r15_c52_3;
  wire [7:0] t_r15_c52_4;
  wire [7:0] t_r15_c52_5;
  wire [7:0] t_r15_c52_6;
  wire [7:0] t_r15_c52_7;
  wire [7:0] t_r15_c52_8;
  wire [7:0] t_r15_c52_9;
  wire [7:0] t_r15_c52_10;
  wire [7:0] t_r15_c52_11;
  wire [7:0] t_r15_c52_12;
  wire [7:0] t_r15_c53_0;
  wire [7:0] t_r15_c53_1;
  wire [7:0] t_r15_c53_2;
  wire [7:0] t_r15_c53_3;
  wire [7:0] t_r15_c53_4;
  wire [7:0] t_r15_c53_5;
  wire [7:0] t_r15_c53_6;
  wire [7:0] t_r15_c53_7;
  wire [7:0] t_r15_c53_8;
  wire [7:0] t_r15_c53_9;
  wire [7:0] t_r15_c53_10;
  wire [7:0] t_r15_c53_11;
  wire [7:0] t_r15_c53_12;
  wire [7:0] t_r15_c54_0;
  wire [7:0] t_r15_c54_1;
  wire [7:0] t_r15_c54_2;
  wire [7:0] t_r15_c54_3;
  wire [7:0] t_r15_c54_4;
  wire [7:0] t_r15_c54_5;
  wire [7:0] t_r15_c54_6;
  wire [7:0] t_r15_c54_7;
  wire [7:0] t_r15_c54_8;
  wire [7:0] t_r15_c54_9;
  wire [7:0] t_r15_c54_10;
  wire [7:0] t_r15_c54_11;
  wire [7:0] t_r15_c54_12;
  wire [7:0] t_r15_c55_0;
  wire [7:0] t_r15_c55_1;
  wire [7:0] t_r15_c55_2;
  wire [7:0] t_r15_c55_3;
  wire [7:0] t_r15_c55_4;
  wire [7:0] t_r15_c55_5;
  wire [7:0] t_r15_c55_6;
  wire [7:0] t_r15_c55_7;
  wire [7:0] t_r15_c55_8;
  wire [7:0] t_r15_c55_9;
  wire [7:0] t_r15_c55_10;
  wire [7:0] t_r15_c55_11;
  wire [7:0] t_r15_c55_12;
  wire [7:0] t_r15_c56_0;
  wire [7:0] t_r15_c56_1;
  wire [7:0] t_r15_c56_2;
  wire [7:0] t_r15_c56_3;
  wire [7:0] t_r15_c56_4;
  wire [7:0] t_r15_c56_5;
  wire [7:0] t_r15_c56_6;
  wire [7:0] t_r15_c56_7;
  wire [7:0] t_r15_c56_8;
  wire [7:0] t_r15_c56_9;
  wire [7:0] t_r15_c56_10;
  wire [7:0] t_r15_c56_11;
  wire [7:0] t_r15_c56_12;
  wire [7:0] t_r15_c57_0;
  wire [7:0] t_r15_c57_1;
  wire [7:0] t_r15_c57_2;
  wire [7:0] t_r15_c57_3;
  wire [7:0] t_r15_c57_4;
  wire [7:0] t_r15_c57_5;
  wire [7:0] t_r15_c57_6;
  wire [7:0] t_r15_c57_7;
  wire [7:0] t_r15_c57_8;
  wire [7:0] t_r15_c57_9;
  wire [7:0] t_r15_c57_10;
  wire [7:0] t_r15_c57_11;
  wire [7:0] t_r15_c57_12;
  wire [7:0] t_r15_c58_0;
  wire [7:0] t_r15_c58_1;
  wire [7:0] t_r15_c58_2;
  wire [7:0] t_r15_c58_3;
  wire [7:0] t_r15_c58_4;
  wire [7:0] t_r15_c58_5;
  wire [7:0] t_r15_c58_6;
  wire [7:0] t_r15_c58_7;
  wire [7:0] t_r15_c58_8;
  wire [7:0] t_r15_c58_9;
  wire [7:0] t_r15_c58_10;
  wire [7:0] t_r15_c58_11;
  wire [7:0] t_r15_c58_12;
  wire [7:0] t_r15_c59_0;
  wire [7:0] t_r15_c59_1;
  wire [7:0] t_r15_c59_2;
  wire [7:0] t_r15_c59_3;
  wire [7:0] t_r15_c59_4;
  wire [7:0] t_r15_c59_5;
  wire [7:0] t_r15_c59_6;
  wire [7:0] t_r15_c59_7;
  wire [7:0] t_r15_c59_8;
  wire [7:0] t_r15_c59_9;
  wire [7:0] t_r15_c59_10;
  wire [7:0] t_r15_c59_11;
  wire [7:0] t_r15_c59_12;
  wire [7:0] t_r15_c60_0;
  wire [7:0] t_r15_c60_1;
  wire [7:0] t_r15_c60_2;
  wire [7:0] t_r15_c60_3;
  wire [7:0] t_r15_c60_4;
  wire [7:0] t_r15_c60_5;
  wire [7:0] t_r15_c60_6;
  wire [7:0] t_r15_c60_7;
  wire [7:0] t_r15_c60_8;
  wire [7:0] t_r15_c60_9;
  wire [7:0] t_r15_c60_10;
  wire [7:0] t_r15_c60_11;
  wire [7:0] t_r15_c60_12;
  wire [7:0] t_r15_c61_0;
  wire [7:0] t_r15_c61_1;
  wire [7:0] t_r15_c61_2;
  wire [7:0] t_r15_c61_3;
  wire [7:0] t_r15_c61_4;
  wire [7:0] t_r15_c61_5;
  wire [7:0] t_r15_c61_6;
  wire [7:0] t_r15_c61_7;
  wire [7:0] t_r15_c61_8;
  wire [7:0] t_r15_c61_9;
  wire [7:0] t_r15_c61_10;
  wire [7:0] t_r15_c61_11;
  wire [7:0] t_r15_c61_12;
  wire [7:0] t_r15_c62_0;
  wire [7:0] t_r15_c62_1;
  wire [7:0] t_r15_c62_2;
  wire [7:0] t_r15_c62_3;
  wire [7:0] t_r15_c62_4;
  wire [7:0] t_r15_c62_5;
  wire [7:0] t_r15_c62_6;
  wire [7:0] t_r15_c62_7;
  wire [7:0] t_r15_c62_8;
  wire [7:0] t_r15_c62_9;
  wire [7:0] t_r15_c62_10;
  wire [7:0] t_r15_c62_11;
  wire [7:0] t_r15_c62_12;
  wire [7:0] t_r15_c63_0;
  wire [7:0] t_r15_c63_1;
  wire [7:0] t_r15_c63_2;
  wire [7:0] t_r15_c63_3;
  wire [7:0] t_r15_c63_4;
  wire [7:0] t_r15_c63_5;
  wire [7:0] t_r15_c63_6;
  wire [7:0] t_r15_c63_7;
  wire [7:0] t_r15_c63_8;
  wire [7:0] t_r15_c63_9;
  wire [7:0] t_r15_c63_10;
  wire [7:0] t_r15_c63_11;
  wire [7:0] t_r15_c63_12;
  wire [7:0] t_r15_c64_0;
  wire [7:0] t_r15_c64_1;
  wire [7:0] t_r15_c64_2;
  wire [7:0] t_r15_c64_3;
  wire [7:0] t_r15_c64_4;
  wire [7:0] t_r15_c64_5;
  wire [7:0] t_r15_c64_6;
  wire [7:0] t_r15_c64_7;
  wire [7:0] t_r15_c64_8;
  wire [7:0] t_r15_c64_9;
  wire [7:0] t_r15_c64_10;
  wire [7:0] t_r15_c64_11;
  wire [7:0] t_r15_c64_12;
  wire [7:0] t_r15_c65_0;
  wire [7:0] t_r15_c65_1;
  wire [7:0] t_r15_c65_2;
  wire [7:0] t_r15_c65_3;
  wire [7:0] t_r15_c65_4;
  wire [7:0] t_r15_c65_5;
  wire [7:0] t_r15_c65_6;
  wire [7:0] t_r15_c65_7;
  wire [7:0] t_r15_c65_8;
  wire [7:0] t_r15_c65_9;
  wire [7:0] t_r15_c65_10;
  wire [7:0] t_r15_c65_11;
  wire [7:0] t_r15_c65_12;
  wire [7:0] t_r16_c0_0;
  wire [7:0] t_r16_c0_1;
  wire [7:0] t_r16_c0_2;
  wire [7:0] t_r16_c0_3;
  wire [7:0] t_r16_c0_4;
  wire [7:0] t_r16_c0_5;
  wire [7:0] t_r16_c0_6;
  wire [7:0] t_r16_c0_7;
  wire [7:0] t_r16_c0_8;
  wire [7:0] t_r16_c0_9;
  wire [7:0] t_r16_c0_10;
  wire [7:0] t_r16_c0_11;
  wire [7:0] t_r16_c0_12;
  wire [7:0] t_r16_c1_0;
  wire [7:0] t_r16_c1_1;
  wire [7:0] t_r16_c1_2;
  wire [7:0] t_r16_c1_3;
  wire [7:0] t_r16_c1_4;
  wire [7:0] t_r16_c1_5;
  wire [7:0] t_r16_c1_6;
  wire [7:0] t_r16_c1_7;
  wire [7:0] t_r16_c1_8;
  wire [7:0] t_r16_c1_9;
  wire [7:0] t_r16_c1_10;
  wire [7:0] t_r16_c1_11;
  wire [7:0] t_r16_c1_12;
  wire [7:0] t_r16_c2_0;
  wire [7:0] t_r16_c2_1;
  wire [7:0] t_r16_c2_2;
  wire [7:0] t_r16_c2_3;
  wire [7:0] t_r16_c2_4;
  wire [7:0] t_r16_c2_5;
  wire [7:0] t_r16_c2_6;
  wire [7:0] t_r16_c2_7;
  wire [7:0] t_r16_c2_8;
  wire [7:0] t_r16_c2_9;
  wire [7:0] t_r16_c2_10;
  wire [7:0] t_r16_c2_11;
  wire [7:0] t_r16_c2_12;
  wire [7:0] t_r16_c3_0;
  wire [7:0] t_r16_c3_1;
  wire [7:0] t_r16_c3_2;
  wire [7:0] t_r16_c3_3;
  wire [7:0] t_r16_c3_4;
  wire [7:0] t_r16_c3_5;
  wire [7:0] t_r16_c3_6;
  wire [7:0] t_r16_c3_7;
  wire [7:0] t_r16_c3_8;
  wire [7:0] t_r16_c3_9;
  wire [7:0] t_r16_c3_10;
  wire [7:0] t_r16_c3_11;
  wire [7:0] t_r16_c3_12;
  wire [7:0] t_r16_c4_0;
  wire [7:0] t_r16_c4_1;
  wire [7:0] t_r16_c4_2;
  wire [7:0] t_r16_c4_3;
  wire [7:0] t_r16_c4_4;
  wire [7:0] t_r16_c4_5;
  wire [7:0] t_r16_c4_6;
  wire [7:0] t_r16_c4_7;
  wire [7:0] t_r16_c4_8;
  wire [7:0] t_r16_c4_9;
  wire [7:0] t_r16_c4_10;
  wire [7:0] t_r16_c4_11;
  wire [7:0] t_r16_c4_12;
  wire [7:0] t_r16_c5_0;
  wire [7:0] t_r16_c5_1;
  wire [7:0] t_r16_c5_2;
  wire [7:0] t_r16_c5_3;
  wire [7:0] t_r16_c5_4;
  wire [7:0] t_r16_c5_5;
  wire [7:0] t_r16_c5_6;
  wire [7:0] t_r16_c5_7;
  wire [7:0] t_r16_c5_8;
  wire [7:0] t_r16_c5_9;
  wire [7:0] t_r16_c5_10;
  wire [7:0] t_r16_c5_11;
  wire [7:0] t_r16_c5_12;
  wire [7:0] t_r16_c6_0;
  wire [7:0] t_r16_c6_1;
  wire [7:0] t_r16_c6_2;
  wire [7:0] t_r16_c6_3;
  wire [7:0] t_r16_c6_4;
  wire [7:0] t_r16_c6_5;
  wire [7:0] t_r16_c6_6;
  wire [7:0] t_r16_c6_7;
  wire [7:0] t_r16_c6_8;
  wire [7:0] t_r16_c6_9;
  wire [7:0] t_r16_c6_10;
  wire [7:0] t_r16_c6_11;
  wire [7:0] t_r16_c6_12;
  wire [7:0] t_r16_c7_0;
  wire [7:0] t_r16_c7_1;
  wire [7:0] t_r16_c7_2;
  wire [7:0] t_r16_c7_3;
  wire [7:0] t_r16_c7_4;
  wire [7:0] t_r16_c7_5;
  wire [7:0] t_r16_c7_6;
  wire [7:0] t_r16_c7_7;
  wire [7:0] t_r16_c7_8;
  wire [7:0] t_r16_c7_9;
  wire [7:0] t_r16_c7_10;
  wire [7:0] t_r16_c7_11;
  wire [7:0] t_r16_c7_12;
  wire [7:0] t_r16_c8_0;
  wire [7:0] t_r16_c8_1;
  wire [7:0] t_r16_c8_2;
  wire [7:0] t_r16_c8_3;
  wire [7:0] t_r16_c8_4;
  wire [7:0] t_r16_c8_5;
  wire [7:0] t_r16_c8_6;
  wire [7:0] t_r16_c8_7;
  wire [7:0] t_r16_c8_8;
  wire [7:0] t_r16_c8_9;
  wire [7:0] t_r16_c8_10;
  wire [7:0] t_r16_c8_11;
  wire [7:0] t_r16_c8_12;
  wire [7:0] t_r16_c9_0;
  wire [7:0] t_r16_c9_1;
  wire [7:0] t_r16_c9_2;
  wire [7:0] t_r16_c9_3;
  wire [7:0] t_r16_c9_4;
  wire [7:0] t_r16_c9_5;
  wire [7:0] t_r16_c9_6;
  wire [7:0] t_r16_c9_7;
  wire [7:0] t_r16_c9_8;
  wire [7:0] t_r16_c9_9;
  wire [7:0] t_r16_c9_10;
  wire [7:0] t_r16_c9_11;
  wire [7:0] t_r16_c9_12;
  wire [7:0] t_r16_c10_0;
  wire [7:0] t_r16_c10_1;
  wire [7:0] t_r16_c10_2;
  wire [7:0] t_r16_c10_3;
  wire [7:0] t_r16_c10_4;
  wire [7:0] t_r16_c10_5;
  wire [7:0] t_r16_c10_6;
  wire [7:0] t_r16_c10_7;
  wire [7:0] t_r16_c10_8;
  wire [7:0] t_r16_c10_9;
  wire [7:0] t_r16_c10_10;
  wire [7:0] t_r16_c10_11;
  wire [7:0] t_r16_c10_12;
  wire [7:0] t_r16_c11_0;
  wire [7:0] t_r16_c11_1;
  wire [7:0] t_r16_c11_2;
  wire [7:0] t_r16_c11_3;
  wire [7:0] t_r16_c11_4;
  wire [7:0] t_r16_c11_5;
  wire [7:0] t_r16_c11_6;
  wire [7:0] t_r16_c11_7;
  wire [7:0] t_r16_c11_8;
  wire [7:0] t_r16_c11_9;
  wire [7:0] t_r16_c11_10;
  wire [7:0] t_r16_c11_11;
  wire [7:0] t_r16_c11_12;
  wire [7:0] t_r16_c12_0;
  wire [7:0] t_r16_c12_1;
  wire [7:0] t_r16_c12_2;
  wire [7:0] t_r16_c12_3;
  wire [7:0] t_r16_c12_4;
  wire [7:0] t_r16_c12_5;
  wire [7:0] t_r16_c12_6;
  wire [7:0] t_r16_c12_7;
  wire [7:0] t_r16_c12_8;
  wire [7:0] t_r16_c12_9;
  wire [7:0] t_r16_c12_10;
  wire [7:0] t_r16_c12_11;
  wire [7:0] t_r16_c12_12;
  wire [7:0] t_r16_c13_0;
  wire [7:0] t_r16_c13_1;
  wire [7:0] t_r16_c13_2;
  wire [7:0] t_r16_c13_3;
  wire [7:0] t_r16_c13_4;
  wire [7:0] t_r16_c13_5;
  wire [7:0] t_r16_c13_6;
  wire [7:0] t_r16_c13_7;
  wire [7:0] t_r16_c13_8;
  wire [7:0] t_r16_c13_9;
  wire [7:0] t_r16_c13_10;
  wire [7:0] t_r16_c13_11;
  wire [7:0] t_r16_c13_12;
  wire [7:0] t_r16_c14_0;
  wire [7:0] t_r16_c14_1;
  wire [7:0] t_r16_c14_2;
  wire [7:0] t_r16_c14_3;
  wire [7:0] t_r16_c14_4;
  wire [7:0] t_r16_c14_5;
  wire [7:0] t_r16_c14_6;
  wire [7:0] t_r16_c14_7;
  wire [7:0] t_r16_c14_8;
  wire [7:0] t_r16_c14_9;
  wire [7:0] t_r16_c14_10;
  wire [7:0] t_r16_c14_11;
  wire [7:0] t_r16_c14_12;
  wire [7:0] t_r16_c15_0;
  wire [7:0] t_r16_c15_1;
  wire [7:0] t_r16_c15_2;
  wire [7:0] t_r16_c15_3;
  wire [7:0] t_r16_c15_4;
  wire [7:0] t_r16_c15_5;
  wire [7:0] t_r16_c15_6;
  wire [7:0] t_r16_c15_7;
  wire [7:0] t_r16_c15_8;
  wire [7:0] t_r16_c15_9;
  wire [7:0] t_r16_c15_10;
  wire [7:0] t_r16_c15_11;
  wire [7:0] t_r16_c15_12;
  wire [7:0] t_r16_c16_0;
  wire [7:0] t_r16_c16_1;
  wire [7:0] t_r16_c16_2;
  wire [7:0] t_r16_c16_3;
  wire [7:0] t_r16_c16_4;
  wire [7:0] t_r16_c16_5;
  wire [7:0] t_r16_c16_6;
  wire [7:0] t_r16_c16_7;
  wire [7:0] t_r16_c16_8;
  wire [7:0] t_r16_c16_9;
  wire [7:0] t_r16_c16_10;
  wire [7:0] t_r16_c16_11;
  wire [7:0] t_r16_c16_12;
  wire [7:0] t_r16_c17_0;
  wire [7:0] t_r16_c17_1;
  wire [7:0] t_r16_c17_2;
  wire [7:0] t_r16_c17_3;
  wire [7:0] t_r16_c17_4;
  wire [7:0] t_r16_c17_5;
  wire [7:0] t_r16_c17_6;
  wire [7:0] t_r16_c17_7;
  wire [7:0] t_r16_c17_8;
  wire [7:0] t_r16_c17_9;
  wire [7:0] t_r16_c17_10;
  wire [7:0] t_r16_c17_11;
  wire [7:0] t_r16_c17_12;
  wire [7:0] t_r16_c18_0;
  wire [7:0] t_r16_c18_1;
  wire [7:0] t_r16_c18_2;
  wire [7:0] t_r16_c18_3;
  wire [7:0] t_r16_c18_4;
  wire [7:0] t_r16_c18_5;
  wire [7:0] t_r16_c18_6;
  wire [7:0] t_r16_c18_7;
  wire [7:0] t_r16_c18_8;
  wire [7:0] t_r16_c18_9;
  wire [7:0] t_r16_c18_10;
  wire [7:0] t_r16_c18_11;
  wire [7:0] t_r16_c18_12;
  wire [7:0] t_r16_c19_0;
  wire [7:0] t_r16_c19_1;
  wire [7:0] t_r16_c19_2;
  wire [7:0] t_r16_c19_3;
  wire [7:0] t_r16_c19_4;
  wire [7:0] t_r16_c19_5;
  wire [7:0] t_r16_c19_6;
  wire [7:0] t_r16_c19_7;
  wire [7:0] t_r16_c19_8;
  wire [7:0] t_r16_c19_9;
  wire [7:0] t_r16_c19_10;
  wire [7:0] t_r16_c19_11;
  wire [7:0] t_r16_c19_12;
  wire [7:0] t_r16_c20_0;
  wire [7:0] t_r16_c20_1;
  wire [7:0] t_r16_c20_2;
  wire [7:0] t_r16_c20_3;
  wire [7:0] t_r16_c20_4;
  wire [7:0] t_r16_c20_5;
  wire [7:0] t_r16_c20_6;
  wire [7:0] t_r16_c20_7;
  wire [7:0] t_r16_c20_8;
  wire [7:0] t_r16_c20_9;
  wire [7:0] t_r16_c20_10;
  wire [7:0] t_r16_c20_11;
  wire [7:0] t_r16_c20_12;
  wire [7:0] t_r16_c21_0;
  wire [7:0] t_r16_c21_1;
  wire [7:0] t_r16_c21_2;
  wire [7:0] t_r16_c21_3;
  wire [7:0] t_r16_c21_4;
  wire [7:0] t_r16_c21_5;
  wire [7:0] t_r16_c21_6;
  wire [7:0] t_r16_c21_7;
  wire [7:0] t_r16_c21_8;
  wire [7:0] t_r16_c21_9;
  wire [7:0] t_r16_c21_10;
  wire [7:0] t_r16_c21_11;
  wire [7:0] t_r16_c21_12;
  wire [7:0] t_r16_c22_0;
  wire [7:0] t_r16_c22_1;
  wire [7:0] t_r16_c22_2;
  wire [7:0] t_r16_c22_3;
  wire [7:0] t_r16_c22_4;
  wire [7:0] t_r16_c22_5;
  wire [7:0] t_r16_c22_6;
  wire [7:0] t_r16_c22_7;
  wire [7:0] t_r16_c22_8;
  wire [7:0] t_r16_c22_9;
  wire [7:0] t_r16_c22_10;
  wire [7:0] t_r16_c22_11;
  wire [7:0] t_r16_c22_12;
  wire [7:0] t_r16_c23_0;
  wire [7:0] t_r16_c23_1;
  wire [7:0] t_r16_c23_2;
  wire [7:0] t_r16_c23_3;
  wire [7:0] t_r16_c23_4;
  wire [7:0] t_r16_c23_5;
  wire [7:0] t_r16_c23_6;
  wire [7:0] t_r16_c23_7;
  wire [7:0] t_r16_c23_8;
  wire [7:0] t_r16_c23_9;
  wire [7:0] t_r16_c23_10;
  wire [7:0] t_r16_c23_11;
  wire [7:0] t_r16_c23_12;
  wire [7:0] t_r16_c24_0;
  wire [7:0] t_r16_c24_1;
  wire [7:0] t_r16_c24_2;
  wire [7:0] t_r16_c24_3;
  wire [7:0] t_r16_c24_4;
  wire [7:0] t_r16_c24_5;
  wire [7:0] t_r16_c24_6;
  wire [7:0] t_r16_c24_7;
  wire [7:0] t_r16_c24_8;
  wire [7:0] t_r16_c24_9;
  wire [7:0] t_r16_c24_10;
  wire [7:0] t_r16_c24_11;
  wire [7:0] t_r16_c24_12;
  wire [7:0] t_r16_c25_0;
  wire [7:0] t_r16_c25_1;
  wire [7:0] t_r16_c25_2;
  wire [7:0] t_r16_c25_3;
  wire [7:0] t_r16_c25_4;
  wire [7:0] t_r16_c25_5;
  wire [7:0] t_r16_c25_6;
  wire [7:0] t_r16_c25_7;
  wire [7:0] t_r16_c25_8;
  wire [7:0] t_r16_c25_9;
  wire [7:0] t_r16_c25_10;
  wire [7:0] t_r16_c25_11;
  wire [7:0] t_r16_c25_12;
  wire [7:0] t_r16_c26_0;
  wire [7:0] t_r16_c26_1;
  wire [7:0] t_r16_c26_2;
  wire [7:0] t_r16_c26_3;
  wire [7:0] t_r16_c26_4;
  wire [7:0] t_r16_c26_5;
  wire [7:0] t_r16_c26_6;
  wire [7:0] t_r16_c26_7;
  wire [7:0] t_r16_c26_8;
  wire [7:0] t_r16_c26_9;
  wire [7:0] t_r16_c26_10;
  wire [7:0] t_r16_c26_11;
  wire [7:0] t_r16_c26_12;
  wire [7:0] t_r16_c27_0;
  wire [7:0] t_r16_c27_1;
  wire [7:0] t_r16_c27_2;
  wire [7:0] t_r16_c27_3;
  wire [7:0] t_r16_c27_4;
  wire [7:0] t_r16_c27_5;
  wire [7:0] t_r16_c27_6;
  wire [7:0] t_r16_c27_7;
  wire [7:0] t_r16_c27_8;
  wire [7:0] t_r16_c27_9;
  wire [7:0] t_r16_c27_10;
  wire [7:0] t_r16_c27_11;
  wire [7:0] t_r16_c27_12;
  wire [7:0] t_r16_c28_0;
  wire [7:0] t_r16_c28_1;
  wire [7:0] t_r16_c28_2;
  wire [7:0] t_r16_c28_3;
  wire [7:0] t_r16_c28_4;
  wire [7:0] t_r16_c28_5;
  wire [7:0] t_r16_c28_6;
  wire [7:0] t_r16_c28_7;
  wire [7:0] t_r16_c28_8;
  wire [7:0] t_r16_c28_9;
  wire [7:0] t_r16_c28_10;
  wire [7:0] t_r16_c28_11;
  wire [7:0] t_r16_c28_12;
  wire [7:0] t_r16_c29_0;
  wire [7:0] t_r16_c29_1;
  wire [7:0] t_r16_c29_2;
  wire [7:0] t_r16_c29_3;
  wire [7:0] t_r16_c29_4;
  wire [7:0] t_r16_c29_5;
  wire [7:0] t_r16_c29_6;
  wire [7:0] t_r16_c29_7;
  wire [7:0] t_r16_c29_8;
  wire [7:0] t_r16_c29_9;
  wire [7:0] t_r16_c29_10;
  wire [7:0] t_r16_c29_11;
  wire [7:0] t_r16_c29_12;
  wire [7:0] t_r16_c30_0;
  wire [7:0] t_r16_c30_1;
  wire [7:0] t_r16_c30_2;
  wire [7:0] t_r16_c30_3;
  wire [7:0] t_r16_c30_4;
  wire [7:0] t_r16_c30_5;
  wire [7:0] t_r16_c30_6;
  wire [7:0] t_r16_c30_7;
  wire [7:0] t_r16_c30_8;
  wire [7:0] t_r16_c30_9;
  wire [7:0] t_r16_c30_10;
  wire [7:0] t_r16_c30_11;
  wire [7:0] t_r16_c30_12;
  wire [7:0] t_r16_c31_0;
  wire [7:0] t_r16_c31_1;
  wire [7:0] t_r16_c31_2;
  wire [7:0] t_r16_c31_3;
  wire [7:0] t_r16_c31_4;
  wire [7:0] t_r16_c31_5;
  wire [7:0] t_r16_c31_6;
  wire [7:0] t_r16_c31_7;
  wire [7:0] t_r16_c31_8;
  wire [7:0] t_r16_c31_9;
  wire [7:0] t_r16_c31_10;
  wire [7:0] t_r16_c31_11;
  wire [7:0] t_r16_c31_12;
  wire [7:0] t_r16_c32_0;
  wire [7:0] t_r16_c32_1;
  wire [7:0] t_r16_c32_2;
  wire [7:0] t_r16_c32_3;
  wire [7:0] t_r16_c32_4;
  wire [7:0] t_r16_c32_5;
  wire [7:0] t_r16_c32_6;
  wire [7:0] t_r16_c32_7;
  wire [7:0] t_r16_c32_8;
  wire [7:0] t_r16_c32_9;
  wire [7:0] t_r16_c32_10;
  wire [7:0] t_r16_c32_11;
  wire [7:0] t_r16_c32_12;
  wire [7:0] t_r16_c33_0;
  wire [7:0] t_r16_c33_1;
  wire [7:0] t_r16_c33_2;
  wire [7:0] t_r16_c33_3;
  wire [7:0] t_r16_c33_4;
  wire [7:0] t_r16_c33_5;
  wire [7:0] t_r16_c33_6;
  wire [7:0] t_r16_c33_7;
  wire [7:0] t_r16_c33_8;
  wire [7:0] t_r16_c33_9;
  wire [7:0] t_r16_c33_10;
  wire [7:0] t_r16_c33_11;
  wire [7:0] t_r16_c33_12;
  wire [7:0] t_r16_c34_0;
  wire [7:0] t_r16_c34_1;
  wire [7:0] t_r16_c34_2;
  wire [7:0] t_r16_c34_3;
  wire [7:0] t_r16_c34_4;
  wire [7:0] t_r16_c34_5;
  wire [7:0] t_r16_c34_6;
  wire [7:0] t_r16_c34_7;
  wire [7:0] t_r16_c34_8;
  wire [7:0] t_r16_c34_9;
  wire [7:0] t_r16_c34_10;
  wire [7:0] t_r16_c34_11;
  wire [7:0] t_r16_c34_12;
  wire [7:0] t_r16_c35_0;
  wire [7:0] t_r16_c35_1;
  wire [7:0] t_r16_c35_2;
  wire [7:0] t_r16_c35_3;
  wire [7:0] t_r16_c35_4;
  wire [7:0] t_r16_c35_5;
  wire [7:0] t_r16_c35_6;
  wire [7:0] t_r16_c35_7;
  wire [7:0] t_r16_c35_8;
  wire [7:0] t_r16_c35_9;
  wire [7:0] t_r16_c35_10;
  wire [7:0] t_r16_c35_11;
  wire [7:0] t_r16_c35_12;
  wire [7:0] t_r16_c36_0;
  wire [7:0] t_r16_c36_1;
  wire [7:0] t_r16_c36_2;
  wire [7:0] t_r16_c36_3;
  wire [7:0] t_r16_c36_4;
  wire [7:0] t_r16_c36_5;
  wire [7:0] t_r16_c36_6;
  wire [7:0] t_r16_c36_7;
  wire [7:0] t_r16_c36_8;
  wire [7:0] t_r16_c36_9;
  wire [7:0] t_r16_c36_10;
  wire [7:0] t_r16_c36_11;
  wire [7:0] t_r16_c36_12;
  wire [7:0] t_r16_c37_0;
  wire [7:0] t_r16_c37_1;
  wire [7:0] t_r16_c37_2;
  wire [7:0] t_r16_c37_3;
  wire [7:0] t_r16_c37_4;
  wire [7:0] t_r16_c37_5;
  wire [7:0] t_r16_c37_6;
  wire [7:0] t_r16_c37_7;
  wire [7:0] t_r16_c37_8;
  wire [7:0] t_r16_c37_9;
  wire [7:0] t_r16_c37_10;
  wire [7:0] t_r16_c37_11;
  wire [7:0] t_r16_c37_12;
  wire [7:0] t_r16_c38_0;
  wire [7:0] t_r16_c38_1;
  wire [7:0] t_r16_c38_2;
  wire [7:0] t_r16_c38_3;
  wire [7:0] t_r16_c38_4;
  wire [7:0] t_r16_c38_5;
  wire [7:0] t_r16_c38_6;
  wire [7:0] t_r16_c38_7;
  wire [7:0] t_r16_c38_8;
  wire [7:0] t_r16_c38_9;
  wire [7:0] t_r16_c38_10;
  wire [7:0] t_r16_c38_11;
  wire [7:0] t_r16_c38_12;
  wire [7:0] t_r16_c39_0;
  wire [7:0] t_r16_c39_1;
  wire [7:0] t_r16_c39_2;
  wire [7:0] t_r16_c39_3;
  wire [7:0] t_r16_c39_4;
  wire [7:0] t_r16_c39_5;
  wire [7:0] t_r16_c39_6;
  wire [7:0] t_r16_c39_7;
  wire [7:0] t_r16_c39_8;
  wire [7:0] t_r16_c39_9;
  wire [7:0] t_r16_c39_10;
  wire [7:0] t_r16_c39_11;
  wire [7:0] t_r16_c39_12;
  wire [7:0] t_r16_c40_0;
  wire [7:0] t_r16_c40_1;
  wire [7:0] t_r16_c40_2;
  wire [7:0] t_r16_c40_3;
  wire [7:0] t_r16_c40_4;
  wire [7:0] t_r16_c40_5;
  wire [7:0] t_r16_c40_6;
  wire [7:0] t_r16_c40_7;
  wire [7:0] t_r16_c40_8;
  wire [7:0] t_r16_c40_9;
  wire [7:0] t_r16_c40_10;
  wire [7:0] t_r16_c40_11;
  wire [7:0] t_r16_c40_12;
  wire [7:0] t_r16_c41_0;
  wire [7:0] t_r16_c41_1;
  wire [7:0] t_r16_c41_2;
  wire [7:0] t_r16_c41_3;
  wire [7:0] t_r16_c41_4;
  wire [7:0] t_r16_c41_5;
  wire [7:0] t_r16_c41_6;
  wire [7:0] t_r16_c41_7;
  wire [7:0] t_r16_c41_8;
  wire [7:0] t_r16_c41_9;
  wire [7:0] t_r16_c41_10;
  wire [7:0] t_r16_c41_11;
  wire [7:0] t_r16_c41_12;
  wire [7:0] t_r16_c42_0;
  wire [7:0] t_r16_c42_1;
  wire [7:0] t_r16_c42_2;
  wire [7:0] t_r16_c42_3;
  wire [7:0] t_r16_c42_4;
  wire [7:0] t_r16_c42_5;
  wire [7:0] t_r16_c42_6;
  wire [7:0] t_r16_c42_7;
  wire [7:0] t_r16_c42_8;
  wire [7:0] t_r16_c42_9;
  wire [7:0] t_r16_c42_10;
  wire [7:0] t_r16_c42_11;
  wire [7:0] t_r16_c42_12;
  wire [7:0] t_r16_c43_0;
  wire [7:0] t_r16_c43_1;
  wire [7:0] t_r16_c43_2;
  wire [7:0] t_r16_c43_3;
  wire [7:0] t_r16_c43_4;
  wire [7:0] t_r16_c43_5;
  wire [7:0] t_r16_c43_6;
  wire [7:0] t_r16_c43_7;
  wire [7:0] t_r16_c43_8;
  wire [7:0] t_r16_c43_9;
  wire [7:0] t_r16_c43_10;
  wire [7:0] t_r16_c43_11;
  wire [7:0] t_r16_c43_12;
  wire [7:0] t_r16_c44_0;
  wire [7:0] t_r16_c44_1;
  wire [7:0] t_r16_c44_2;
  wire [7:0] t_r16_c44_3;
  wire [7:0] t_r16_c44_4;
  wire [7:0] t_r16_c44_5;
  wire [7:0] t_r16_c44_6;
  wire [7:0] t_r16_c44_7;
  wire [7:0] t_r16_c44_8;
  wire [7:0] t_r16_c44_9;
  wire [7:0] t_r16_c44_10;
  wire [7:0] t_r16_c44_11;
  wire [7:0] t_r16_c44_12;
  wire [7:0] t_r16_c45_0;
  wire [7:0] t_r16_c45_1;
  wire [7:0] t_r16_c45_2;
  wire [7:0] t_r16_c45_3;
  wire [7:0] t_r16_c45_4;
  wire [7:0] t_r16_c45_5;
  wire [7:0] t_r16_c45_6;
  wire [7:0] t_r16_c45_7;
  wire [7:0] t_r16_c45_8;
  wire [7:0] t_r16_c45_9;
  wire [7:0] t_r16_c45_10;
  wire [7:0] t_r16_c45_11;
  wire [7:0] t_r16_c45_12;
  wire [7:0] t_r16_c46_0;
  wire [7:0] t_r16_c46_1;
  wire [7:0] t_r16_c46_2;
  wire [7:0] t_r16_c46_3;
  wire [7:0] t_r16_c46_4;
  wire [7:0] t_r16_c46_5;
  wire [7:0] t_r16_c46_6;
  wire [7:0] t_r16_c46_7;
  wire [7:0] t_r16_c46_8;
  wire [7:0] t_r16_c46_9;
  wire [7:0] t_r16_c46_10;
  wire [7:0] t_r16_c46_11;
  wire [7:0] t_r16_c46_12;
  wire [7:0] t_r16_c47_0;
  wire [7:0] t_r16_c47_1;
  wire [7:0] t_r16_c47_2;
  wire [7:0] t_r16_c47_3;
  wire [7:0] t_r16_c47_4;
  wire [7:0] t_r16_c47_5;
  wire [7:0] t_r16_c47_6;
  wire [7:0] t_r16_c47_7;
  wire [7:0] t_r16_c47_8;
  wire [7:0] t_r16_c47_9;
  wire [7:0] t_r16_c47_10;
  wire [7:0] t_r16_c47_11;
  wire [7:0] t_r16_c47_12;
  wire [7:0] t_r16_c48_0;
  wire [7:0] t_r16_c48_1;
  wire [7:0] t_r16_c48_2;
  wire [7:0] t_r16_c48_3;
  wire [7:0] t_r16_c48_4;
  wire [7:0] t_r16_c48_5;
  wire [7:0] t_r16_c48_6;
  wire [7:0] t_r16_c48_7;
  wire [7:0] t_r16_c48_8;
  wire [7:0] t_r16_c48_9;
  wire [7:0] t_r16_c48_10;
  wire [7:0] t_r16_c48_11;
  wire [7:0] t_r16_c48_12;
  wire [7:0] t_r16_c49_0;
  wire [7:0] t_r16_c49_1;
  wire [7:0] t_r16_c49_2;
  wire [7:0] t_r16_c49_3;
  wire [7:0] t_r16_c49_4;
  wire [7:0] t_r16_c49_5;
  wire [7:0] t_r16_c49_6;
  wire [7:0] t_r16_c49_7;
  wire [7:0] t_r16_c49_8;
  wire [7:0] t_r16_c49_9;
  wire [7:0] t_r16_c49_10;
  wire [7:0] t_r16_c49_11;
  wire [7:0] t_r16_c49_12;
  wire [7:0] t_r16_c50_0;
  wire [7:0] t_r16_c50_1;
  wire [7:0] t_r16_c50_2;
  wire [7:0] t_r16_c50_3;
  wire [7:0] t_r16_c50_4;
  wire [7:0] t_r16_c50_5;
  wire [7:0] t_r16_c50_6;
  wire [7:0] t_r16_c50_7;
  wire [7:0] t_r16_c50_8;
  wire [7:0] t_r16_c50_9;
  wire [7:0] t_r16_c50_10;
  wire [7:0] t_r16_c50_11;
  wire [7:0] t_r16_c50_12;
  wire [7:0] t_r16_c51_0;
  wire [7:0] t_r16_c51_1;
  wire [7:0] t_r16_c51_2;
  wire [7:0] t_r16_c51_3;
  wire [7:0] t_r16_c51_4;
  wire [7:0] t_r16_c51_5;
  wire [7:0] t_r16_c51_6;
  wire [7:0] t_r16_c51_7;
  wire [7:0] t_r16_c51_8;
  wire [7:0] t_r16_c51_9;
  wire [7:0] t_r16_c51_10;
  wire [7:0] t_r16_c51_11;
  wire [7:0] t_r16_c51_12;
  wire [7:0] t_r16_c52_0;
  wire [7:0] t_r16_c52_1;
  wire [7:0] t_r16_c52_2;
  wire [7:0] t_r16_c52_3;
  wire [7:0] t_r16_c52_4;
  wire [7:0] t_r16_c52_5;
  wire [7:0] t_r16_c52_6;
  wire [7:0] t_r16_c52_7;
  wire [7:0] t_r16_c52_8;
  wire [7:0] t_r16_c52_9;
  wire [7:0] t_r16_c52_10;
  wire [7:0] t_r16_c52_11;
  wire [7:0] t_r16_c52_12;
  wire [7:0] t_r16_c53_0;
  wire [7:0] t_r16_c53_1;
  wire [7:0] t_r16_c53_2;
  wire [7:0] t_r16_c53_3;
  wire [7:0] t_r16_c53_4;
  wire [7:0] t_r16_c53_5;
  wire [7:0] t_r16_c53_6;
  wire [7:0] t_r16_c53_7;
  wire [7:0] t_r16_c53_8;
  wire [7:0] t_r16_c53_9;
  wire [7:0] t_r16_c53_10;
  wire [7:0] t_r16_c53_11;
  wire [7:0] t_r16_c53_12;
  wire [7:0] t_r16_c54_0;
  wire [7:0] t_r16_c54_1;
  wire [7:0] t_r16_c54_2;
  wire [7:0] t_r16_c54_3;
  wire [7:0] t_r16_c54_4;
  wire [7:0] t_r16_c54_5;
  wire [7:0] t_r16_c54_6;
  wire [7:0] t_r16_c54_7;
  wire [7:0] t_r16_c54_8;
  wire [7:0] t_r16_c54_9;
  wire [7:0] t_r16_c54_10;
  wire [7:0] t_r16_c54_11;
  wire [7:0] t_r16_c54_12;
  wire [7:0] t_r16_c55_0;
  wire [7:0] t_r16_c55_1;
  wire [7:0] t_r16_c55_2;
  wire [7:0] t_r16_c55_3;
  wire [7:0] t_r16_c55_4;
  wire [7:0] t_r16_c55_5;
  wire [7:0] t_r16_c55_6;
  wire [7:0] t_r16_c55_7;
  wire [7:0] t_r16_c55_8;
  wire [7:0] t_r16_c55_9;
  wire [7:0] t_r16_c55_10;
  wire [7:0] t_r16_c55_11;
  wire [7:0] t_r16_c55_12;
  wire [7:0] t_r16_c56_0;
  wire [7:0] t_r16_c56_1;
  wire [7:0] t_r16_c56_2;
  wire [7:0] t_r16_c56_3;
  wire [7:0] t_r16_c56_4;
  wire [7:0] t_r16_c56_5;
  wire [7:0] t_r16_c56_6;
  wire [7:0] t_r16_c56_7;
  wire [7:0] t_r16_c56_8;
  wire [7:0] t_r16_c56_9;
  wire [7:0] t_r16_c56_10;
  wire [7:0] t_r16_c56_11;
  wire [7:0] t_r16_c56_12;
  wire [7:0] t_r16_c57_0;
  wire [7:0] t_r16_c57_1;
  wire [7:0] t_r16_c57_2;
  wire [7:0] t_r16_c57_3;
  wire [7:0] t_r16_c57_4;
  wire [7:0] t_r16_c57_5;
  wire [7:0] t_r16_c57_6;
  wire [7:0] t_r16_c57_7;
  wire [7:0] t_r16_c57_8;
  wire [7:0] t_r16_c57_9;
  wire [7:0] t_r16_c57_10;
  wire [7:0] t_r16_c57_11;
  wire [7:0] t_r16_c57_12;
  wire [7:0] t_r16_c58_0;
  wire [7:0] t_r16_c58_1;
  wire [7:0] t_r16_c58_2;
  wire [7:0] t_r16_c58_3;
  wire [7:0] t_r16_c58_4;
  wire [7:0] t_r16_c58_5;
  wire [7:0] t_r16_c58_6;
  wire [7:0] t_r16_c58_7;
  wire [7:0] t_r16_c58_8;
  wire [7:0] t_r16_c58_9;
  wire [7:0] t_r16_c58_10;
  wire [7:0] t_r16_c58_11;
  wire [7:0] t_r16_c58_12;
  wire [7:0] t_r16_c59_0;
  wire [7:0] t_r16_c59_1;
  wire [7:0] t_r16_c59_2;
  wire [7:0] t_r16_c59_3;
  wire [7:0] t_r16_c59_4;
  wire [7:0] t_r16_c59_5;
  wire [7:0] t_r16_c59_6;
  wire [7:0] t_r16_c59_7;
  wire [7:0] t_r16_c59_8;
  wire [7:0] t_r16_c59_9;
  wire [7:0] t_r16_c59_10;
  wire [7:0] t_r16_c59_11;
  wire [7:0] t_r16_c59_12;
  wire [7:0] t_r16_c60_0;
  wire [7:0] t_r16_c60_1;
  wire [7:0] t_r16_c60_2;
  wire [7:0] t_r16_c60_3;
  wire [7:0] t_r16_c60_4;
  wire [7:0] t_r16_c60_5;
  wire [7:0] t_r16_c60_6;
  wire [7:0] t_r16_c60_7;
  wire [7:0] t_r16_c60_8;
  wire [7:0] t_r16_c60_9;
  wire [7:0] t_r16_c60_10;
  wire [7:0] t_r16_c60_11;
  wire [7:0] t_r16_c60_12;
  wire [7:0] t_r16_c61_0;
  wire [7:0] t_r16_c61_1;
  wire [7:0] t_r16_c61_2;
  wire [7:0] t_r16_c61_3;
  wire [7:0] t_r16_c61_4;
  wire [7:0] t_r16_c61_5;
  wire [7:0] t_r16_c61_6;
  wire [7:0] t_r16_c61_7;
  wire [7:0] t_r16_c61_8;
  wire [7:0] t_r16_c61_9;
  wire [7:0] t_r16_c61_10;
  wire [7:0] t_r16_c61_11;
  wire [7:0] t_r16_c61_12;
  wire [7:0] t_r16_c62_0;
  wire [7:0] t_r16_c62_1;
  wire [7:0] t_r16_c62_2;
  wire [7:0] t_r16_c62_3;
  wire [7:0] t_r16_c62_4;
  wire [7:0] t_r16_c62_5;
  wire [7:0] t_r16_c62_6;
  wire [7:0] t_r16_c62_7;
  wire [7:0] t_r16_c62_8;
  wire [7:0] t_r16_c62_9;
  wire [7:0] t_r16_c62_10;
  wire [7:0] t_r16_c62_11;
  wire [7:0] t_r16_c62_12;
  wire [7:0] t_r16_c63_0;
  wire [7:0] t_r16_c63_1;
  wire [7:0] t_r16_c63_2;
  wire [7:0] t_r16_c63_3;
  wire [7:0] t_r16_c63_4;
  wire [7:0] t_r16_c63_5;
  wire [7:0] t_r16_c63_6;
  wire [7:0] t_r16_c63_7;
  wire [7:0] t_r16_c63_8;
  wire [7:0] t_r16_c63_9;
  wire [7:0] t_r16_c63_10;
  wire [7:0] t_r16_c63_11;
  wire [7:0] t_r16_c63_12;
  wire [7:0] t_r16_c64_0;
  wire [7:0] t_r16_c64_1;
  wire [7:0] t_r16_c64_2;
  wire [7:0] t_r16_c64_3;
  wire [7:0] t_r16_c64_4;
  wire [7:0] t_r16_c64_5;
  wire [7:0] t_r16_c64_6;
  wire [7:0] t_r16_c64_7;
  wire [7:0] t_r16_c64_8;
  wire [7:0] t_r16_c64_9;
  wire [7:0] t_r16_c64_10;
  wire [7:0] t_r16_c64_11;
  wire [7:0] t_r16_c64_12;
  wire [7:0] t_r16_c65_0;
  wire [7:0] t_r16_c65_1;
  wire [7:0] t_r16_c65_2;
  wire [7:0] t_r16_c65_3;
  wire [7:0] t_r16_c65_4;
  wire [7:0] t_r16_c65_5;
  wire [7:0] t_r16_c65_6;
  wire [7:0] t_r16_c65_7;
  wire [7:0] t_r16_c65_8;
  wire [7:0] t_r16_c65_9;
  wire [7:0] t_r16_c65_10;
  wire [7:0] t_r16_c65_11;
  wire [7:0] t_r16_c65_12;
  wire [7:0] t_r17_c0_0;
  wire [7:0] t_r17_c0_1;
  wire [7:0] t_r17_c0_2;
  wire [7:0] t_r17_c0_3;
  wire [7:0] t_r17_c0_4;
  wire [7:0] t_r17_c0_5;
  wire [7:0] t_r17_c0_6;
  wire [7:0] t_r17_c0_7;
  wire [7:0] t_r17_c0_8;
  wire [7:0] t_r17_c0_9;
  wire [7:0] t_r17_c0_10;
  wire [7:0] t_r17_c0_11;
  wire [7:0] t_r17_c0_12;
  wire [7:0] t_r17_c1_0;
  wire [7:0] t_r17_c1_1;
  wire [7:0] t_r17_c1_2;
  wire [7:0] t_r17_c1_3;
  wire [7:0] t_r17_c1_4;
  wire [7:0] t_r17_c1_5;
  wire [7:0] t_r17_c1_6;
  wire [7:0] t_r17_c1_7;
  wire [7:0] t_r17_c1_8;
  wire [7:0] t_r17_c1_9;
  wire [7:0] t_r17_c1_10;
  wire [7:0] t_r17_c1_11;
  wire [7:0] t_r17_c1_12;
  wire [7:0] t_r17_c2_0;
  wire [7:0] t_r17_c2_1;
  wire [7:0] t_r17_c2_2;
  wire [7:0] t_r17_c2_3;
  wire [7:0] t_r17_c2_4;
  wire [7:0] t_r17_c2_5;
  wire [7:0] t_r17_c2_6;
  wire [7:0] t_r17_c2_7;
  wire [7:0] t_r17_c2_8;
  wire [7:0] t_r17_c2_9;
  wire [7:0] t_r17_c2_10;
  wire [7:0] t_r17_c2_11;
  wire [7:0] t_r17_c2_12;
  wire [7:0] t_r17_c3_0;
  wire [7:0] t_r17_c3_1;
  wire [7:0] t_r17_c3_2;
  wire [7:0] t_r17_c3_3;
  wire [7:0] t_r17_c3_4;
  wire [7:0] t_r17_c3_5;
  wire [7:0] t_r17_c3_6;
  wire [7:0] t_r17_c3_7;
  wire [7:0] t_r17_c3_8;
  wire [7:0] t_r17_c3_9;
  wire [7:0] t_r17_c3_10;
  wire [7:0] t_r17_c3_11;
  wire [7:0] t_r17_c3_12;
  wire [7:0] t_r17_c4_0;
  wire [7:0] t_r17_c4_1;
  wire [7:0] t_r17_c4_2;
  wire [7:0] t_r17_c4_3;
  wire [7:0] t_r17_c4_4;
  wire [7:0] t_r17_c4_5;
  wire [7:0] t_r17_c4_6;
  wire [7:0] t_r17_c4_7;
  wire [7:0] t_r17_c4_8;
  wire [7:0] t_r17_c4_9;
  wire [7:0] t_r17_c4_10;
  wire [7:0] t_r17_c4_11;
  wire [7:0] t_r17_c4_12;
  wire [7:0] t_r17_c5_0;
  wire [7:0] t_r17_c5_1;
  wire [7:0] t_r17_c5_2;
  wire [7:0] t_r17_c5_3;
  wire [7:0] t_r17_c5_4;
  wire [7:0] t_r17_c5_5;
  wire [7:0] t_r17_c5_6;
  wire [7:0] t_r17_c5_7;
  wire [7:0] t_r17_c5_8;
  wire [7:0] t_r17_c5_9;
  wire [7:0] t_r17_c5_10;
  wire [7:0] t_r17_c5_11;
  wire [7:0] t_r17_c5_12;
  wire [7:0] t_r17_c6_0;
  wire [7:0] t_r17_c6_1;
  wire [7:0] t_r17_c6_2;
  wire [7:0] t_r17_c6_3;
  wire [7:0] t_r17_c6_4;
  wire [7:0] t_r17_c6_5;
  wire [7:0] t_r17_c6_6;
  wire [7:0] t_r17_c6_7;
  wire [7:0] t_r17_c6_8;
  wire [7:0] t_r17_c6_9;
  wire [7:0] t_r17_c6_10;
  wire [7:0] t_r17_c6_11;
  wire [7:0] t_r17_c6_12;
  wire [7:0] t_r17_c7_0;
  wire [7:0] t_r17_c7_1;
  wire [7:0] t_r17_c7_2;
  wire [7:0] t_r17_c7_3;
  wire [7:0] t_r17_c7_4;
  wire [7:0] t_r17_c7_5;
  wire [7:0] t_r17_c7_6;
  wire [7:0] t_r17_c7_7;
  wire [7:0] t_r17_c7_8;
  wire [7:0] t_r17_c7_9;
  wire [7:0] t_r17_c7_10;
  wire [7:0] t_r17_c7_11;
  wire [7:0] t_r17_c7_12;
  wire [7:0] t_r17_c8_0;
  wire [7:0] t_r17_c8_1;
  wire [7:0] t_r17_c8_2;
  wire [7:0] t_r17_c8_3;
  wire [7:0] t_r17_c8_4;
  wire [7:0] t_r17_c8_5;
  wire [7:0] t_r17_c8_6;
  wire [7:0] t_r17_c8_7;
  wire [7:0] t_r17_c8_8;
  wire [7:0] t_r17_c8_9;
  wire [7:0] t_r17_c8_10;
  wire [7:0] t_r17_c8_11;
  wire [7:0] t_r17_c8_12;
  wire [7:0] t_r17_c9_0;
  wire [7:0] t_r17_c9_1;
  wire [7:0] t_r17_c9_2;
  wire [7:0] t_r17_c9_3;
  wire [7:0] t_r17_c9_4;
  wire [7:0] t_r17_c9_5;
  wire [7:0] t_r17_c9_6;
  wire [7:0] t_r17_c9_7;
  wire [7:0] t_r17_c9_8;
  wire [7:0] t_r17_c9_9;
  wire [7:0] t_r17_c9_10;
  wire [7:0] t_r17_c9_11;
  wire [7:0] t_r17_c9_12;
  wire [7:0] t_r17_c10_0;
  wire [7:0] t_r17_c10_1;
  wire [7:0] t_r17_c10_2;
  wire [7:0] t_r17_c10_3;
  wire [7:0] t_r17_c10_4;
  wire [7:0] t_r17_c10_5;
  wire [7:0] t_r17_c10_6;
  wire [7:0] t_r17_c10_7;
  wire [7:0] t_r17_c10_8;
  wire [7:0] t_r17_c10_9;
  wire [7:0] t_r17_c10_10;
  wire [7:0] t_r17_c10_11;
  wire [7:0] t_r17_c10_12;
  wire [7:0] t_r17_c11_0;
  wire [7:0] t_r17_c11_1;
  wire [7:0] t_r17_c11_2;
  wire [7:0] t_r17_c11_3;
  wire [7:0] t_r17_c11_4;
  wire [7:0] t_r17_c11_5;
  wire [7:0] t_r17_c11_6;
  wire [7:0] t_r17_c11_7;
  wire [7:0] t_r17_c11_8;
  wire [7:0] t_r17_c11_9;
  wire [7:0] t_r17_c11_10;
  wire [7:0] t_r17_c11_11;
  wire [7:0] t_r17_c11_12;
  wire [7:0] t_r17_c12_0;
  wire [7:0] t_r17_c12_1;
  wire [7:0] t_r17_c12_2;
  wire [7:0] t_r17_c12_3;
  wire [7:0] t_r17_c12_4;
  wire [7:0] t_r17_c12_5;
  wire [7:0] t_r17_c12_6;
  wire [7:0] t_r17_c12_7;
  wire [7:0] t_r17_c12_8;
  wire [7:0] t_r17_c12_9;
  wire [7:0] t_r17_c12_10;
  wire [7:0] t_r17_c12_11;
  wire [7:0] t_r17_c12_12;
  wire [7:0] t_r17_c13_0;
  wire [7:0] t_r17_c13_1;
  wire [7:0] t_r17_c13_2;
  wire [7:0] t_r17_c13_3;
  wire [7:0] t_r17_c13_4;
  wire [7:0] t_r17_c13_5;
  wire [7:0] t_r17_c13_6;
  wire [7:0] t_r17_c13_7;
  wire [7:0] t_r17_c13_8;
  wire [7:0] t_r17_c13_9;
  wire [7:0] t_r17_c13_10;
  wire [7:0] t_r17_c13_11;
  wire [7:0] t_r17_c13_12;
  wire [7:0] t_r17_c14_0;
  wire [7:0] t_r17_c14_1;
  wire [7:0] t_r17_c14_2;
  wire [7:0] t_r17_c14_3;
  wire [7:0] t_r17_c14_4;
  wire [7:0] t_r17_c14_5;
  wire [7:0] t_r17_c14_6;
  wire [7:0] t_r17_c14_7;
  wire [7:0] t_r17_c14_8;
  wire [7:0] t_r17_c14_9;
  wire [7:0] t_r17_c14_10;
  wire [7:0] t_r17_c14_11;
  wire [7:0] t_r17_c14_12;
  wire [7:0] t_r17_c15_0;
  wire [7:0] t_r17_c15_1;
  wire [7:0] t_r17_c15_2;
  wire [7:0] t_r17_c15_3;
  wire [7:0] t_r17_c15_4;
  wire [7:0] t_r17_c15_5;
  wire [7:0] t_r17_c15_6;
  wire [7:0] t_r17_c15_7;
  wire [7:0] t_r17_c15_8;
  wire [7:0] t_r17_c15_9;
  wire [7:0] t_r17_c15_10;
  wire [7:0] t_r17_c15_11;
  wire [7:0] t_r17_c15_12;
  wire [7:0] t_r17_c16_0;
  wire [7:0] t_r17_c16_1;
  wire [7:0] t_r17_c16_2;
  wire [7:0] t_r17_c16_3;
  wire [7:0] t_r17_c16_4;
  wire [7:0] t_r17_c16_5;
  wire [7:0] t_r17_c16_6;
  wire [7:0] t_r17_c16_7;
  wire [7:0] t_r17_c16_8;
  wire [7:0] t_r17_c16_9;
  wire [7:0] t_r17_c16_10;
  wire [7:0] t_r17_c16_11;
  wire [7:0] t_r17_c16_12;
  wire [7:0] t_r17_c17_0;
  wire [7:0] t_r17_c17_1;
  wire [7:0] t_r17_c17_2;
  wire [7:0] t_r17_c17_3;
  wire [7:0] t_r17_c17_4;
  wire [7:0] t_r17_c17_5;
  wire [7:0] t_r17_c17_6;
  wire [7:0] t_r17_c17_7;
  wire [7:0] t_r17_c17_8;
  wire [7:0] t_r17_c17_9;
  wire [7:0] t_r17_c17_10;
  wire [7:0] t_r17_c17_11;
  wire [7:0] t_r17_c17_12;
  wire [7:0] t_r17_c18_0;
  wire [7:0] t_r17_c18_1;
  wire [7:0] t_r17_c18_2;
  wire [7:0] t_r17_c18_3;
  wire [7:0] t_r17_c18_4;
  wire [7:0] t_r17_c18_5;
  wire [7:0] t_r17_c18_6;
  wire [7:0] t_r17_c18_7;
  wire [7:0] t_r17_c18_8;
  wire [7:0] t_r17_c18_9;
  wire [7:0] t_r17_c18_10;
  wire [7:0] t_r17_c18_11;
  wire [7:0] t_r17_c18_12;
  wire [7:0] t_r17_c19_0;
  wire [7:0] t_r17_c19_1;
  wire [7:0] t_r17_c19_2;
  wire [7:0] t_r17_c19_3;
  wire [7:0] t_r17_c19_4;
  wire [7:0] t_r17_c19_5;
  wire [7:0] t_r17_c19_6;
  wire [7:0] t_r17_c19_7;
  wire [7:0] t_r17_c19_8;
  wire [7:0] t_r17_c19_9;
  wire [7:0] t_r17_c19_10;
  wire [7:0] t_r17_c19_11;
  wire [7:0] t_r17_c19_12;
  wire [7:0] t_r17_c20_0;
  wire [7:0] t_r17_c20_1;
  wire [7:0] t_r17_c20_2;
  wire [7:0] t_r17_c20_3;
  wire [7:0] t_r17_c20_4;
  wire [7:0] t_r17_c20_5;
  wire [7:0] t_r17_c20_6;
  wire [7:0] t_r17_c20_7;
  wire [7:0] t_r17_c20_8;
  wire [7:0] t_r17_c20_9;
  wire [7:0] t_r17_c20_10;
  wire [7:0] t_r17_c20_11;
  wire [7:0] t_r17_c20_12;
  wire [7:0] t_r17_c21_0;
  wire [7:0] t_r17_c21_1;
  wire [7:0] t_r17_c21_2;
  wire [7:0] t_r17_c21_3;
  wire [7:0] t_r17_c21_4;
  wire [7:0] t_r17_c21_5;
  wire [7:0] t_r17_c21_6;
  wire [7:0] t_r17_c21_7;
  wire [7:0] t_r17_c21_8;
  wire [7:0] t_r17_c21_9;
  wire [7:0] t_r17_c21_10;
  wire [7:0] t_r17_c21_11;
  wire [7:0] t_r17_c21_12;
  wire [7:0] t_r17_c22_0;
  wire [7:0] t_r17_c22_1;
  wire [7:0] t_r17_c22_2;
  wire [7:0] t_r17_c22_3;
  wire [7:0] t_r17_c22_4;
  wire [7:0] t_r17_c22_5;
  wire [7:0] t_r17_c22_6;
  wire [7:0] t_r17_c22_7;
  wire [7:0] t_r17_c22_8;
  wire [7:0] t_r17_c22_9;
  wire [7:0] t_r17_c22_10;
  wire [7:0] t_r17_c22_11;
  wire [7:0] t_r17_c22_12;
  wire [7:0] t_r17_c23_0;
  wire [7:0] t_r17_c23_1;
  wire [7:0] t_r17_c23_2;
  wire [7:0] t_r17_c23_3;
  wire [7:0] t_r17_c23_4;
  wire [7:0] t_r17_c23_5;
  wire [7:0] t_r17_c23_6;
  wire [7:0] t_r17_c23_7;
  wire [7:0] t_r17_c23_8;
  wire [7:0] t_r17_c23_9;
  wire [7:0] t_r17_c23_10;
  wire [7:0] t_r17_c23_11;
  wire [7:0] t_r17_c23_12;
  wire [7:0] t_r17_c24_0;
  wire [7:0] t_r17_c24_1;
  wire [7:0] t_r17_c24_2;
  wire [7:0] t_r17_c24_3;
  wire [7:0] t_r17_c24_4;
  wire [7:0] t_r17_c24_5;
  wire [7:0] t_r17_c24_6;
  wire [7:0] t_r17_c24_7;
  wire [7:0] t_r17_c24_8;
  wire [7:0] t_r17_c24_9;
  wire [7:0] t_r17_c24_10;
  wire [7:0] t_r17_c24_11;
  wire [7:0] t_r17_c24_12;
  wire [7:0] t_r17_c25_0;
  wire [7:0] t_r17_c25_1;
  wire [7:0] t_r17_c25_2;
  wire [7:0] t_r17_c25_3;
  wire [7:0] t_r17_c25_4;
  wire [7:0] t_r17_c25_5;
  wire [7:0] t_r17_c25_6;
  wire [7:0] t_r17_c25_7;
  wire [7:0] t_r17_c25_8;
  wire [7:0] t_r17_c25_9;
  wire [7:0] t_r17_c25_10;
  wire [7:0] t_r17_c25_11;
  wire [7:0] t_r17_c25_12;
  wire [7:0] t_r17_c26_0;
  wire [7:0] t_r17_c26_1;
  wire [7:0] t_r17_c26_2;
  wire [7:0] t_r17_c26_3;
  wire [7:0] t_r17_c26_4;
  wire [7:0] t_r17_c26_5;
  wire [7:0] t_r17_c26_6;
  wire [7:0] t_r17_c26_7;
  wire [7:0] t_r17_c26_8;
  wire [7:0] t_r17_c26_9;
  wire [7:0] t_r17_c26_10;
  wire [7:0] t_r17_c26_11;
  wire [7:0] t_r17_c26_12;
  wire [7:0] t_r17_c27_0;
  wire [7:0] t_r17_c27_1;
  wire [7:0] t_r17_c27_2;
  wire [7:0] t_r17_c27_3;
  wire [7:0] t_r17_c27_4;
  wire [7:0] t_r17_c27_5;
  wire [7:0] t_r17_c27_6;
  wire [7:0] t_r17_c27_7;
  wire [7:0] t_r17_c27_8;
  wire [7:0] t_r17_c27_9;
  wire [7:0] t_r17_c27_10;
  wire [7:0] t_r17_c27_11;
  wire [7:0] t_r17_c27_12;
  wire [7:0] t_r17_c28_0;
  wire [7:0] t_r17_c28_1;
  wire [7:0] t_r17_c28_2;
  wire [7:0] t_r17_c28_3;
  wire [7:0] t_r17_c28_4;
  wire [7:0] t_r17_c28_5;
  wire [7:0] t_r17_c28_6;
  wire [7:0] t_r17_c28_7;
  wire [7:0] t_r17_c28_8;
  wire [7:0] t_r17_c28_9;
  wire [7:0] t_r17_c28_10;
  wire [7:0] t_r17_c28_11;
  wire [7:0] t_r17_c28_12;
  wire [7:0] t_r17_c29_0;
  wire [7:0] t_r17_c29_1;
  wire [7:0] t_r17_c29_2;
  wire [7:0] t_r17_c29_3;
  wire [7:0] t_r17_c29_4;
  wire [7:0] t_r17_c29_5;
  wire [7:0] t_r17_c29_6;
  wire [7:0] t_r17_c29_7;
  wire [7:0] t_r17_c29_8;
  wire [7:0] t_r17_c29_9;
  wire [7:0] t_r17_c29_10;
  wire [7:0] t_r17_c29_11;
  wire [7:0] t_r17_c29_12;
  wire [7:0] t_r17_c30_0;
  wire [7:0] t_r17_c30_1;
  wire [7:0] t_r17_c30_2;
  wire [7:0] t_r17_c30_3;
  wire [7:0] t_r17_c30_4;
  wire [7:0] t_r17_c30_5;
  wire [7:0] t_r17_c30_6;
  wire [7:0] t_r17_c30_7;
  wire [7:0] t_r17_c30_8;
  wire [7:0] t_r17_c30_9;
  wire [7:0] t_r17_c30_10;
  wire [7:0] t_r17_c30_11;
  wire [7:0] t_r17_c30_12;
  wire [7:0] t_r17_c31_0;
  wire [7:0] t_r17_c31_1;
  wire [7:0] t_r17_c31_2;
  wire [7:0] t_r17_c31_3;
  wire [7:0] t_r17_c31_4;
  wire [7:0] t_r17_c31_5;
  wire [7:0] t_r17_c31_6;
  wire [7:0] t_r17_c31_7;
  wire [7:0] t_r17_c31_8;
  wire [7:0] t_r17_c31_9;
  wire [7:0] t_r17_c31_10;
  wire [7:0] t_r17_c31_11;
  wire [7:0] t_r17_c31_12;
  wire [7:0] t_r17_c32_0;
  wire [7:0] t_r17_c32_1;
  wire [7:0] t_r17_c32_2;
  wire [7:0] t_r17_c32_3;
  wire [7:0] t_r17_c32_4;
  wire [7:0] t_r17_c32_5;
  wire [7:0] t_r17_c32_6;
  wire [7:0] t_r17_c32_7;
  wire [7:0] t_r17_c32_8;
  wire [7:0] t_r17_c32_9;
  wire [7:0] t_r17_c32_10;
  wire [7:0] t_r17_c32_11;
  wire [7:0] t_r17_c32_12;
  wire [7:0] t_r17_c33_0;
  wire [7:0] t_r17_c33_1;
  wire [7:0] t_r17_c33_2;
  wire [7:0] t_r17_c33_3;
  wire [7:0] t_r17_c33_4;
  wire [7:0] t_r17_c33_5;
  wire [7:0] t_r17_c33_6;
  wire [7:0] t_r17_c33_7;
  wire [7:0] t_r17_c33_8;
  wire [7:0] t_r17_c33_9;
  wire [7:0] t_r17_c33_10;
  wire [7:0] t_r17_c33_11;
  wire [7:0] t_r17_c33_12;
  wire [7:0] t_r17_c34_0;
  wire [7:0] t_r17_c34_1;
  wire [7:0] t_r17_c34_2;
  wire [7:0] t_r17_c34_3;
  wire [7:0] t_r17_c34_4;
  wire [7:0] t_r17_c34_5;
  wire [7:0] t_r17_c34_6;
  wire [7:0] t_r17_c34_7;
  wire [7:0] t_r17_c34_8;
  wire [7:0] t_r17_c34_9;
  wire [7:0] t_r17_c34_10;
  wire [7:0] t_r17_c34_11;
  wire [7:0] t_r17_c34_12;
  wire [7:0] t_r17_c35_0;
  wire [7:0] t_r17_c35_1;
  wire [7:0] t_r17_c35_2;
  wire [7:0] t_r17_c35_3;
  wire [7:0] t_r17_c35_4;
  wire [7:0] t_r17_c35_5;
  wire [7:0] t_r17_c35_6;
  wire [7:0] t_r17_c35_7;
  wire [7:0] t_r17_c35_8;
  wire [7:0] t_r17_c35_9;
  wire [7:0] t_r17_c35_10;
  wire [7:0] t_r17_c35_11;
  wire [7:0] t_r17_c35_12;
  wire [7:0] t_r17_c36_0;
  wire [7:0] t_r17_c36_1;
  wire [7:0] t_r17_c36_2;
  wire [7:0] t_r17_c36_3;
  wire [7:0] t_r17_c36_4;
  wire [7:0] t_r17_c36_5;
  wire [7:0] t_r17_c36_6;
  wire [7:0] t_r17_c36_7;
  wire [7:0] t_r17_c36_8;
  wire [7:0] t_r17_c36_9;
  wire [7:0] t_r17_c36_10;
  wire [7:0] t_r17_c36_11;
  wire [7:0] t_r17_c36_12;
  wire [7:0] t_r17_c37_0;
  wire [7:0] t_r17_c37_1;
  wire [7:0] t_r17_c37_2;
  wire [7:0] t_r17_c37_3;
  wire [7:0] t_r17_c37_4;
  wire [7:0] t_r17_c37_5;
  wire [7:0] t_r17_c37_6;
  wire [7:0] t_r17_c37_7;
  wire [7:0] t_r17_c37_8;
  wire [7:0] t_r17_c37_9;
  wire [7:0] t_r17_c37_10;
  wire [7:0] t_r17_c37_11;
  wire [7:0] t_r17_c37_12;
  wire [7:0] t_r17_c38_0;
  wire [7:0] t_r17_c38_1;
  wire [7:0] t_r17_c38_2;
  wire [7:0] t_r17_c38_3;
  wire [7:0] t_r17_c38_4;
  wire [7:0] t_r17_c38_5;
  wire [7:0] t_r17_c38_6;
  wire [7:0] t_r17_c38_7;
  wire [7:0] t_r17_c38_8;
  wire [7:0] t_r17_c38_9;
  wire [7:0] t_r17_c38_10;
  wire [7:0] t_r17_c38_11;
  wire [7:0] t_r17_c38_12;
  wire [7:0] t_r17_c39_0;
  wire [7:0] t_r17_c39_1;
  wire [7:0] t_r17_c39_2;
  wire [7:0] t_r17_c39_3;
  wire [7:0] t_r17_c39_4;
  wire [7:0] t_r17_c39_5;
  wire [7:0] t_r17_c39_6;
  wire [7:0] t_r17_c39_7;
  wire [7:0] t_r17_c39_8;
  wire [7:0] t_r17_c39_9;
  wire [7:0] t_r17_c39_10;
  wire [7:0] t_r17_c39_11;
  wire [7:0] t_r17_c39_12;
  wire [7:0] t_r17_c40_0;
  wire [7:0] t_r17_c40_1;
  wire [7:0] t_r17_c40_2;
  wire [7:0] t_r17_c40_3;
  wire [7:0] t_r17_c40_4;
  wire [7:0] t_r17_c40_5;
  wire [7:0] t_r17_c40_6;
  wire [7:0] t_r17_c40_7;
  wire [7:0] t_r17_c40_8;
  wire [7:0] t_r17_c40_9;
  wire [7:0] t_r17_c40_10;
  wire [7:0] t_r17_c40_11;
  wire [7:0] t_r17_c40_12;
  wire [7:0] t_r17_c41_0;
  wire [7:0] t_r17_c41_1;
  wire [7:0] t_r17_c41_2;
  wire [7:0] t_r17_c41_3;
  wire [7:0] t_r17_c41_4;
  wire [7:0] t_r17_c41_5;
  wire [7:0] t_r17_c41_6;
  wire [7:0] t_r17_c41_7;
  wire [7:0] t_r17_c41_8;
  wire [7:0] t_r17_c41_9;
  wire [7:0] t_r17_c41_10;
  wire [7:0] t_r17_c41_11;
  wire [7:0] t_r17_c41_12;
  wire [7:0] t_r17_c42_0;
  wire [7:0] t_r17_c42_1;
  wire [7:0] t_r17_c42_2;
  wire [7:0] t_r17_c42_3;
  wire [7:0] t_r17_c42_4;
  wire [7:0] t_r17_c42_5;
  wire [7:0] t_r17_c42_6;
  wire [7:0] t_r17_c42_7;
  wire [7:0] t_r17_c42_8;
  wire [7:0] t_r17_c42_9;
  wire [7:0] t_r17_c42_10;
  wire [7:0] t_r17_c42_11;
  wire [7:0] t_r17_c42_12;
  wire [7:0] t_r17_c43_0;
  wire [7:0] t_r17_c43_1;
  wire [7:0] t_r17_c43_2;
  wire [7:0] t_r17_c43_3;
  wire [7:0] t_r17_c43_4;
  wire [7:0] t_r17_c43_5;
  wire [7:0] t_r17_c43_6;
  wire [7:0] t_r17_c43_7;
  wire [7:0] t_r17_c43_8;
  wire [7:0] t_r17_c43_9;
  wire [7:0] t_r17_c43_10;
  wire [7:0] t_r17_c43_11;
  wire [7:0] t_r17_c43_12;
  wire [7:0] t_r17_c44_0;
  wire [7:0] t_r17_c44_1;
  wire [7:0] t_r17_c44_2;
  wire [7:0] t_r17_c44_3;
  wire [7:0] t_r17_c44_4;
  wire [7:0] t_r17_c44_5;
  wire [7:0] t_r17_c44_6;
  wire [7:0] t_r17_c44_7;
  wire [7:0] t_r17_c44_8;
  wire [7:0] t_r17_c44_9;
  wire [7:0] t_r17_c44_10;
  wire [7:0] t_r17_c44_11;
  wire [7:0] t_r17_c44_12;
  wire [7:0] t_r17_c45_0;
  wire [7:0] t_r17_c45_1;
  wire [7:0] t_r17_c45_2;
  wire [7:0] t_r17_c45_3;
  wire [7:0] t_r17_c45_4;
  wire [7:0] t_r17_c45_5;
  wire [7:0] t_r17_c45_6;
  wire [7:0] t_r17_c45_7;
  wire [7:0] t_r17_c45_8;
  wire [7:0] t_r17_c45_9;
  wire [7:0] t_r17_c45_10;
  wire [7:0] t_r17_c45_11;
  wire [7:0] t_r17_c45_12;
  wire [7:0] t_r17_c46_0;
  wire [7:0] t_r17_c46_1;
  wire [7:0] t_r17_c46_2;
  wire [7:0] t_r17_c46_3;
  wire [7:0] t_r17_c46_4;
  wire [7:0] t_r17_c46_5;
  wire [7:0] t_r17_c46_6;
  wire [7:0] t_r17_c46_7;
  wire [7:0] t_r17_c46_8;
  wire [7:0] t_r17_c46_9;
  wire [7:0] t_r17_c46_10;
  wire [7:0] t_r17_c46_11;
  wire [7:0] t_r17_c46_12;
  wire [7:0] t_r17_c47_0;
  wire [7:0] t_r17_c47_1;
  wire [7:0] t_r17_c47_2;
  wire [7:0] t_r17_c47_3;
  wire [7:0] t_r17_c47_4;
  wire [7:0] t_r17_c47_5;
  wire [7:0] t_r17_c47_6;
  wire [7:0] t_r17_c47_7;
  wire [7:0] t_r17_c47_8;
  wire [7:0] t_r17_c47_9;
  wire [7:0] t_r17_c47_10;
  wire [7:0] t_r17_c47_11;
  wire [7:0] t_r17_c47_12;
  wire [7:0] t_r17_c48_0;
  wire [7:0] t_r17_c48_1;
  wire [7:0] t_r17_c48_2;
  wire [7:0] t_r17_c48_3;
  wire [7:0] t_r17_c48_4;
  wire [7:0] t_r17_c48_5;
  wire [7:0] t_r17_c48_6;
  wire [7:0] t_r17_c48_7;
  wire [7:0] t_r17_c48_8;
  wire [7:0] t_r17_c48_9;
  wire [7:0] t_r17_c48_10;
  wire [7:0] t_r17_c48_11;
  wire [7:0] t_r17_c48_12;
  wire [7:0] t_r17_c49_0;
  wire [7:0] t_r17_c49_1;
  wire [7:0] t_r17_c49_2;
  wire [7:0] t_r17_c49_3;
  wire [7:0] t_r17_c49_4;
  wire [7:0] t_r17_c49_5;
  wire [7:0] t_r17_c49_6;
  wire [7:0] t_r17_c49_7;
  wire [7:0] t_r17_c49_8;
  wire [7:0] t_r17_c49_9;
  wire [7:0] t_r17_c49_10;
  wire [7:0] t_r17_c49_11;
  wire [7:0] t_r17_c49_12;
  wire [7:0] t_r17_c50_0;
  wire [7:0] t_r17_c50_1;
  wire [7:0] t_r17_c50_2;
  wire [7:0] t_r17_c50_3;
  wire [7:0] t_r17_c50_4;
  wire [7:0] t_r17_c50_5;
  wire [7:0] t_r17_c50_6;
  wire [7:0] t_r17_c50_7;
  wire [7:0] t_r17_c50_8;
  wire [7:0] t_r17_c50_9;
  wire [7:0] t_r17_c50_10;
  wire [7:0] t_r17_c50_11;
  wire [7:0] t_r17_c50_12;
  wire [7:0] t_r17_c51_0;
  wire [7:0] t_r17_c51_1;
  wire [7:0] t_r17_c51_2;
  wire [7:0] t_r17_c51_3;
  wire [7:0] t_r17_c51_4;
  wire [7:0] t_r17_c51_5;
  wire [7:0] t_r17_c51_6;
  wire [7:0] t_r17_c51_7;
  wire [7:0] t_r17_c51_8;
  wire [7:0] t_r17_c51_9;
  wire [7:0] t_r17_c51_10;
  wire [7:0] t_r17_c51_11;
  wire [7:0] t_r17_c51_12;
  wire [7:0] t_r17_c52_0;
  wire [7:0] t_r17_c52_1;
  wire [7:0] t_r17_c52_2;
  wire [7:0] t_r17_c52_3;
  wire [7:0] t_r17_c52_4;
  wire [7:0] t_r17_c52_5;
  wire [7:0] t_r17_c52_6;
  wire [7:0] t_r17_c52_7;
  wire [7:0] t_r17_c52_8;
  wire [7:0] t_r17_c52_9;
  wire [7:0] t_r17_c52_10;
  wire [7:0] t_r17_c52_11;
  wire [7:0] t_r17_c52_12;
  wire [7:0] t_r17_c53_0;
  wire [7:0] t_r17_c53_1;
  wire [7:0] t_r17_c53_2;
  wire [7:0] t_r17_c53_3;
  wire [7:0] t_r17_c53_4;
  wire [7:0] t_r17_c53_5;
  wire [7:0] t_r17_c53_6;
  wire [7:0] t_r17_c53_7;
  wire [7:0] t_r17_c53_8;
  wire [7:0] t_r17_c53_9;
  wire [7:0] t_r17_c53_10;
  wire [7:0] t_r17_c53_11;
  wire [7:0] t_r17_c53_12;
  wire [7:0] t_r17_c54_0;
  wire [7:0] t_r17_c54_1;
  wire [7:0] t_r17_c54_2;
  wire [7:0] t_r17_c54_3;
  wire [7:0] t_r17_c54_4;
  wire [7:0] t_r17_c54_5;
  wire [7:0] t_r17_c54_6;
  wire [7:0] t_r17_c54_7;
  wire [7:0] t_r17_c54_8;
  wire [7:0] t_r17_c54_9;
  wire [7:0] t_r17_c54_10;
  wire [7:0] t_r17_c54_11;
  wire [7:0] t_r17_c54_12;
  wire [7:0] t_r17_c55_0;
  wire [7:0] t_r17_c55_1;
  wire [7:0] t_r17_c55_2;
  wire [7:0] t_r17_c55_3;
  wire [7:0] t_r17_c55_4;
  wire [7:0] t_r17_c55_5;
  wire [7:0] t_r17_c55_6;
  wire [7:0] t_r17_c55_7;
  wire [7:0] t_r17_c55_8;
  wire [7:0] t_r17_c55_9;
  wire [7:0] t_r17_c55_10;
  wire [7:0] t_r17_c55_11;
  wire [7:0] t_r17_c55_12;
  wire [7:0] t_r17_c56_0;
  wire [7:0] t_r17_c56_1;
  wire [7:0] t_r17_c56_2;
  wire [7:0] t_r17_c56_3;
  wire [7:0] t_r17_c56_4;
  wire [7:0] t_r17_c56_5;
  wire [7:0] t_r17_c56_6;
  wire [7:0] t_r17_c56_7;
  wire [7:0] t_r17_c56_8;
  wire [7:0] t_r17_c56_9;
  wire [7:0] t_r17_c56_10;
  wire [7:0] t_r17_c56_11;
  wire [7:0] t_r17_c56_12;
  wire [7:0] t_r17_c57_0;
  wire [7:0] t_r17_c57_1;
  wire [7:0] t_r17_c57_2;
  wire [7:0] t_r17_c57_3;
  wire [7:0] t_r17_c57_4;
  wire [7:0] t_r17_c57_5;
  wire [7:0] t_r17_c57_6;
  wire [7:0] t_r17_c57_7;
  wire [7:0] t_r17_c57_8;
  wire [7:0] t_r17_c57_9;
  wire [7:0] t_r17_c57_10;
  wire [7:0] t_r17_c57_11;
  wire [7:0] t_r17_c57_12;
  wire [7:0] t_r17_c58_0;
  wire [7:0] t_r17_c58_1;
  wire [7:0] t_r17_c58_2;
  wire [7:0] t_r17_c58_3;
  wire [7:0] t_r17_c58_4;
  wire [7:0] t_r17_c58_5;
  wire [7:0] t_r17_c58_6;
  wire [7:0] t_r17_c58_7;
  wire [7:0] t_r17_c58_8;
  wire [7:0] t_r17_c58_9;
  wire [7:0] t_r17_c58_10;
  wire [7:0] t_r17_c58_11;
  wire [7:0] t_r17_c58_12;
  wire [7:0] t_r17_c59_0;
  wire [7:0] t_r17_c59_1;
  wire [7:0] t_r17_c59_2;
  wire [7:0] t_r17_c59_3;
  wire [7:0] t_r17_c59_4;
  wire [7:0] t_r17_c59_5;
  wire [7:0] t_r17_c59_6;
  wire [7:0] t_r17_c59_7;
  wire [7:0] t_r17_c59_8;
  wire [7:0] t_r17_c59_9;
  wire [7:0] t_r17_c59_10;
  wire [7:0] t_r17_c59_11;
  wire [7:0] t_r17_c59_12;
  wire [7:0] t_r17_c60_0;
  wire [7:0] t_r17_c60_1;
  wire [7:0] t_r17_c60_2;
  wire [7:0] t_r17_c60_3;
  wire [7:0] t_r17_c60_4;
  wire [7:0] t_r17_c60_5;
  wire [7:0] t_r17_c60_6;
  wire [7:0] t_r17_c60_7;
  wire [7:0] t_r17_c60_8;
  wire [7:0] t_r17_c60_9;
  wire [7:0] t_r17_c60_10;
  wire [7:0] t_r17_c60_11;
  wire [7:0] t_r17_c60_12;
  wire [7:0] t_r17_c61_0;
  wire [7:0] t_r17_c61_1;
  wire [7:0] t_r17_c61_2;
  wire [7:0] t_r17_c61_3;
  wire [7:0] t_r17_c61_4;
  wire [7:0] t_r17_c61_5;
  wire [7:0] t_r17_c61_6;
  wire [7:0] t_r17_c61_7;
  wire [7:0] t_r17_c61_8;
  wire [7:0] t_r17_c61_9;
  wire [7:0] t_r17_c61_10;
  wire [7:0] t_r17_c61_11;
  wire [7:0] t_r17_c61_12;
  wire [7:0] t_r17_c62_0;
  wire [7:0] t_r17_c62_1;
  wire [7:0] t_r17_c62_2;
  wire [7:0] t_r17_c62_3;
  wire [7:0] t_r17_c62_4;
  wire [7:0] t_r17_c62_5;
  wire [7:0] t_r17_c62_6;
  wire [7:0] t_r17_c62_7;
  wire [7:0] t_r17_c62_8;
  wire [7:0] t_r17_c62_9;
  wire [7:0] t_r17_c62_10;
  wire [7:0] t_r17_c62_11;
  wire [7:0] t_r17_c62_12;
  wire [7:0] t_r17_c63_0;
  wire [7:0] t_r17_c63_1;
  wire [7:0] t_r17_c63_2;
  wire [7:0] t_r17_c63_3;
  wire [7:0] t_r17_c63_4;
  wire [7:0] t_r17_c63_5;
  wire [7:0] t_r17_c63_6;
  wire [7:0] t_r17_c63_7;
  wire [7:0] t_r17_c63_8;
  wire [7:0] t_r17_c63_9;
  wire [7:0] t_r17_c63_10;
  wire [7:0] t_r17_c63_11;
  wire [7:0] t_r17_c63_12;
  wire [7:0] t_r17_c64_0;
  wire [7:0] t_r17_c64_1;
  wire [7:0] t_r17_c64_2;
  wire [7:0] t_r17_c64_3;
  wire [7:0] t_r17_c64_4;
  wire [7:0] t_r17_c64_5;
  wire [7:0] t_r17_c64_6;
  wire [7:0] t_r17_c64_7;
  wire [7:0] t_r17_c64_8;
  wire [7:0] t_r17_c64_9;
  wire [7:0] t_r17_c64_10;
  wire [7:0] t_r17_c64_11;
  wire [7:0] t_r17_c64_12;
  wire [7:0] t_r17_c65_0;
  wire [7:0] t_r17_c65_1;
  wire [7:0] t_r17_c65_2;
  wire [7:0] t_r17_c65_3;
  wire [7:0] t_r17_c65_4;
  wire [7:0] t_r17_c65_5;
  wire [7:0] t_r17_c65_6;
  wire [7:0] t_r17_c65_7;
  wire [7:0] t_r17_c65_8;
  wire [7:0] t_r17_c65_9;
  wire [7:0] t_r17_c65_10;
  wire [7:0] t_r17_c65_11;
  wire [7:0] t_r17_c65_12;
  wire [7:0] t_r18_c0_0;
  wire [7:0] t_r18_c0_1;
  wire [7:0] t_r18_c0_2;
  wire [7:0] t_r18_c0_3;
  wire [7:0] t_r18_c0_4;
  wire [7:0] t_r18_c0_5;
  wire [7:0] t_r18_c0_6;
  wire [7:0] t_r18_c0_7;
  wire [7:0] t_r18_c0_8;
  wire [7:0] t_r18_c0_9;
  wire [7:0] t_r18_c0_10;
  wire [7:0] t_r18_c0_11;
  wire [7:0] t_r18_c0_12;
  wire [7:0] t_r18_c1_0;
  wire [7:0] t_r18_c1_1;
  wire [7:0] t_r18_c1_2;
  wire [7:0] t_r18_c1_3;
  wire [7:0] t_r18_c1_4;
  wire [7:0] t_r18_c1_5;
  wire [7:0] t_r18_c1_6;
  wire [7:0] t_r18_c1_7;
  wire [7:0] t_r18_c1_8;
  wire [7:0] t_r18_c1_9;
  wire [7:0] t_r18_c1_10;
  wire [7:0] t_r18_c1_11;
  wire [7:0] t_r18_c1_12;
  wire [7:0] t_r18_c2_0;
  wire [7:0] t_r18_c2_1;
  wire [7:0] t_r18_c2_2;
  wire [7:0] t_r18_c2_3;
  wire [7:0] t_r18_c2_4;
  wire [7:0] t_r18_c2_5;
  wire [7:0] t_r18_c2_6;
  wire [7:0] t_r18_c2_7;
  wire [7:0] t_r18_c2_8;
  wire [7:0] t_r18_c2_9;
  wire [7:0] t_r18_c2_10;
  wire [7:0] t_r18_c2_11;
  wire [7:0] t_r18_c2_12;
  wire [7:0] t_r18_c3_0;
  wire [7:0] t_r18_c3_1;
  wire [7:0] t_r18_c3_2;
  wire [7:0] t_r18_c3_3;
  wire [7:0] t_r18_c3_4;
  wire [7:0] t_r18_c3_5;
  wire [7:0] t_r18_c3_6;
  wire [7:0] t_r18_c3_7;
  wire [7:0] t_r18_c3_8;
  wire [7:0] t_r18_c3_9;
  wire [7:0] t_r18_c3_10;
  wire [7:0] t_r18_c3_11;
  wire [7:0] t_r18_c3_12;
  wire [7:0] t_r18_c4_0;
  wire [7:0] t_r18_c4_1;
  wire [7:0] t_r18_c4_2;
  wire [7:0] t_r18_c4_3;
  wire [7:0] t_r18_c4_4;
  wire [7:0] t_r18_c4_5;
  wire [7:0] t_r18_c4_6;
  wire [7:0] t_r18_c4_7;
  wire [7:0] t_r18_c4_8;
  wire [7:0] t_r18_c4_9;
  wire [7:0] t_r18_c4_10;
  wire [7:0] t_r18_c4_11;
  wire [7:0] t_r18_c4_12;
  wire [7:0] t_r18_c5_0;
  wire [7:0] t_r18_c5_1;
  wire [7:0] t_r18_c5_2;
  wire [7:0] t_r18_c5_3;
  wire [7:0] t_r18_c5_4;
  wire [7:0] t_r18_c5_5;
  wire [7:0] t_r18_c5_6;
  wire [7:0] t_r18_c5_7;
  wire [7:0] t_r18_c5_8;
  wire [7:0] t_r18_c5_9;
  wire [7:0] t_r18_c5_10;
  wire [7:0] t_r18_c5_11;
  wire [7:0] t_r18_c5_12;
  wire [7:0] t_r18_c6_0;
  wire [7:0] t_r18_c6_1;
  wire [7:0] t_r18_c6_2;
  wire [7:0] t_r18_c6_3;
  wire [7:0] t_r18_c6_4;
  wire [7:0] t_r18_c6_5;
  wire [7:0] t_r18_c6_6;
  wire [7:0] t_r18_c6_7;
  wire [7:0] t_r18_c6_8;
  wire [7:0] t_r18_c6_9;
  wire [7:0] t_r18_c6_10;
  wire [7:0] t_r18_c6_11;
  wire [7:0] t_r18_c6_12;
  wire [7:0] t_r18_c7_0;
  wire [7:0] t_r18_c7_1;
  wire [7:0] t_r18_c7_2;
  wire [7:0] t_r18_c7_3;
  wire [7:0] t_r18_c7_4;
  wire [7:0] t_r18_c7_5;
  wire [7:0] t_r18_c7_6;
  wire [7:0] t_r18_c7_7;
  wire [7:0] t_r18_c7_8;
  wire [7:0] t_r18_c7_9;
  wire [7:0] t_r18_c7_10;
  wire [7:0] t_r18_c7_11;
  wire [7:0] t_r18_c7_12;
  wire [7:0] t_r18_c8_0;
  wire [7:0] t_r18_c8_1;
  wire [7:0] t_r18_c8_2;
  wire [7:0] t_r18_c8_3;
  wire [7:0] t_r18_c8_4;
  wire [7:0] t_r18_c8_5;
  wire [7:0] t_r18_c8_6;
  wire [7:0] t_r18_c8_7;
  wire [7:0] t_r18_c8_8;
  wire [7:0] t_r18_c8_9;
  wire [7:0] t_r18_c8_10;
  wire [7:0] t_r18_c8_11;
  wire [7:0] t_r18_c8_12;
  wire [7:0] t_r18_c9_0;
  wire [7:0] t_r18_c9_1;
  wire [7:0] t_r18_c9_2;
  wire [7:0] t_r18_c9_3;
  wire [7:0] t_r18_c9_4;
  wire [7:0] t_r18_c9_5;
  wire [7:0] t_r18_c9_6;
  wire [7:0] t_r18_c9_7;
  wire [7:0] t_r18_c9_8;
  wire [7:0] t_r18_c9_9;
  wire [7:0] t_r18_c9_10;
  wire [7:0] t_r18_c9_11;
  wire [7:0] t_r18_c9_12;
  wire [7:0] t_r18_c10_0;
  wire [7:0] t_r18_c10_1;
  wire [7:0] t_r18_c10_2;
  wire [7:0] t_r18_c10_3;
  wire [7:0] t_r18_c10_4;
  wire [7:0] t_r18_c10_5;
  wire [7:0] t_r18_c10_6;
  wire [7:0] t_r18_c10_7;
  wire [7:0] t_r18_c10_8;
  wire [7:0] t_r18_c10_9;
  wire [7:0] t_r18_c10_10;
  wire [7:0] t_r18_c10_11;
  wire [7:0] t_r18_c10_12;
  wire [7:0] t_r18_c11_0;
  wire [7:0] t_r18_c11_1;
  wire [7:0] t_r18_c11_2;
  wire [7:0] t_r18_c11_3;
  wire [7:0] t_r18_c11_4;
  wire [7:0] t_r18_c11_5;
  wire [7:0] t_r18_c11_6;
  wire [7:0] t_r18_c11_7;
  wire [7:0] t_r18_c11_8;
  wire [7:0] t_r18_c11_9;
  wire [7:0] t_r18_c11_10;
  wire [7:0] t_r18_c11_11;
  wire [7:0] t_r18_c11_12;
  wire [7:0] t_r18_c12_0;
  wire [7:0] t_r18_c12_1;
  wire [7:0] t_r18_c12_2;
  wire [7:0] t_r18_c12_3;
  wire [7:0] t_r18_c12_4;
  wire [7:0] t_r18_c12_5;
  wire [7:0] t_r18_c12_6;
  wire [7:0] t_r18_c12_7;
  wire [7:0] t_r18_c12_8;
  wire [7:0] t_r18_c12_9;
  wire [7:0] t_r18_c12_10;
  wire [7:0] t_r18_c12_11;
  wire [7:0] t_r18_c12_12;
  wire [7:0] t_r18_c13_0;
  wire [7:0] t_r18_c13_1;
  wire [7:0] t_r18_c13_2;
  wire [7:0] t_r18_c13_3;
  wire [7:0] t_r18_c13_4;
  wire [7:0] t_r18_c13_5;
  wire [7:0] t_r18_c13_6;
  wire [7:0] t_r18_c13_7;
  wire [7:0] t_r18_c13_8;
  wire [7:0] t_r18_c13_9;
  wire [7:0] t_r18_c13_10;
  wire [7:0] t_r18_c13_11;
  wire [7:0] t_r18_c13_12;
  wire [7:0] t_r18_c14_0;
  wire [7:0] t_r18_c14_1;
  wire [7:0] t_r18_c14_2;
  wire [7:0] t_r18_c14_3;
  wire [7:0] t_r18_c14_4;
  wire [7:0] t_r18_c14_5;
  wire [7:0] t_r18_c14_6;
  wire [7:0] t_r18_c14_7;
  wire [7:0] t_r18_c14_8;
  wire [7:0] t_r18_c14_9;
  wire [7:0] t_r18_c14_10;
  wire [7:0] t_r18_c14_11;
  wire [7:0] t_r18_c14_12;
  wire [7:0] t_r18_c15_0;
  wire [7:0] t_r18_c15_1;
  wire [7:0] t_r18_c15_2;
  wire [7:0] t_r18_c15_3;
  wire [7:0] t_r18_c15_4;
  wire [7:0] t_r18_c15_5;
  wire [7:0] t_r18_c15_6;
  wire [7:0] t_r18_c15_7;
  wire [7:0] t_r18_c15_8;
  wire [7:0] t_r18_c15_9;
  wire [7:0] t_r18_c15_10;
  wire [7:0] t_r18_c15_11;
  wire [7:0] t_r18_c15_12;
  wire [7:0] t_r18_c16_0;
  wire [7:0] t_r18_c16_1;
  wire [7:0] t_r18_c16_2;
  wire [7:0] t_r18_c16_3;
  wire [7:0] t_r18_c16_4;
  wire [7:0] t_r18_c16_5;
  wire [7:0] t_r18_c16_6;
  wire [7:0] t_r18_c16_7;
  wire [7:0] t_r18_c16_8;
  wire [7:0] t_r18_c16_9;
  wire [7:0] t_r18_c16_10;
  wire [7:0] t_r18_c16_11;
  wire [7:0] t_r18_c16_12;
  wire [7:0] t_r18_c17_0;
  wire [7:0] t_r18_c17_1;
  wire [7:0] t_r18_c17_2;
  wire [7:0] t_r18_c17_3;
  wire [7:0] t_r18_c17_4;
  wire [7:0] t_r18_c17_5;
  wire [7:0] t_r18_c17_6;
  wire [7:0] t_r18_c17_7;
  wire [7:0] t_r18_c17_8;
  wire [7:0] t_r18_c17_9;
  wire [7:0] t_r18_c17_10;
  wire [7:0] t_r18_c17_11;
  wire [7:0] t_r18_c17_12;
  wire [7:0] t_r18_c18_0;
  wire [7:0] t_r18_c18_1;
  wire [7:0] t_r18_c18_2;
  wire [7:0] t_r18_c18_3;
  wire [7:0] t_r18_c18_4;
  wire [7:0] t_r18_c18_5;
  wire [7:0] t_r18_c18_6;
  wire [7:0] t_r18_c18_7;
  wire [7:0] t_r18_c18_8;
  wire [7:0] t_r18_c18_9;
  wire [7:0] t_r18_c18_10;
  wire [7:0] t_r18_c18_11;
  wire [7:0] t_r18_c18_12;
  wire [7:0] t_r18_c19_0;
  wire [7:0] t_r18_c19_1;
  wire [7:0] t_r18_c19_2;
  wire [7:0] t_r18_c19_3;
  wire [7:0] t_r18_c19_4;
  wire [7:0] t_r18_c19_5;
  wire [7:0] t_r18_c19_6;
  wire [7:0] t_r18_c19_7;
  wire [7:0] t_r18_c19_8;
  wire [7:0] t_r18_c19_9;
  wire [7:0] t_r18_c19_10;
  wire [7:0] t_r18_c19_11;
  wire [7:0] t_r18_c19_12;
  wire [7:0] t_r18_c20_0;
  wire [7:0] t_r18_c20_1;
  wire [7:0] t_r18_c20_2;
  wire [7:0] t_r18_c20_3;
  wire [7:0] t_r18_c20_4;
  wire [7:0] t_r18_c20_5;
  wire [7:0] t_r18_c20_6;
  wire [7:0] t_r18_c20_7;
  wire [7:0] t_r18_c20_8;
  wire [7:0] t_r18_c20_9;
  wire [7:0] t_r18_c20_10;
  wire [7:0] t_r18_c20_11;
  wire [7:0] t_r18_c20_12;
  wire [7:0] t_r18_c21_0;
  wire [7:0] t_r18_c21_1;
  wire [7:0] t_r18_c21_2;
  wire [7:0] t_r18_c21_3;
  wire [7:0] t_r18_c21_4;
  wire [7:0] t_r18_c21_5;
  wire [7:0] t_r18_c21_6;
  wire [7:0] t_r18_c21_7;
  wire [7:0] t_r18_c21_8;
  wire [7:0] t_r18_c21_9;
  wire [7:0] t_r18_c21_10;
  wire [7:0] t_r18_c21_11;
  wire [7:0] t_r18_c21_12;
  wire [7:0] t_r18_c22_0;
  wire [7:0] t_r18_c22_1;
  wire [7:0] t_r18_c22_2;
  wire [7:0] t_r18_c22_3;
  wire [7:0] t_r18_c22_4;
  wire [7:0] t_r18_c22_5;
  wire [7:0] t_r18_c22_6;
  wire [7:0] t_r18_c22_7;
  wire [7:0] t_r18_c22_8;
  wire [7:0] t_r18_c22_9;
  wire [7:0] t_r18_c22_10;
  wire [7:0] t_r18_c22_11;
  wire [7:0] t_r18_c22_12;
  wire [7:0] t_r18_c23_0;
  wire [7:0] t_r18_c23_1;
  wire [7:0] t_r18_c23_2;
  wire [7:0] t_r18_c23_3;
  wire [7:0] t_r18_c23_4;
  wire [7:0] t_r18_c23_5;
  wire [7:0] t_r18_c23_6;
  wire [7:0] t_r18_c23_7;
  wire [7:0] t_r18_c23_8;
  wire [7:0] t_r18_c23_9;
  wire [7:0] t_r18_c23_10;
  wire [7:0] t_r18_c23_11;
  wire [7:0] t_r18_c23_12;
  wire [7:0] t_r18_c24_0;
  wire [7:0] t_r18_c24_1;
  wire [7:0] t_r18_c24_2;
  wire [7:0] t_r18_c24_3;
  wire [7:0] t_r18_c24_4;
  wire [7:0] t_r18_c24_5;
  wire [7:0] t_r18_c24_6;
  wire [7:0] t_r18_c24_7;
  wire [7:0] t_r18_c24_8;
  wire [7:0] t_r18_c24_9;
  wire [7:0] t_r18_c24_10;
  wire [7:0] t_r18_c24_11;
  wire [7:0] t_r18_c24_12;
  wire [7:0] t_r18_c25_0;
  wire [7:0] t_r18_c25_1;
  wire [7:0] t_r18_c25_2;
  wire [7:0] t_r18_c25_3;
  wire [7:0] t_r18_c25_4;
  wire [7:0] t_r18_c25_5;
  wire [7:0] t_r18_c25_6;
  wire [7:0] t_r18_c25_7;
  wire [7:0] t_r18_c25_8;
  wire [7:0] t_r18_c25_9;
  wire [7:0] t_r18_c25_10;
  wire [7:0] t_r18_c25_11;
  wire [7:0] t_r18_c25_12;
  wire [7:0] t_r18_c26_0;
  wire [7:0] t_r18_c26_1;
  wire [7:0] t_r18_c26_2;
  wire [7:0] t_r18_c26_3;
  wire [7:0] t_r18_c26_4;
  wire [7:0] t_r18_c26_5;
  wire [7:0] t_r18_c26_6;
  wire [7:0] t_r18_c26_7;
  wire [7:0] t_r18_c26_8;
  wire [7:0] t_r18_c26_9;
  wire [7:0] t_r18_c26_10;
  wire [7:0] t_r18_c26_11;
  wire [7:0] t_r18_c26_12;
  wire [7:0] t_r18_c27_0;
  wire [7:0] t_r18_c27_1;
  wire [7:0] t_r18_c27_2;
  wire [7:0] t_r18_c27_3;
  wire [7:0] t_r18_c27_4;
  wire [7:0] t_r18_c27_5;
  wire [7:0] t_r18_c27_6;
  wire [7:0] t_r18_c27_7;
  wire [7:0] t_r18_c27_8;
  wire [7:0] t_r18_c27_9;
  wire [7:0] t_r18_c27_10;
  wire [7:0] t_r18_c27_11;
  wire [7:0] t_r18_c27_12;
  wire [7:0] t_r18_c28_0;
  wire [7:0] t_r18_c28_1;
  wire [7:0] t_r18_c28_2;
  wire [7:0] t_r18_c28_3;
  wire [7:0] t_r18_c28_4;
  wire [7:0] t_r18_c28_5;
  wire [7:0] t_r18_c28_6;
  wire [7:0] t_r18_c28_7;
  wire [7:0] t_r18_c28_8;
  wire [7:0] t_r18_c28_9;
  wire [7:0] t_r18_c28_10;
  wire [7:0] t_r18_c28_11;
  wire [7:0] t_r18_c28_12;
  wire [7:0] t_r18_c29_0;
  wire [7:0] t_r18_c29_1;
  wire [7:0] t_r18_c29_2;
  wire [7:0] t_r18_c29_3;
  wire [7:0] t_r18_c29_4;
  wire [7:0] t_r18_c29_5;
  wire [7:0] t_r18_c29_6;
  wire [7:0] t_r18_c29_7;
  wire [7:0] t_r18_c29_8;
  wire [7:0] t_r18_c29_9;
  wire [7:0] t_r18_c29_10;
  wire [7:0] t_r18_c29_11;
  wire [7:0] t_r18_c29_12;
  wire [7:0] t_r18_c30_0;
  wire [7:0] t_r18_c30_1;
  wire [7:0] t_r18_c30_2;
  wire [7:0] t_r18_c30_3;
  wire [7:0] t_r18_c30_4;
  wire [7:0] t_r18_c30_5;
  wire [7:0] t_r18_c30_6;
  wire [7:0] t_r18_c30_7;
  wire [7:0] t_r18_c30_8;
  wire [7:0] t_r18_c30_9;
  wire [7:0] t_r18_c30_10;
  wire [7:0] t_r18_c30_11;
  wire [7:0] t_r18_c30_12;
  wire [7:0] t_r18_c31_0;
  wire [7:0] t_r18_c31_1;
  wire [7:0] t_r18_c31_2;
  wire [7:0] t_r18_c31_3;
  wire [7:0] t_r18_c31_4;
  wire [7:0] t_r18_c31_5;
  wire [7:0] t_r18_c31_6;
  wire [7:0] t_r18_c31_7;
  wire [7:0] t_r18_c31_8;
  wire [7:0] t_r18_c31_9;
  wire [7:0] t_r18_c31_10;
  wire [7:0] t_r18_c31_11;
  wire [7:0] t_r18_c31_12;
  wire [7:0] t_r18_c32_0;
  wire [7:0] t_r18_c32_1;
  wire [7:0] t_r18_c32_2;
  wire [7:0] t_r18_c32_3;
  wire [7:0] t_r18_c32_4;
  wire [7:0] t_r18_c32_5;
  wire [7:0] t_r18_c32_6;
  wire [7:0] t_r18_c32_7;
  wire [7:0] t_r18_c32_8;
  wire [7:0] t_r18_c32_9;
  wire [7:0] t_r18_c32_10;
  wire [7:0] t_r18_c32_11;
  wire [7:0] t_r18_c32_12;
  wire [7:0] t_r18_c33_0;
  wire [7:0] t_r18_c33_1;
  wire [7:0] t_r18_c33_2;
  wire [7:0] t_r18_c33_3;
  wire [7:0] t_r18_c33_4;
  wire [7:0] t_r18_c33_5;
  wire [7:0] t_r18_c33_6;
  wire [7:0] t_r18_c33_7;
  wire [7:0] t_r18_c33_8;
  wire [7:0] t_r18_c33_9;
  wire [7:0] t_r18_c33_10;
  wire [7:0] t_r18_c33_11;
  wire [7:0] t_r18_c33_12;
  wire [7:0] t_r18_c34_0;
  wire [7:0] t_r18_c34_1;
  wire [7:0] t_r18_c34_2;
  wire [7:0] t_r18_c34_3;
  wire [7:0] t_r18_c34_4;
  wire [7:0] t_r18_c34_5;
  wire [7:0] t_r18_c34_6;
  wire [7:0] t_r18_c34_7;
  wire [7:0] t_r18_c34_8;
  wire [7:0] t_r18_c34_9;
  wire [7:0] t_r18_c34_10;
  wire [7:0] t_r18_c34_11;
  wire [7:0] t_r18_c34_12;
  wire [7:0] t_r18_c35_0;
  wire [7:0] t_r18_c35_1;
  wire [7:0] t_r18_c35_2;
  wire [7:0] t_r18_c35_3;
  wire [7:0] t_r18_c35_4;
  wire [7:0] t_r18_c35_5;
  wire [7:0] t_r18_c35_6;
  wire [7:0] t_r18_c35_7;
  wire [7:0] t_r18_c35_8;
  wire [7:0] t_r18_c35_9;
  wire [7:0] t_r18_c35_10;
  wire [7:0] t_r18_c35_11;
  wire [7:0] t_r18_c35_12;
  wire [7:0] t_r18_c36_0;
  wire [7:0] t_r18_c36_1;
  wire [7:0] t_r18_c36_2;
  wire [7:0] t_r18_c36_3;
  wire [7:0] t_r18_c36_4;
  wire [7:0] t_r18_c36_5;
  wire [7:0] t_r18_c36_6;
  wire [7:0] t_r18_c36_7;
  wire [7:0] t_r18_c36_8;
  wire [7:0] t_r18_c36_9;
  wire [7:0] t_r18_c36_10;
  wire [7:0] t_r18_c36_11;
  wire [7:0] t_r18_c36_12;
  wire [7:0] t_r18_c37_0;
  wire [7:0] t_r18_c37_1;
  wire [7:0] t_r18_c37_2;
  wire [7:0] t_r18_c37_3;
  wire [7:0] t_r18_c37_4;
  wire [7:0] t_r18_c37_5;
  wire [7:0] t_r18_c37_6;
  wire [7:0] t_r18_c37_7;
  wire [7:0] t_r18_c37_8;
  wire [7:0] t_r18_c37_9;
  wire [7:0] t_r18_c37_10;
  wire [7:0] t_r18_c37_11;
  wire [7:0] t_r18_c37_12;
  wire [7:0] t_r18_c38_0;
  wire [7:0] t_r18_c38_1;
  wire [7:0] t_r18_c38_2;
  wire [7:0] t_r18_c38_3;
  wire [7:0] t_r18_c38_4;
  wire [7:0] t_r18_c38_5;
  wire [7:0] t_r18_c38_6;
  wire [7:0] t_r18_c38_7;
  wire [7:0] t_r18_c38_8;
  wire [7:0] t_r18_c38_9;
  wire [7:0] t_r18_c38_10;
  wire [7:0] t_r18_c38_11;
  wire [7:0] t_r18_c38_12;
  wire [7:0] t_r18_c39_0;
  wire [7:0] t_r18_c39_1;
  wire [7:0] t_r18_c39_2;
  wire [7:0] t_r18_c39_3;
  wire [7:0] t_r18_c39_4;
  wire [7:0] t_r18_c39_5;
  wire [7:0] t_r18_c39_6;
  wire [7:0] t_r18_c39_7;
  wire [7:0] t_r18_c39_8;
  wire [7:0] t_r18_c39_9;
  wire [7:0] t_r18_c39_10;
  wire [7:0] t_r18_c39_11;
  wire [7:0] t_r18_c39_12;
  wire [7:0] t_r18_c40_0;
  wire [7:0] t_r18_c40_1;
  wire [7:0] t_r18_c40_2;
  wire [7:0] t_r18_c40_3;
  wire [7:0] t_r18_c40_4;
  wire [7:0] t_r18_c40_5;
  wire [7:0] t_r18_c40_6;
  wire [7:0] t_r18_c40_7;
  wire [7:0] t_r18_c40_8;
  wire [7:0] t_r18_c40_9;
  wire [7:0] t_r18_c40_10;
  wire [7:0] t_r18_c40_11;
  wire [7:0] t_r18_c40_12;
  wire [7:0] t_r18_c41_0;
  wire [7:0] t_r18_c41_1;
  wire [7:0] t_r18_c41_2;
  wire [7:0] t_r18_c41_3;
  wire [7:0] t_r18_c41_4;
  wire [7:0] t_r18_c41_5;
  wire [7:0] t_r18_c41_6;
  wire [7:0] t_r18_c41_7;
  wire [7:0] t_r18_c41_8;
  wire [7:0] t_r18_c41_9;
  wire [7:0] t_r18_c41_10;
  wire [7:0] t_r18_c41_11;
  wire [7:0] t_r18_c41_12;
  wire [7:0] t_r18_c42_0;
  wire [7:0] t_r18_c42_1;
  wire [7:0] t_r18_c42_2;
  wire [7:0] t_r18_c42_3;
  wire [7:0] t_r18_c42_4;
  wire [7:0] t_r18_c42_5;
  wire [7:0] t_r18_c42_6;
  wire [7:0] t_r18_c42_7;
  wire [7:0] t_r18_c42_8;
  wire [7:0] t_r18_c42_9;
  wire [7:0] t_r18_c42_10;
  wire [7:0] t_r18_c42_11;
  wire [7:0] t_r18_c42_12;
  wire [7:0] t_r18_c43_0;
  wire [7:0] t_r18_c43_1;
  wire [7:0] t_r18_c43_2;
  wire [7:0] t_r18_c43_3;
  wire [7:0] t_r18_c43_4;
  wire [7:0] t_r18_c43_5;
  wire [7:0] t_r18_c43_6;
  wire [7:0] t_r18_c43_7;
  wire [7:0] t_r18_c43_8;
  wire [7:0] t_r18_c43_9;
  wire [7:0] t_r18_c43_10;
  wire [7:0] t_r18_c43_11;
  wire [7:0] t_r18_c43_12;
  wire [7:0] t_r18_c44_0;
  wire [7:0] t_r18_c44_1;
  wire [7:0] t_r18_c44_2;
  wire [7:0] t_r18_c44_3;
  wire [7:0] t_r18_c44_4;
  wire [7:0] t_r18_c44_5;
  wire [7:0] t_r18_c44_6;
  wire [7:0] t_r18_c44_7;
  wire [7:0] t_r18_c44_8;
  wire [7:0] t_r18_c44_9;
  wire [7:0] t_r18_c44_10;
  wire [7:0] t_r18_c44_11;
  wire [7:0] t_r18_c44_12;
  wire [7:0] t_r18_c45_0;
  wire [7:0] t_r18_c45_1;
  wire [7:0] t_r18_c45_2;
  wire [7:0] t_r18_c45_3;
  wire [7:0] t_r18_c45_4;
  wire [7:0] t_r18_c45_5;
  wire [7:0] t_r18_c45_6;
  wire [7:0] t_r18_c45_7;
  wire [7:0] t_r18_c45_8;
  wire [7:0] t_r18_c45_9;
  wire [7:0] t_r18_c45_10;
  wire [7:0] t_r18_c45_11;
  wire [7:0] t_r18_c45_12;
  wire [7:0] t_r18_c46_0;
  wire [7:0] t_r18_c46_1;
  wire [7:0] t_r18_c46_2;
  wire [7:0] t_r18_c46_3;
  wire [7:0] t_r18_c46_4;
  wire [7:0] t_r18_c46_5;
  wire [7:0] t_r18_c46_6;
  wire [7:0] t_r18_c46_7;
  wire [7:0] t_r18_c46_8;
  wire [7:0] t_r18_c46_9;
  wire [7:0] t_r18_c46_10;
  wire [7:0] t_r18_c46_11;
  wire [7:0] t_r18_c46_12;
  wire [7:0] t_r18_c47_0;
  wire [7:0] t_r18_c47_1;
  wire [7:0] t_r18_c47_2;
  wire [7:0] t_r18_c47_3;
  wire [7:0] t_r18_c47_4;
  wire [7:0] t_r18_c47_5;
  wire [7:0] t_r18_c47_6;
  wire [7:0] t_r18_c47_7;
  wire [7:0] t_r18_c47_8;
  wire [7:0] t_r18_c47_9;
  wire [7:0] t_r18_c47_10;
  wire [7:0] t_r18_c47_11;
  wire [7:0] t_r18_c47_12;
  wire [7:0] t_r18_c48_0;
  wire [7:0] t_r18_c48_1;
  wire [7:0] t_r18_c48_2;
  wire [7:0] t_r18_c48_3;
  wire [7:0] t_r18_c48_4;
  wire [7:0] t_r18_c48_5;
  wire [7:0] t_r18_c48_6;
  wire [7:0] t_r18_c48_7;
  wire [7:0] t_r18_c48_8;
  wire [7:0] t_r18_c48_9;
  wire [7:0] t_r18_c48_10;
  wire [7:0] t_r18_c48_11;
  wire [7:0] t_r18_c48_12;
  wire [7:0] t_r18_c49_0;
  wire [7:0] t_r18_c49_1;
  wire [7:0] t_r18_c49_2;
  wire [7:0] t_r18_c49_3;
  wire [7:0] t_r18_c49_4;
  wire [7:0] t_r18_c49_5;
  wire [7:0] t_r18_c49_6;
  wire [7:0] t_r18_c49_7;
  wire [7:0] t_r18_c49_8;
  wire [7:0] t_r18_c49_9;
  wire [7:0] t_r18_c49_10;
  wire [7:0] t_r18_c49_11;
  wire [7:0] t_r18_c49_12;
  wire [7:0] t_r18_c50_0;
  wire [7:0] t_r18_c50_1;
  wire [7:0] t_r18_c50_2;
  wire [7:0] t_r18_c50_3;
  wire [7:0] t_r18_c50_4;
  wire [7:0] t_r18_c50_5;
  wire [7:0] t_r18_c50_6;
  wire [7:0] t_r18_c50_7;
  wire [7:0] t_r18_c50_8;
  wire [7:0] t_r18_c50_9;
  wire [7:0] t_r18_c50_10;
  wire [7:0] t_r18_c50_11;
  wire [7:0] t_r18_c50_12;
  wire [7:0] t_r18_c51_0;
  wire [7:0] t_r18_c51_1;
  wire [7:0] t_r18_c51_2;
  wire [7:0] t_r18_c51_3;
  wire [7:0] t_r18_c51_4;
  wire [7:0] t_r18_c51_5;
  wire [7:0] t_r18_c51_6;
  wire [7:0] t_r18_c51_7;
  wire [7:0] t_r18_c51_8;
  wire [7:0] t_r18_c51_9;
  wire [7:0] t_r18_c51_10;
  wire [7:0] t_r18_c51_11;
  wire [7:0] t_r18_c51_12;
  wire [7:0] t_r18_c52_0;
  wire [7:0] t_r18_c52_1;
  wire [7:0] t_r18_c52_2;
  wire [7:0] t_r18_c52_3;
  wire [7:0] t_r18_c52_4;
  wire [7:0] t_r18_c52_5;
  wire [7:0] t_r18_c52_6;
  wire [7:0] t_r18_c52_7;
  wire [7:0] t_r18_c52_8;
  wire [7:0] t_r18_c52_9;
  wire [7:0] t_r18_c52_10;
  wire [7:0] t_r18_c52_11;
  wire [7:0] t_r18_c52_12;
  wire [7:0] t_r18_c53_0;
  wire [7:0] t_r18_c53_1;
  wire [7:0] t_r18_c53_2;
  wire [7:0] t_r18_c53_3;
  wire [7:0] t_r18_c53_4;
  wire [7:0] t_r18_c53_5;
  wire [7:0] t_r18_c53_6;
  wire [7:0] t_r18_c53_7;
  wire [7:0] t_r18_c53_8;
  wire [7:0] t_r18_c53_9;
  wire [7:0] t_r18_c53_10;
  wire [7:0] t_r18_c53_11;
  wire [7:0] t_r18_c53_12;
  wire [7:0] t_r18_c54_0;
  wire [7:0] t_r18_c54_1;
  wire [7:0] t_r18_c54_2;
  wire [7:0] t_r18_c54_3;
  wire [7:0] t_r18_c54_4;
  wire [7:0] t_r18_c54_5;
  wire [7:0] t_r18_c54_6;
  wire [7:0] t_r18_c54_7;
  wire [7:0] t_r18_c54_8;
  wire [7:0] t_r18_c54_9;
  wire [7:0] t_r18_c54_10;
  wire [7:0] t_r18_c54_11;
  wire [7:0] t_r18_c54_12;
  wire [7:0] t_r18_c55_0;
  wire [7:0] t_r18_c55_1;
  wire [7:0] t_r18_c55_2;
  wire [7:0] t_r18_c55_3;
  wire [7:0] t_r18_c55_4;
  wire [7:0] t_r18_c55_5;
  wire [7:0] t_r18_c55_6;
  wire [7:0] t_r18_c55_7;
  wire [7:0] t_r18_c55_8;
  wire [7:0] t_r18_c55_9;
  wire [7:0] t_r18_c55_10;
  wire [7:0] t_r18_c55_11;
  wire [7:0] t_r18_c55_12;
  wire [7:0] t_r18_c56_0;
  wire [7:0] t_r18_c56_1;
  wire [7:0] t_r18_c56_2;
  wire [7:0] t_r18_c56_3;
  wire [7:0] t_r18_c56_4;
  wire [7:0] t_r18_c56_5;
  wire [7:0] t_r18_c56_6;
  wire [7:0] t_r18_c56_7;
  wire [7:0] t_r18_c56_8;
  wire [7:0] t_r18_c56_9;
  wire [7:0] t_r18_c56_10;
  wire [7:0] t_r18_c56_11;
  wire [7:0] t_r18_c56_12;
  wire [7:0] t_r18_c57_0;
  wire [7:0] t_r18_c57_1;
  wire [7:0] t_r18_c57_2;
  wire [7:0] t_r18_c57_3;
  wire [7:0] t_r18_c57_4;
  wire [7:0] t_r18_c57_5;
  wire [7:0] t_r18_c57_6;
  wire [7:0] t_r18_c57_7;
  wire [7:0] t_r18_c57_8;
  wire [7:0] t_r18_c57_9;
  wire [7:0] t_r18_c57_10;
  wire [7:0] t_r18_c57_11;
  wire [7:0] t_r18_c57_12;
  wire [7:0] t_r18_c58_0;
  wire [7:0] t_r18_c58_1;
  wire [7:0] t_r18_c58_2;
  wire [7:0] t_r18_c58_3;
  wire [7:0] t_r18_c58_4;
  wire [7:0] t_r18_c58_5;
  wire [7:0] t_r18_c58_6;
  wire [7:0] t_r18_c58_7;
  wire [7:0] t_r18_c58_8;
  wire [7:0] t_r18_c58_9;
  wire [7:0] t_r18_c58_10;
  wire [7:0] t_r18_c58_11;
  wire [7:0] t_r18_c58_12;
  wire [7:0] t_r18_c59_0;
  wire [7:0] t_r18_c59_1;
  wire [7:0] t_r18_c59_2;
  wire [7:0] t_r18_c59_3;
  wire [7:0] t_r18_c59_4;
  wire [7:0] t_r18_c59_5;
  wire [7:0] t_r18_c59_6;
  wire [7:0] t_r18_c59_7;
  wire [7:0] t_r18_c59_8;
  wire [7:0] t_r18_c59_9;
  wire [7:0] t_r18_c59_10;
  wire [7:0] t_r18_c59_11;
  wire [7:0] t_r18_c59_12;
  wire [7:0] t_r18_c60_0;
  wire [7:0] t_r18_c60_1;
  wire [7:0] t_r18_c60_2;
  wire [7:0] t_r18_c60_3;
  wire [7:0] t_r18_c60_4;
  wire [7:0] t_r18_c60_5;
  wire [7:0] t_r18_c60_6;
  wire [7:0] t_r18_c60_7;
  wire [7:0] t_r18_c60_8;
  wire [7:0] t_r18_c60_9;
  wire [7:0] t_r18_c60_10;
  wire [7:0] t_r18_c60_11;
  wire [7:0] t_r18_c60_12;
  wire [7:0] t_r18_c61_0;
  wire [7:0] t_r18_c61_1;
  wire [7:0] t_r18_c61_2;
  wire [7:0] t_r18_c61_3;
  wire [7:0] t_r18_c61_4;
  wire [7:0] t_r18_c61_5;
  wire [7:0] t_r18_c61_6;
  wire [7:0] t_r18_c61_7;
  wire [7:0] t_r18_c61_8;
  wire [7:0] t_r18_c61_9;
  wire [7:0] t_r18_c61_10;
  wire [7:0] t_r18_c61_11;
  wire [7:0] t_r18_c61_12;
  wire [7:0] t_r18_c62_0;
  wire [7:0] t_r18_c62_1;
  wire [7:0] t_r18_c62_2;
  wire [7:0] t_r18_c62_3;
  wire [7:0] t_r18_c62_4;
  wire [7:0] t_r18_c62_5;
  wire [7:0] t_r18_c62_6;
  wire [7:0] t_r18_c62_7;
  wire [7:0] t_r18_c62_8;
  wire [7:0] t_r18_c62_9;
  wire [7:0] t_r18_c62_10;
  wire [7:0] t_r18_c62_11;
  wire [7:0] t_r18_c62_12;
  wire [7:0] t_r18_c63_0;
  wire [7:0] t_r18_c63_1;
  wire [7:0] t_r18_c63_2;
  wire [7:0] t_r18_c63_3;
  wire [7:0] t_r18_c63_4;
  wire [7:0] t_r18_c63_5;
  wire [7:0] t_r18_c63_6;
  wire [7:0] t_r18_c63_7;
  wire [7:0] t_r18_c63_8;
  wire [7:0] t_r18_c63_9;
  wire [7:0] t_r18_c63_10;
  wire [7:0] t_r18_c63_11;
  wire [7:0] t_r18_c63_12;
  wire [7:0] t_r18_c64_0;
  wire [7:0] t_r18_c64_1;
  wire [7:0] t_r18_c64_2;
  wire [7:0] t_r18_c64_3;
  wire [7:0] t_r18_c64_4;
  wire [7:0] t_r18_c64_5;
  wire [7:0] t_r18_c64_6;
  wire [7:0] t_r18_c64_7;
  wire [7:0] t_r18_c64_8;
  wire [7:0] t_r18_c64_9;
  wire [7:0] t_r18_c64_10;
  wire [7:0] t_r18_c64_11;
  wire [7:0] t_r18_c64_12;
  wire [7:0] t_r18_c65_0;
  wire [7:0] t_r18_c65_1;
  wire [7:0] t_r18_c65_2;
  wire [7:0] t_r18_c65_3;
  wire [7:0] t_r18_c65_4;
  wire [7:0] t_r18_c65_5;
  wire [7:0] t_r18_c65_6;
  wire [7:0] t_r18_c65_7;
  wire [7:0] t_r18_c65_8;
  wire [7:0] t_r18_c65_9;
  wire [7:0] t_r18_c65_10;
  wire [7:0] t_r18_c65_11;
  wire [7:0] t_r18_c65_12;
  wire [7:0] t_r19_c0_0;
  wire [7:0] t_r19_c0_1;
  wire [7:0] t_r19_c0_2;
  wire [7:0] t_r19_c0_3;
  wire [7:0] t_r19_c0_4;
  wire [7:0] t_r19_c0_5;
  wire [7:0] t_r19_c0_6;
  wire [7:0] t_r19_c0_7;
  wire [7:0] t_r19_c0_8;
  wire [7:0] t_r19_c0_9;
  wire [7:0] t_r19_c0_10;
  wire [7:0] t_r19_c0_11;
  wire [7:0] t_r19_c0_12;
  wire [7:0] t_r19_c1_0;
  wire [7:0] t_r19_c1_1;
  wire [7:0] t_r19_c1_2;
  wire [7:0] t_r19_c1_3;
  wire [7:0] t_r19_c1_4;
  wire [7:0] t_r19_c1_5;
  wire [7:0] t_r19_c1_6;
  wire [7:0] t_r19_c1_7;
  wire [7:0] t_r19_c1_8;
  wire [7:0] t_r19_c1_9;
  wire [7:0] t_r19_c1_10;
  wire [7:0] t_r19_c1_11;
  wire [7:0] t_r19_c1_12;
  wire [7:0] t_r19_c2_0;
  wire [7:0] t_r19_c2_1;
  wire [7:0] t_r19_c2_2;
  wire [7:0] t_r19_c2_3;
  wire [7:0] t_r19_c2_4;
  wire [7:0] t_r19_c2_5;
  wire [7:0] t_r19_c2_6;
  wire [7:0] t_r19_c2_7;
  wire [7:0] t_r19_c2_8;
  wire [7:0] t_r19_c2_9;
  wire [7:0] t_r19_c2_10;
  wire [7:0] t_r19_c2_11;
  wire [7:0] t_r19_c2_12;
  wire [7:0] t_r19_c3_0;
  wire [7:0] t_r19_c3_1;
  wire [7:0] t_r19_c3_2;
  wire [7:0] t_r19_c3_3;
  wire [7:0] t_r19_c3_4;
  wire [7:0] t_r19_c3_5;
  wire [7:0] t_r19_c3_6;
  wire [7:0] t_r19_c3_7;
  wire [7:0] t_r19_c3_8;
  wire [7:0] t_r19_c3_9;
  wire [7:0] t_r19_c3_10;
  wire [7:0] t_r19_c3_11;
  wire [7:0] t_r19_c3_12;
  wire [7:0] t_r19_c4_0;
  wire [7:0] t_r19_c4_1;
  wire [7:0] t_r19_c4_2;
  wire [7:0] t_r19_c4_3;
  wire [7:0] t_r19_c4_4;
  wire [7:0] t_r19_c4_5;
  wire [7:0] t_r19_c4_6;
  wire [7:0] t_r19_c4_7;
  wire [7:0] t_r19_c4_8;
  wire [7:0] t_r19_c4_9;
  wire [7:0] t_r19_c4_10;
  wire [7:0] t_r19_c4_11;
  wire [7:0] t_r19_c4_12;
  wire [7:0] t_r19_c5_0;
  wire [7:0] t_r19_c5_1;
  wire [7:0] t_r19_c5_2;
  wire [7:0] t_r19_c5_3;
  wire [7:0] t_r19_c5_4;
  wire [7:0] t_r19_c5_5;
  wire [7:0] t_r19_c5_6;
  wire [7:0] t_r19_c5_7;
  wire [7:0] t_r19_c5_8;
  wire [7:0] t_r19_c5_9;
  wire [7:0] t_r19_c5_10;
  wire [7:0] t_r19_c5_11;
  wire [7:0] t_r19_c5_12;
  wire [7:0] t_r19_c6_0;
  wire [7:0] t_r19_c6_1;
  wire [7:0] t_r19_c6_2;
  wire [7:0] t_r19_c6_3;
  wire [7:0] t_r19_c6_4;
  wire [7:0] t_r19_c6_5;
  wire [7:0] t_r19_c6_6;
  wire [7:0] t_r19_c6_7;
  wire [7:0] t_r19_c6_8;
  wire [7:0] t_r19_c6_9;
  wire [7:0] t_r19_c6_10;
  wire [7:0] t_r19_c6_11;
  wire [7:0] t_r19_c6_12;
  wire [7:0] t_r19_c7_0;
  wire [7:0] t_r19_c7_1;
  wire [7:0] t_r19_c7_2;
  wire [7:0] t_r19_c7_3;
  wire [7:0] t_r19_c7_4;
  wire [7:0] t_r19_c7_5;
  wire [7:0] t_r19_c7_6;
  wire [7:0] t_r19_c7_7;
  wire [7:0] t_r19_c7_8;
  wire [7:0] t_r19_c7_9;
  wire [7:0] t_r19_c7_10;
  wire [7:0] t_r19_c7_11;
  wire [7:0] t_r19_c7_12;
  wire [7:0] t_r19_c8_0;
  wire [7:0] t_r19_c8_1;
  wire [7:0] t_r19_c8_2;
  wire [7:0] t_r19_c8_3;
  wire [7:0] t_r19_c8_4;
  wire [7:0] t_r19_c8_5;
  wire [7:0] t_r19_c8_6;
  wire [7:0] t_r19_c8_7;
  wire [7:0] t_r19_c8_8;
  wire [7:0] t_r19_c8_9;
  wire [7:0] t_r19_c8_10;
  wire [7:0] t_r19_c8_11;
  wire [7:0] t_r19_c8_12;
  wire [7:0] t_r19_c9_0;
  wire [7:0] t_r19_c9_1;
  wire [7:0] t_r19_c9_2;
  wire [7:0] t_r19_c9_3;
  wire [7:0] t_r19_c9_4;
  wire [7:0] t_r19_c9_5;
  wire [7:0] t_r19_c9_6;
  wire [7:0] t_r19_c9_7;
  wire [7:0] t_r19_c9_8;
  wire [7:0] t_r19_c9_9;
  wire [7:0] t_r19_c9_10;
  wire [7:0] t_r19_c9_11;
  wire [7:0] t_r19_c9_12;
  wire [7:0] t_r19_c10_0;
  wire [7:0] t_r19_c10_1;
  wire [7:0] t_r19_c10_2;
  wire [7:0] t_r19_c10_3;
  wire [7:0] t_r19_c10_4;
  wire [7:0] t_r19_c10_5;
  wire [7:0] t_r19_c10_6;
  wire [7:0] t_r19_c10_7;
  wire [7:0] t_r19_c10_8;
  wire [7:0] t_r19_c10_9;
  wire [7:0] t_r19_c10_10;
  wire [7:0] t_r19_c10_11;
  wire [7:0] t_r19_c10_12;
  wire [7:0] t_r19_c11_0;
  wire [7:0] t_r19_c11_1;
  wire [7:0] t_r19_c11_2;
  wire [7:0] t_r19_c11_3;
  wire [7:0] t_r19_c11_4;
  wire [7:0] t_r19_c11_5;
  wire [7:0] t_r19_c11_6;
  wire [7:0] t_r19_c11_7;
  wire [7:0] t_r19_c11_8;
  wire [7:0] t_r19_c11_9;
  wire [7:0] t_r19_c11_10;
  wire [7:0] t_r19_c11_11;
  wire [7:0] t_r19_c11_12;
  wire [7:0] t_r19_c12_0;
  wire [7:0] t_r19_c12_1;
  wire [7:0] t_r19_c12_2;
  wire [7:0] t_r19_c12_3;
  wire [7:0] t_r19_c12_4;
  wire [7:0] t_r19_c12_5;
  wire [7:0] t_r19_c12_6;
  wire [7:0] t_r19_c12_7;
  wire [7:0] t_r19_c12_8;
  wire [7:0] t_r19_c12_9;
  wire [7:0] t_r19_c12_10;
  wire [7:0] t_r19_c12_11;
  wire [7:0] t_r19_c12_12;
  wire [7:0] t_r19_c13_0;
  wire [7:0] t_r19_c13_1;
  wire [7:0] t_r19_c13_2;
  wire [7:0] t_r19_c13_3;
  wire [7:0] t_r19_c13_4;
  wire [7:0] t_r19_c13_5;
  wire [7:0] t_r19_c13_6;
  wire [7:0] t_r19_c13_7;
  wire [7:0] t_r19_c13_8;
  wire [7:0] t_r19_c13_9;
  wire [7:0] t_r19_c13_10;
  wire [7:0] t_r19_c13_11;
  wire [7:0] t_r19_c13_12;
  wire [7:0] t_r19_c14_0;
  wire [7:0] t_r19_c14_1;
  wire [7:0] t_r19_c14_2;
  wire [7:0] t_r19_c14_3;
  wire [7:0] t_r19_c14_4;
  wire [7:0] t_r19_c14_5;
  wire [7:0] t_r19_c14_6;
  wire [7:0] t_r19_c14_7;
  wire [7:0] t_r19_c14_8;
  wire [7:0] t_r19_c14_9;
  wire [7:0] t_r19_c14_10;
  wire [7:0] t_r19_c14_11;
  wire [7:0] t_r19_c14_12;
  wire [7:0] t_r19_c15_0;
  wire [7:0] t_r19_c15_1;
  wire [7:0] t_r19_c15_2;
  wire [7:0] t_r19_c15_3;
  wire [7:0] t_r19_c15_4;
  wire [7:0] t_r19_c15_5;
  wire [7:0] t_r19_c15_6;
  wire [7:0] t_r19_c15_7;
  wire [7:0] t_r19_c15_8;
  wire [7:0] t_r19_c15_9;
  wire [7:0] t_r19_c15_10;
  wire [7:0] t_r19_c15_11;
  wire [7:0] t_r19_c15_12;
  wire [7:0] t_r19_c16_0;
  wire [7:0] t_r19_c16_1;
  wire [7:0] t_r19_c16_2;
  wire [7:0] t_r19_c16_3;
  wire [7:0] t_r19_c16_4;
  wire [7:0] t_r19_c16_5;
  wire [7:0] t_r19_c16_6;
  wire [7:0] t_r19_c16_7;
  wire [7:0] t_r19_c16_8;
  wire [7:0] t_r19_c16_9;
  wire [7:0] t_r19_c16_10;
  wire [7:0] t_r19_c16_11;
  wire [7:0] t_r19_c16_12;
  wire [7:0] t_r19_c17_0;
  wire [7:0] t_r19_c17_1;
  wire [7:0] t_r19_c17_2;
  wire [7:0] t_r19_c17_3;
  wire [7:0] t_r19_c17_4;
  wire [7:0] t_r19_c17_5;
  wire [7:0] t_r19_c17_6;
  wire [7:0] t_r19_c17_7;
  wire [7:0] t_r19_c17_8;
  wire [7:0] t_r19_c17_9;
  wire [7:0] t_r19_c17_10;
  wire [7:0] t_r19_c17_11;
  wire [7:0] t_r19_c17_12;
  wire [7:0] t_r19_c18_0;
  wire [7:0] t_r19_c18_1;
  wire [7:0] t_r19_c18_2;
  wire [7:0] t_r19_c18_3;
  wire [7:0] t_r19_c18_4;
  wire [7:0] t_r19_c18_5;
  wire [7:0] t_r19_c18_6;
  wire [7:0] t_r19_c18_7;
  wire [7:0] t_r19_c18_8;
  wire [7:0] t_r19_c18_9;
  wire [7:0] t_r19_c18_10;
  wire [7:0] t_r19_c18_11;
  wire [7:0] t_r19_c18_12;
  wire [7:0] t_r19_c19_0;
  wire [7:0] t_r19_c19_1;
  wire [7:0] t_r19_c19_2;
  wire [7:0] t_r19_c19_3;
  wire [7:0] t_r19_c19_4;
  wire [7:0] t_r19_c19_5;
  wire [7:0] t_r19_c19_6;
  wire [7:0] t_r19_c19_7;
  wire [7:0] t_r19_c19_8;
  wire [7:0] t_r19_c19_9;
  wire [7:0] t_r19_c19_10;
  wire [7:0] t_r19_c19_11;
  wire [7:0] t_r19_c19_12;
  wire [7:0] t_r19_c20_0;
  wire [7:0] t_r19_c20_1;
  wire [7:0] t_r19_c20_2;
  wire [7:0] t_r19_c20_3;
  wire [7:0] t_r19_c20_4;
  wire [7:0] t_r19_c20_5;
  wire [7:0] t_r19_c20_6;
  wire [7:0] t_r19_c20_7;
  wire [7:0] t_r19_c20_8;
  wire [7:0] t_r19_c20_9;
  wire [7:0] t_r19_c20_10;
  wire [7:0] t_r19_c20_11;
  wire [7:0] t_r19_c20_12;
  wire [7:0] t_r19_c21_0;
  wire [7:0] t_r19_c21_1;
  wire [7:0] t_r19_c21_2;
  wire [7:0] t_r19_c21_3;
  wire [7:0] t_r19_c21_4;
  wire [7:0] t_r19_c21_5;
  wire [7:0] t_r19_c21_6;
  wire [7:0] t_r19_c21_7;
  wire [7:0] t_r19_c21_8;
  wire [7:0] t_r19_c21_9;
  wire [7:0] t_r19_c21_10;
  wire [7:0] t_r19_c21_11;
  wire [7:0] t_r19_c21_12;
  wire [7:0] t_r19_c22_0;
  wire [7:0] t_r19_c22_1;
  wire [7:0] t_r19_c22_2;
  wire [7:0] t_r19_c22_3;
  wire [7:0] t_r19_c22_4;
  wire [7:0] t_r19_c22_5;
  wire [7:0] t_r19_c22_6;
  wire [7:0] t_r19_c22_7;
  wire [7:0] t_r19_c22_8;
  wire [7:0] t_r19_c22_9;
  wire [7:0] t_r19_c22_10;
  wire [7:0] t_r19_c22_11;
  wire [7:0] t_r19_c22_12;
  wire [7:0] t_r19_c23_0;
  wire [7:0] t_r19_c23_1;
  wire [7:0] t_r19_c23_2;
  wire [7:0] t_r19_c23_3;
  wire [7:0] t_r19_c23_4;
  wire [7:0] t_r19_c23_5;
  wire [7:0] t_r19_c23_6;
  wire [7:0] t_r19_c23_7;
  wire [7:0] t_r19_c23_8;
  wire [7:0] t_r19_c23_9;
  wire [7:0] t_r19_c23_10;
  wire [7:0] t_r19_c23_11;
  wire [7:0] t_r19_c23_12;
  wire [7:0] t_r19_c24_0;
  wire [7:0] t_r19_c24_1;
  wire [7:0] t_r19_c24_2;
  wire [7:0] t_r19_c24_3;
  wire [7:0] t_r19_c24_4;
  wire [7:0] t_r19_c24_5;
  wire [7:0] t_r19_c24_6;
  wire [7:0] t_r19_c24_7;
  wire [7:0] t_r19_c24_8;
  wire [7:0] t_r19_c24_9;
  wire [7:0] t_r19_c24_10;
  wire [7:0] t_r19_c24_11;
  wire [7:0] t_r19_c24_12;
  wire [7:0] t_r19_c25_0;
  wire [7:0] t_r19_c25_1;
  wire [7:0] t_r19_c25_2;
  wire [7:0] t_r19_c25_3;
  wire [7:0] t_r19_c25_4;
  wire [7:0] t_r19_c25_5;
  wire [7:0] t_r19_c25_6;
  wire [7:0] t_r19_c25_7;
  wire [7:0] t_r19_c25_8;
  wire [7:0] t_r19_c25_9;
  wire [7:0] t_r19_c25_10;
  wire [7:0] t_r19_c25_11;
  wire [7:0] t_r19_c25_12;
  wire [7:0] t_r19_c26_0;
  wire [7:0] t_r19_c26_1;
  wire [7:0] t_r19_c26_2;
  wire [7:0] t_r19_c26_3;
  wire [7:0] t_r19_c26_4;
  wire [7:0] t_r19_c26_5;
  wire [7:0] t_r19_c26_6;
  wire [7:0] t_r19_c26_7;
  wire [7:0] t_r19_c26_8;
  wire [7:0] t_r19_c26_9;
  wire [7:0] t_r19_c26_10;
  wire [7:0] t_r19_c26_11;
  wire [7:0] t_r19_c26_12;
  wire [7:0] t_r19_c27_0;
  wire [7:0] t_r19_c27_1;
  wire [7:0] t_r19_c27_2;
  wire [7:0] t_r19_c27_3;
  wire [7:0] t_r19_c27_4;
  wire [7:0] t_r19_c27_5;
  wire [7:0] t_r19_c27_6;
  wire [7:0] t_r19_c27_7;
  wire [7:0] t_r19_c27_8;
  wire [7:0] t_r19_c27_9;
  wire [7:0] t_r19_c27_10;
  wire [7:0] t_r19_c27_11;
  wire [7:0] t_r19_c27_12;
  wire [7:0] t_r19_c28_0;
  wire [7:0] t_r19_c28_1;
  wire [7:0] t_r19_c28_2;
  wire [7:0] t_r19_c28_3;
  wire [7:0] t_r19_c28_4;
  wire [7:0] t_r19_c28_5;
  wire [7:0] t_r19_c28_6;
  wire [7:0] t_r19_c28_7;
  wire [7:0] t_r19_c28_8;
  wire [7:0] t_r19_c28_9;
  wire [7:0] t_r19_c28_10;
  wire [7:0] t_r19_c28_11;
  wire [7:0] t_r19_c28_12;
  wire [7:0] t_r19_c29_0;
  wire [7:0] t_r19_c29_1;
  wire [7:0] t_r19_c29_2;
  wire [7:0] t_r19_c29_3;
  wire [7:0] t_r19_c29_4;
  wire [7:0] t_r19_c29_5;
  wire [7:0] t_r19_c29_6;
  wire [7:0] t_r19_c29_7;
  wire [7:0] t_r19_c29_8;
  wire [7:0] t_r19_c29_9;
  wire [7:0] t_r19_c29_10;
  wire [7:0] t_r19_c29_11;
  wire [7:0] t_r19_c29_12;
  wire [7:0] t_r19_c30_0;
  wire [7:0] t_r19_c30_1;
  wire [7:0] t_r19_c30_2;
  wire [7:0] t_r19_c30_3;
  wire [7:0] t_r19_c30_4;
  wire [7:0] t_r19_c30_5;
  wire [7:0] t_r19_c30_6;
  wire [7:0] t_r19_c30_7;
  wire [7:0] t_r19_c30_8;
  wire [7:0] t_r19_c30_9;
  wire [7:0] t_r19_c30_10;
  wire [7:0] t_r19_c30_11;
  wire [7:0] t_r19_c30_12;
  wire [7:0] t_r19_c31_0;
  wire [7:0] t_r19_c31_1;
  wire [7:0] t_r19_c31_2;
  wire [7:0] t_r19_c31_3;
  wire [7:0] t_r19_c31_4;
  wire [7:0] t_r19_c31_5;
  wire [7:0] t_r19_c31_6;
  wire [7:0] t_r19_c31_7;
  wire [7:0] t_r19_c31_8;
  wire [7:0] t_r19_c31_9;
  wire [7:0] t_r19_c31_10;
  wire [7:0] t_r19_c31_11;
  wire [7:0] t_r19_c31_12;
  wire [7:0] t_r19_c32_0;
  wire [7:0] t_r19_c32_1;
  wire [7:0] t_r19_c32_2;
  wire [7:0] t_r19_c32_3;
  wire [7:0] t_r19_c32_4;
  wire [7:0] t_r19_c32_5;
  wire [7:0] t_r19_c32_6;
  wire [7:0] t_r19_c32_7;
  wire [7:0] t_r19_c32_8;
  wire [7:0] t_r19_c32_9;
  wire [7:0] t_r19_c32_10;
  wire [7:0] t_r19_c32_11;
  wire [7:0] t_r19_c32_12;
  wire [7:0] t_r19_c33_0;
  wire [7:0] t_r19_c33_1;
  wire [7:0] t_r19_c33_2;
  wire [7:0] t_r19_c33_3;
  wire [7:0] t_r19_c33_4;
  wire [7:0] t_r19_c33_5;
  wire [7:0] t_r19_c33_6;
  wire [7:0] t_r19_c33_7;
  wire [7:0] t_r19_c33_8;
  wire [7:0] t_r19_c33_9;
  wire [7:0] t_r19_c33_10;
  wire [7:0] t_r19_c33_11;
  wire [7:0] t_r19_c33_12;
  wire [7:0] t_r19_c34_0;
  wire [7:0] t_r19_c34_1;
  wire [7:0] t_r19_c34_2;
  wire [7:0] t_r19_c34_3;
  wire [7:0] t_r19_c34_4;
  wire [7:0] t_r19_c34_5;
  wire [7:0] t_r19_c34_6;
  wire [7:0] t_r19_c34_7;
  wire [7:0] t_r19_c34_8;
  wire [7:0] t_r19_c34_9;
  wire [7:0] t_r19_c34_10;
  wire [7:0] t_r19_c34_11;
  wire [7:0] t_r19_c34_12;
  wire [7:0] t_r19_c35_0;
  wire [7:0] t_r19_c35_1;
  wire [7:0] t_r19_c35_2;
  wire [7:0] t_r19_c35_3;
  wire [7:0] t_r19_c35_4;
  wire [7:0] t_r19_c35_5;
  wire [7:0] t_r19_c35_6;
  wire [7:0] t_r19_c35_7;
  wire [7:0] t_r19_c35_8;
  wire [7:0] t_r19_c35_9;
  wire [7:0] t_r19_c35_10;
  wire [7:0] t_r19_c35_11;
  wire [7:0] t_r19_c35_12;
  wire [7:0] t_r19_c36_0;
  wire [7:0] t_r19_c36_1;
  wire [7:0] t_r19_c36_2;
  wire [7:0] t_r19_c36_3;
  wire [7:0] t_r19_c36_4;
  wire [7:0] t_r19_c36_5;
  wire [7:0] t_r19_c36_6;
  wire [7:0] t_r19_c36_7;
  wire [7:0] t_r19_c36_8;
  wire [7:0] t_r19_c36_9;
  wire [7:0] t_r19_c36_10;
  wire [7:0] t_r19_c36_11;
  wire [7:0] t_r19_c36_12;
  wire [7:0] t_r19_c37_0;
  wire [7:0] t_r19_c37_1;
  wire [7:0] t_r19_c37_2;
  wire [7:0] t_r19_c37_3;
  wire [7:0] t_r19_c37_4;
  wire [7:0] t_r19_c37_5;
  wire [7:0] t_r19_c37_6;
  wire [7:0] t_r19_c37_7;
  wire [7:0] t_r19_c37_8;
  wire [7:0] t_r19_c37_9;
  wire [7:0] t_r19_c37_10;
  wire [7:0] t_r19_c37_11;
  wire [7:0] t_r19_c37_12;
  wire [7:0] t_r19_c38_0;
  wire [7:0] t_r19_c38_1;
  wire [7:0] t_r19_c38_2;
  wire [7:0] t_r19_c38_3;
  wire [7:0] t_r19_c38_4;
  wire [7:0] t_r19_c38_5;
  wire [7:0] t_r19_c38_6;
  wire [7:0] t_r19_c38_7;
  wire [7:0] t_r19_c38_8;
  wire [7:0] t_r19_c38_9;
  wire [7:0] t_r19_c38_10;
  wire [7:0] t_r19_c38_11;
  wire [7:0] t_r19_c38_12;
  wire [7:0] t_r19_c39_0;
  wire [7:0] t_r19_c39_1;
  wire [7:0] t_r19_c39_2;
  wire [7:0] t_r19_c39_3;
  wire [7:0] t_r19_c39_4;
  wire [7:0] t_r19_c39_5;
  wire [7:0] t_r19_c39_6;
  wire [7:0] t_r19_c39_7;
  wire [7:0] t_r19_c39_8;
  wire [7:0] t_r19_c39_9;
  wire [7:0] t_r19_c39_10;
  wire [7:0] t_r19_c39_11;
  wire [7:0] t_r19_c39_12;
  wire [7:0] t_r19_c40_0;
  wire [7:0] t_r19_c40_1;
  wire [7:0] t_r19_c40_2;
  wire [7:0] t_r19_c40_3;
  wire [7:0] t_r19_c40_4;
  wire [7:0] t_r19_c40_5;
  wire [7:0] t_r19_c40_6;
  wire [7:0] t_r19_c40_7;
  wire [7:0] t_r19_c40_8;
  wire [7:0] t_r19_c40_9;
  wire [7:0] t_r19_c40_10;
  wire [7:0] t_r19_c40_11;
  wire [7:0] t_r19_c40_12;
  wire [7:0] t_r19_c41_0;
  wire [7:0] t_r19_c41_1;
  wire [7:0] t_r19_c41_2;
  wire [7:0] t_r19_c41_3;
  wire [7:0] t_r19_c41_4;
  wire [7:0] t_r19_c41_5;
  wire [7:0] t_r19_c41_6;
  wire [7:0] t_r19_c41_7;
  wire [7:0] t_r19_c41_8;
  wire [7:0] t_r19_c41_9;
  wire [7:0] t_r19_c41_10;
  wire [7:0] t_r19_c41_11;
  wire [7:0] t_r19_c41_12;
  wire [7:0] t_r19_c42_0;
  wire [7:0] t_r19_c42_1;
  wire [7:0] t_r19_c42_2;
  wire [7:0] t_r19_c42_3;
  wire [7:0] t_r19_c42_4;
  wire [7:0] t_r19_c42_5;
  wire [7:0] t_r19_c42_6;
  wire [7:0] t_r19_c42_7;
  wire [7:0] t_r19_c42_8;
  wire [7:0] t_r19_c42_9;
  wire [7:0] t_r19_c42_10;
  wire [7:0] t_r19_c42_11;
  wire [7:0] t_r19_c42_12;
  wire [7:0] t_r19_c43_0;
  wire [7:0] t_r19_c43_1;
  wire [7:0] t_r19_c43_2;
  wire [7:0] t_r19_c43_3;
  wire [7:0] t_r19_c43_4;
  wire [7:0] t_r19_c43_5;
  wire [7:0] t_r19_c43_6;
  wire [7:0] t_r19_c43_7;
  wire [7:0] t_r19_c43_8;
  wire [7:0] t_r19_c43_9;
  wire [7:0] t_r19_c43_10;
  wire [7:0] t_r19_c43_11;
  wire [7:0] t_r19_c43_12;
  wire [7:0] t_r19_c44_0;
  wire [7:0] t_r19_c44_1;
  wire [7:0] t_r19_c44_2;
  wire [7:0] t_r19_c44_3;
  wire [7:0] t_r19_c44_4;
  wire [7:0] t_r19_c44_5;
  wire [7:0] t_r19_c44_6;
  wire [7:0] t_r19_c44_7;
  wire [7:0] t_r19_c44_8;
  wire [7:0] t_r19_c44_9;
  wire [7:0] t_r19_c44_10;
  wire [7:0] t_r19_c44_11;
  wire [7:0] t_r19_c44_12;
  wire [7:0] t_r19_c45_0;
  wire [7:0] t_r19_c45_1;
  wire [7:0] t_r19_c45_2;
  wire [7:0] t_r19_c45_3;
  wire [7:0] t_r19_c45_4;
  wire [7:0] t_r19_c45_5;
  wire [7:0] t_r19_c45_6;
  wire [7:0] t_r19_c45_7;
  wire [7:0] t_r19_c45_8;
  wire [7:0] t_r19_c45_9;
  wire [7:0] t_r19_c45_10;
  wire [7:0] t_r19_c45_11;
  wire [7:0] t_r19_c45_12;
  wire [7:0] t_r19_c46_0;
  wire [7:0] t_r19_c46_1;
  wire [7:0] t_r19_c46_2;
  wire [7:0] t_r19_c46_3;
  wire [7:0] t_r19_c46_4;
  wire [7:0] t_r19_c46_5;
  wire [7:0] t_r19_c46_6;
  wire [7:0] t_r19_c46_7;
  wire [7:0] t_r19_c46_8;
  wire [7:0] t_r19_c46_9;
  wire [7:0] t_r19_c46_10;
  wire [7:0] t_r19_c46_11;
  wire [7:0] t_r19_c46_12;
  wire [7:0] t_r19_c47_0;
  wire [7:0] t_r19_c47_1;
  wire [7:0] t_r19_c47_2;
  wire [7:0] t_r19_c47_3;
  wire [7:0] t_r19_c47_4;
  wire [7:0] t_r19_c47_5;
  wire [7:0] t_r19_c47_6;
  wire [7:0] t_r19_c47_7;
  wire [7:0] t_r19_c47_8;
  wire [7:0] t_r19_c47_9;
  wire [7:0] t_r19_c47_10;
  wire [7:0] t_r19_c47_11;
  wire [7:0] t_r19_c47_12;
  wire [7:0] t_r19_c48_0;
  wire [7:0] t_r19_c48_1;
  wire [7:0] t_r19_c48_2;
  wire [7:0] t_r19_c48_3;
  wire [7:0] t_r19_c48_4;
  wire [7:0] t_r19_c48_5;
  wire [7:0] t_r19_c48_6;
  wire [7:0] t_r19_c48_7;
  wire [7:0] t_r19_c48_8;
  wire [7:0] t_r19_c48_9;
  wire [7:0] t_r19_c48_10;
  wire [7:0] t_r19_c48_11;
  wire [7:0] t_r19_c48_12;
  wire [7:0] t_r19_c49_0;
  wire [7:0] t_r19_c49_1;
  wire [7:0] t_r19_c49_2;
  wire [7:0] t_r19_c49_3;
  wire [7:0] t_r19_c49_4;
  wire [7:0] t_r19_c49_5;
  wire [7:0] t_r19_c49_6;
  wire [7:0] t_r19_c49_7;
  wire [7:0] t_r19_c49_8;
  wire [7:0] t_r19_c49_9;
  wire [7:0] t_r19_c49_10;
  wire [7:0] t_r19_c49_11;
  wire [7:0] t_r19_c49_12;
  wire [7:0] t_r19_c50_0;
  wire [7:0] t_r19_c50_1;
  wire [7:0] t_r19_c50_2;
  wire [7:0] t_r19_c50_3;
  wire [7:0] t_r19_c50_4;
  wire [7:0] t_r19_c50_5;
  wire [7:0] t_r19_c50_6;
  wire [7:0] t_r19_c50_7;
  wire [7:0] t_r19_c50_8;
  wire [7:0] t_r19_c50_9;
  wire [7:0] t_r19_c50_10;
  wire [7:0] t_r19_c50_11;
  wire [7:0] t_r19_c50_12;
  wire [7:0] t_r19_c51_0;
  wire [7:0] t_r19_c51_1;
  wire [7:0] t_r19_c51_2;
  wire [7:0] t_r19_c51_3;
  wire [7:0] t_r19_c51_4;
  wire [7:0] t_r19_c51_5;
  wire [7:0] t_r19_c51_6;
  wire [7:0] t_r19_c51_7;
  wire [7:0] t_r19_c51_8;
  wire [7:0] t_r19_c51_9;
  wire [7:0] t_r19_c51_10;
  wire [7:0] t_r19_c51_11;
  wire [7:0] t_r19_c51_12;
  wire [7:0] t_r19_c52_0;
  wire [7:0] t_r19_c52_1;
  wire [7:0] t_r19_c52_2;
  wire [7:0] t_r19_c52_3;
  wire [7:0] t_r19_c52_4;
  wire [7:0] t_r19_c52_5;
  wire [7:0] t_r19_c52_6;
  wire [7:0] t_r19_c52_7;
  wire [7:0] t_r19_c52_8;
  wire [7:0] t_r19_c52_9;
  wire [7:0] t_r19_c52_10;
  wire [7:0] t_r19_c52_11;
  wire [7:0] t_r19_c52_12;
  wire [7:0] t_r19_c53_0;
  wire [7:0] t_r19_c53_1;
  wire [7:0] t_r19_c53_2;
  wire [7:0] t_r19_c53_3;
  wire [7:0] t_r19_c53_4;
  wire [7:0] t_r19_c53_5;
  wire [7:0] t_r19_c53_6;
  wire [7:0] t_r19_c53_7;
  wire [7:0] t_r19_c53_8;
  wire [7:0] t_r19_c53_9;
  wire [7:0] t_r19_c53_10;
  wire [7:0] t_r19_c53_11;
  wire [7:0] t_r19_c53_12;
  wire [7:0] t_r19_c54_0;
  wire [7:0] t_r19_c54_1;
  wire [7:0] t_r19_c54_2;
  wire [7:0] t_r19_c54_3;
  wire [7:0] t_r19_c54_4;
  wire [7:0] t_r19_c54_5;
  wire [7:0] t_r19_c54_6;
  wire [7:0] t_r19_c54_7;
  wire [7:0] t_r19_c54_8;
  wire [7:0] t_r19_c54_9;
  wire [7:0] t_r19_c54_10;
  wire [7:0] t_r19_c54_11;
  wire [7:0] t_r19_c54_12;
  wire [7:0] t_r19_c55_0;
  wire [7:0] t_r19_c55_1;
  wire [7:0] t_r19_c55_2;
  wire [7:0] t_r19_c55_3;
  wire [7:0] t_r19_c55_4;
  wire [7:0] t_r19_c55_5;
  wire [7:0] t_r19_c55_6;
  wire [7:0] t_r19_c55_7;
  wire [7:0] t_r19_c55_8;
  wire [7:0] t_r19_c55_9;
  wire [7:0] t_r19_c55_10;
  wire [7:0] t_r19_c55_11;
  wire [7:0] t_r19_c55_12;
  wire [7:0] t_r19_c56_0;
  wire [7:0] t_r19_c56_1;
  wire [7:0] t_r19_c56_2;
  wire [7:0] t_r19_c56_3;
  wire [7:0] t_r19_c56_4;
  wire [7:0] t_r19_c56_5;
  wire [7:0] t_r19_c56_6;
  wire [7:0] t_r19_c56_7;
  wire [7:0] t_r19_c56_8;
  wire [7:0] t_r19_c56_9;
  wire [7:0] t_r19_c56_10;
  wire [7:0] t_r19_c56_11;
  wire [7:0] t_r19_c56_12;
  wire [7:0] t_r19_c57_0;
  wire [7:0] t_r19_c57_1;
  wire [7:0] t_r19_c57_2;
  wire [7:0] t_r19_c57_3;
  wire [7:0] t_r19_c57_4;
  wire [7:0] t_r19_c57_5;
  wire [7:0] t_r19_c57_6;
  wire [7:0] t_r19_c57_7;
  wire [7:0] t_r19_c57_8;
  wire [7:0] t_r19_c57_9;
  wire [7:0] t_r19_c57_10;
  wire [7:0] t_r19_c57_11;
  wire [7:0] t_r19_c57_12;
  wire [7:0] t_r19_c58_0;
  wire [7:0] t_r19_c58_1;
  wire [7:0] t_r19_c58_2;
  wire [7:0] t_r19_c58_3;
  wire [7:0] t_r19_c58_4;
  wire [7:0] t_r19_c58_5;
  wire [7:0] t_r19_c58_6;
  wire [7:0] t_r19_c58_7;
  wire [7:0] t_r19_c58_8;
  wire [7:0] t_r19_c58_9;
  wire [7:0] t_r19_c58_10;
  wire [7:0] t_r19_c58_11;
  wire [7:0] t_r19_c58_12;
  wire [7:0] t_r19_c59_0;
  wire [7:0] t_r19_c59_1;
  wire [7:0] t_r19_c59_2;
  wire [7:0] t_r19_c59_3;
  wire [7:0] t_r19_c59_4;
  wire [7:0] t_r19_c59_5;
  wire [7:0] t_r19_c59_6;
  wire [7:0] t_r19_c59_7;
  wire [7:0] t_r19_c59_8;
  wire [7:0] t_r19_c59_9;
  wire [7:0] t_r19_c59_10;
  wire [7:0] t_r19_c59_11;
  wire [7:0] t_r19_c59_12;
  wire [7:0] t_r19_c60_0;
  wire [7:0] t_r19_c60_1;
  wire [7:0] t_r19_c60_2;
  wire [7:0] t_r19_c60_3;
  wire [7:0] t_r19_c60_4;
  wire [7:0] t_r19_c60_5;
  wire [7:0] t_r19_c60_6;
  wire [7:0] t_r19_c60_7;
  wire [7:0] t_r19_c60_8;
  wire [7:0] t_r19_c60_9;
  wire [7:0] t_r19_c60_10;
  wire [7:0] t_r19_c60_11;
  wire [7:0] t_r19_c60_12;
  wire [7:0] t_r19_c61_0;
  wire [7:0] t_r19_c61_1;
  wire [7:0] t_r19_c61_2;
  wire [7:0] t_r19_c61_3;
  wire [7:0] t_r19_c61_4;
  wire [7:0] t_r19_c61_5;
  wire [7:0] t_r19_c61_6;
  wire [7:0] t_r19_c61_7;
  wire [7:0] t_r19_c61_8;
  wire [7:0] t_r19_c61_9;
  wire [7:0] t_r19_c61_10;
  wire [7:0] t_r19_c61_11;
  wire [7:0] t_r19_c61_12;
  wire [7:0] t_r19_c62_0;
  wire [7:0] t_r19_c62_1;
  wire [7:0] t_r19_c62_2;
  wire [7:0] t_r19_c62_3;
  wire [7:0] t_r19_c62_4;
  wire [7:0] t_r19_c62_5;
  wire [7:0] t_r19_c62_6;
  wire [7:0] t_r19_c62_7;
  wire [7:0] t_r19_c62_8;
  wire [7:0] t_r19_c62_9;
  wire [7:0] t_r19_c62_10;
  wire [7:0] t_r19_c62_11;
  wire [7:0] t_r19_c62_12;
  wire [7:0] t_r19_c63_0;
  wire [7:0] t_r19_c63_1;
  wire [7:0] t_r19_c63_2;
  wire [7:0] t_r19_c63_3;
  wire [7:0] t_r19_c63_4;
  wire [7:0] t_r19_c63_5;
  wire [7:0] t_r19_c63_6;
  wire [7:0] t_r19_c63_7;
  wire [7:0] t_r19_c63_8;
  wire [7:0] t_r19_c63_9;
  wire [7:0] t_r19_c63_10;
  wire [7:0] t_r19_c63_11;
  wire [7:0] t_r19_c63_12;
  wire [7:0] t_r19_c64_0;
  wire [7:0] t_r19_c64_1;
  wire [7:0] t_r19_c64_2;
  wire [7:0] t_r19_c64_3;
  wire [7:0] t_r19_c64_4;
  wire [7:0] t_r19_c64_5;
  wire [7:0] t_r19_c64_6;
  wire [7:0] t_r19_c64_7;
  wire [7:0] t_r19_c64_8;
  wire [7:0] t_r19_c64_9;
  wire [7:0] t_r19_c64_10;
  wire [7:0] t_r19_c64_11;
  wire [7:0] t_r19_c64_12;
  wire [7:0] t_r19_c65_0;
  wire [7:0] t_r19_c65_1;
  wire [7:0] t_r19_c65_2;
  wire [7:0] t_r19_c65_3;
  wire [7:0] t_r19_c65_4;
  wire [7:0] t_r19_c65_5;
  wire [7:0] t_r19_c65_6;
  wire [7:0] t_r19_c65_7;
  wire [7:0] t_r19_c65_8;
  wire [7:0] t_r19_c65_9;
  wire [7:0] t_r19_c65_10;
  wire [7:0] t_r19_c65_11;
  wire [7:0] t_r19_c65_12;
  wire [7:0] t_r20_c0_0;
  wire [7:0] t_r20_c0_1;
  wire [7:0] t_r20_c0_2;
  wire [7:0] t_r20_c0_3;
  wire [7:0] t_r20_c0_4;
  wire [7:0] t_r20_c0_5;
  wire [7:0] t_r20_c0_6;
  wire [7:0] t_r20_c0_7;
  wire [7:0] t_r20_c0_8;
  wire [7:0] t_r20_c0_9;
  wire [7:0] t_r20_c0_10;
  wire [7:0] t_r20_c0_11;
  wire [7:0] t_r20_c0_12;
  wire [7:0] t_r20_c1_0;
  wire [7:0] t_r20_c1_1;
  wire [7:0] t_r20_c1_2;
  wire [7:0] t_r20_c1_3;
  wire [7:0] t_r20_c1_4;
  wire [7:0] t_r20_c1_5;
  wire [7:0] t_r20_c1_6;
  wire [7:0] t_r20_c1_7;
  wire [7:0] t_r20_c1_8;
  wire [7:0] t_r20_c1_9;
  wire [7:0] t_r20_c1_10;
  wire [7:0] t_r20_c1_11;
  wire [7:0] t_r20_c1_12;
  wire [7:0] t_r20_c2_0;
  wire [7:0] t_r20_c2_1;
  wire [7:0] t_r20_c2_2;
  wire [7:0] t_r20_c2_3;
  wire [7:0] t_r20_c2_4;
  wire [7:0] t_r20_c2_5;
  wire [7:0] t_r20_c2_6;
  wire [7:0] t_r20_c2_7;
  wire [7:0] t_r20_c2_8;
  wire [7:0] t_r20_c2_9;
  wire [7:0] t_r20_c2_10;
  wire [7:0] t_r20_c2_11;
  wire [7:0] t_r20_c2_12;
  wire [7:0] t_r20_c3_0;
  wire [7:0] t_r20_c3_1;
  wire [7:0] t_r20_c3_2;
  wire [7:0] t_r20_c3_3;
  wire [7:0] t_r20_c3_4;
  wire [7:0] t_r20_c3_5;
  wire [7:0] t_r20_c3_6;
  wire [7:0] t_r20_c3_7;
  wire [7:0] t_r20_c3_8;
  wire [7:0] t_r20_c3_9;
  wire [7:0] t_r20_c3_10;
  wire [7:0] t_r20_c3_11;
  wire [7:0] t_r20_c3_12;
  wire [7:0] t_r20_c4_0;
  wire [7:0] t_r20_c4_1;
  wire [7:0] t_r20_c4_2;
  wire [7:0] t_r20_c4_3;
  wire [7:0] t_r20_c4_4;
  wire [7:0] t_r20_c4_5;
  wire [7:0] t_r20_c4_6;
  wire [7:0] t_r20_c4_7;
  wire [7:0] t_r20_c4_8;
  wire [7:0] t_r20_c4_9;
  wire [7:0] t_r20_c4_10;
  wire [7:0] t_r20_c4_11;
  wire [7:0] t_r20_c4_12;
  wire [7:0] t_r20_c5_0;
  wire [7:0] t_r20_c5_1;
  wire [7:0] t_r20_c5_2;
  wire [7:0] t_r20_c5_3;
  wire [7:0] t_r20_c5_4;
  wire [7:0] t_r20_c5_5;
  wire [7:0] t_r20_c5_6;
  wire [7:0] t_r20_c5_7;
  wire [7:0] t_r20_c5_8;
  wire [7:0] t_r20_c5_9;
  wire [7:0] t_r20_c5_10;
  wire [7:0] t_r20_c5_11;
  wire [7:0] t_r20_c5_12;
  wire [7:0] t_r20_c6_0;
  wire [7:0] t_r20_c6_1;
  wire [7:0] t_r20_c6_2;
  wire [7:0] t_r20_c6_3;
  wire [7:0] t_r20_c6_4;
  wire [7:0] t_r20_c6_5;
  wire [7:0] t_r20_c6_6;
  wire [7:0] t_r20_c6_7;
  wire [7:0] t_r20_c6_8;
  wire [7:0] t_r20_c6_9;
  wire [7:0] t_r20_c6_10;
  wire [7:0] t_r20_c6_11;
  wire [7:0] t_r20_c6_12;
  wire [7:0] t_r20_c7_0;
  wire [7:0] t_r20_c7_1;
  wire [7:0] t_r20_c7_2;
  wire [7:0] t_r20_c7_3;
  wire [7:0] t_r20_c7_4;
  wire [7:0] t_r20_c7_5;
  wire [7:0] t_r20_c7_6;
  wire [7:0] t_r20_c7_7;
  wire [7:0] t_r20_c7_8;
  wire [7:0] t_r20_c7_9;
  wire [7:0] t_r20_c7_10;
  wire [7:0] t_r20_c7_11;
  wire [7:0] t_r20_c7_12;
  wire [7:0] t_r20_c8_0;
  wire [7:0] t_r20_c8_1;
  wire [7:0] t_r20_c8_2;
  wire [7:0] t_r20_c8_3;
  wire [7:0] t_r20_c8_4;
  wire [7:0] t_r20_c8_5;
  wire [7:0] t_r20_c8_6;
  wire [7:0] t_r20_c8_7;
  wire [7:0] t_r20_c8_8;
  wire [7:0] t_r20_c8_9;
  wire [7:0] t_r20_c8_10;
  wire [7:0] t_r20_c8_11;
  wire [7:0] t_r20_c8_12;
  wire [7:0] t_r20_c9_0;
  wire [7:0] t_r20_c9_1;
  wire [7:0] t_r20_c9_2;
  wire [7:0] t_r20_c9_3;
  wire [7:0] t_r20_c9_4;
  wire [7:0] t_r20_c9_5;
  wire [7:0] t_r20_c9_6;
  wire [7:0] t_r20_c9_7;
  wire [7:0] t_r20_c9_8;
  wire [7:0] t_r20_c9_9;
  wire [7:0] t_r20_c9_10;
  wire [7:0] t_r20_c9_11;
  wire [7:0] t_r20_c9_12;
  wire [7:0] t_r20_c10_0;
  wire [7:0] t_r20_c10_1;
  wire [7:0] t_r20_c10_2;
  wire [7:0] t_r20_c10_3;
  wire [7:0] t_r20_c10_4;
  wire [7:0] t_r20_c10_5;
  wire [7:0] t_r20_c10_6;
  wire [7:0] t_r20_c10_7;
  wire [7:0] t_r20_c10_8;
  wire [7:0] t_r20_c10_9;
  wire [7:0] t_r20_c10_10;
  wire [7:0] t_r20_c10_11;
  wire [7:0] t_r20_c10_12;
  wire [7:0] t_r20_c11_0;
  wire [7:0] t_r20_c11_1;
  wire [7:0] t_r20_c11_2;
  wire [7:0] t_r20_c11_3;
  wire [7:0] t_r20_c11_4;
  wire [7:0] t_r20_c11_5;
  wire [7:0] t_r20_c11_6;
  wire [7:0] t_r20_c11_7;
  wire [7:0] t_r20_c11_8;
  wire [7:0] t_r20_c11_9;
  wire [7:0] t_r20_c11_10;
  wire [7:0] t_r20_c11_11;
  wire [7:0] t_r20_c11_12;
  wire [7:0] t_r20_c12_0;
  wire [7:0] t_r20_c12_1;
  wire [7:0] t_r20_c12_2;
  wire [7:0] t_r20_c12_3;
  wire [7:0] t_r20_c12_4;
  wire [7:0] t_r20_c12_5;
  wire [7:0] t_r20_c12_6;
  wire [7:0] t_r20_c12_7;
  wire [7:0] t_r20_c12_8;
  wire [7:0] t_r20_c12_9;
  wire [7:0] t_r20_c12_10;
  wire [7:0] t_r20_c12_11;
  wire [7:0] t_r20_c12_12;
  wire [7:0] t_r20_c13_0;
  wire [7:0] t_r20_c13_1;
  wire [7:0] t_r20_c13_2;
  wire [7:0] t_r20_c13_3;
  wire [7:0] t_r20_c13_4;
  wire [7:0] t_r20_c13_5;
  wire [7:0] t_r20_c13_6;
  wire [7:0] t_r20_c13_7;
  wire [7:0] t_r20_c13_8;
  wire [7:0] t_r20_c13_9;
  wire [7:0] t_r20_c13_10;
  wire [7:0] t_r20_c13_11;
  wire [7:0] t_r20_c13_12;
  wire [7:0] t_r20_c14_0;
  wire [7:0] t_r20_c14_1;
  wire [7:0] t_r20_c14_2;
  wire [7:0] t_r20_c14_3;
  wire [7:0] t_r20_c14_4;
  wire [7:0] t_r20_c14_5;
  wire [7:0] t_r20_c14_6;
  wire [7:0] t_r20_c14_7;
  wire [7:0] t_r20_c14_8;
  wire [7:0] t_r20_c14_9;
  wire [7:0] t_r20_c14_10;
  wire [7:0] t_r20_c14_11;
  wire [7:0] t_r20_c14_12;
  wire [7:0] t_r20_c15_0;
  wire [7:0] t_r20_c15_1;
  wire [7:0] t_r20_c15_2;
  wire [7:0] t_r20_c15_3;
  wire [7:0] t_r20_c15_4;
  wire [7:0] t_r20_c15_5;
  wire [7:0] t_r20_c15_6;
  wire [7:0] t_r20_c15_7;
  wire [7:0] t_r20_c15_8;
  wire [7:0] t_r20_c15_9;
  wire [7:0] t_r20_c15_10;
  wire [7:0] t_r20_c15_11;
  wire [7:0] t_r20_c15_12;
  wire [7:0] t_r20_c16_0;
  wire [7:0] t_r20_c16_1;
  wire [7:0] t_r20_c16_2;
  wire [7:0] t_r20_c16_3;
  wire [7:0] t_r20_c16_4;
  wire [7:0] t_r20_c16_5;
  wire [7:0] t_r20_c16_6;
  wire [7:0] t_r20_c16_7;
  wire [7:0] t_r20_c16_8;
  wire [7:0] t_r20_c16_9;
  wire [7:0] t_r20_c16_10;
  wire [7:0] t_r20_c16_11;
  wire [7:0] t_r20_c16_12;
  wire [7:0] t_r20_c17_0;
  wire [7:0] t_r20_c17_1;
  wire [7:0] t_r20_c17_2;
  wire [7:0] t_r20_c17_3;
  wire [7:0] t_r20_c17_4;
  wire [7:0] t_r20_c17_5;
  wire [7:0] t_r20_c17_6;
  wire [7:0] t_r20_c17_7;
  wire [7:0] t_r20_c17_8;
  wire [7:0] t_r20_c17_9;
  wire [7:0] t_r20_c17_10;
  wire [7:0] t_r20_c17_11;
  wire [7:0] t_r20_c17_12;
  wire [7:0] t_r20_c18_0;
  wire [7:0] t_r20_c18_1;
  wire [7:0] t_r20_c18_2;
  wire [7:0] t_r20_c18_3;
  wire [7:0] t_r20_c18_4;
  wire [7:0] t_r20_c18_5;
  wire [7:0] t_r20_c18_6;
  wire [7:0] t_r20_c18_7;
  wire [7:0] t_r20_c18_8;
  wire [7:0] t_r20_c18_9;
  wire [7:0] t_r20_c18_10;
  wire [7:0] t_r20_c18_11;
  wire [7:0] t_r20_c18_12;
  wire [7:0] t_r20_c19_0;
  wire [7:0] t_r20_c19_1;
  wire [7:0] t_r20_c19_2;
  wire [7:0] t_r20_c19_3;
  wire [7:0] t_r20_c19_4;
  wire [7:0] t_r20_c19_5;
  wire [7:0] t_r20_c19_6;
  wire [7:0] t_r20_c19_7;
  wire [7:0] t_r20_c19_8;
  wire [7:0] t_r20_c19_9;
  wire [7:0] t_r20_c19_10;
  wire [7:0] t_r20_c19_11;
  wire [7:0] t_r20_c19_12;
  wire [7:0] t_r20_c20_0;
  wire [7:0] t_r20_c20_1;
  wire [7:0] t_r20_c20_2;
  wire [7:0] t_r20_c20_3;
  wire [7:0] t_r20_c20_4;
  wire [7:0] t_r20_c20_5;
  wire [7:0] t_r20_c20_6;
  wire [7:0] t_r20_c20_7;
  wire [7:0] t_r20_c20_8;
  wire [7:0] t_r20_c20_9;
  wire [7:0] t_r20_c20_10;
  wire [7:0] t_r20_c20_11;
  wire [7:0] t_r20_c20_12;
  wire [7:0] t_r20_c21_0;
  wire [7:0] t_r20_c21_1;
  wire [7:0] t_r20_c21_2;
  wire [7:0] t_r20_c21_3;
  wire [7:0] t_r20_c21_4;
  wire [7:0] t_r20_c21_5;
  wire [7:0] t_r20_c21_6;
  wire [7:0] t_r20_c21_7;
  wire [7:0] t_r20_c21_8;
  wire [7:0] t_r20_c21_9;
  wire [7:0] t_r20_c21_10;
  wire [7:0] t_r20_c21_11;
  wire [7:0] t_r20_c21_12;
  wire [7:0] t_r20_c22_0;
  wire [7:0] t_r20_c22_1;
  wire [7:0] t_r20_c22_2;
  wire [7:0] t_r20_c22_3;
  wire [7:0] t_r20_c22_4;
  wire [7:0] t_r20_c22_5;
  wire [7:0] t_r20_c22_6;
  wire [7:0] t_r20_c22_7;
  wire [7:0] t_r20_c22_8;
  wire [7:0] t_r20_c22_9;
  wire [7:0] t_r20_c22_10;
  wire [7:0] t_r20_c22_11;
  wire [7:0] t_r20_c22_12;
  wire [7:0] t_r20_c23_0;
  wire [7:0] t_r20_c23_1;
  wire [7:0] t_r20_c23_2;
  wire [7:0] t_r20_c23_3;
  wire [7:0] t_r20_c23_4;
  wire [7:0] t_r20_c23_5;
  wire [7:0] t_r20_c23_6;
  wire [7:0] t_r20_c23_7;
  wire [7:0] t_r20_c23_8;
  wire [7:0] t_r20_c23_9;
  wire [7:0] t_r20_c23_10;
  wire [7:0] t_r20_c23_11;
  wire [7:0] t_r20_c23_12;
  wire [7:0] t_r20_c24_0;
  wire [7:0] t_r20_c24_1;
  wire [7:0] t_r20_c24_2;
  wire [7:0] t_r20_c24_3;
  wire [7:0] t_r20_c24_4;
  wire [7:0] t_r20_c24_5;
  wire [7:0] t_r20_c24_6;
  wire [7:0] t_r20_c24_7;
  wire [7:0] t_r20_c24_8;
  wire [7:0] t_r20_c24_9;
  wire [7:0] t_r20_c24_10;
  wire [7:0] t_r20_c24_11;
  wire [7:0] t_r20_c24_12;
  wire [7:0] t_r20_c25_0;
  wire [7:0] t_r20_c25_1;
  wire [7:0] t_r20_c25_2;
  wire [7:0] t_r20_c25_3;
  wire [7:0] t_r20_c25_4;
  wire [7:0] t_r20_c25_5;
  wire [7:0] t_r20_c25_6;
  wire [7:0] t_r20_c25_7;
  wire [7:0] t_r20_c25_8;
  wire [7:0] t_r20_c25_9;
  wire [7:0] t_r20_c25_10;
  wire [7:0] t_r20_c25_11;
  wire [7:0] t_r20_c25_12;
  wire [7:0] t_r20_c26_0;
  wire [7:0] t_r20_c26_1;
  wire [7:0] t_r20_c26_2;
  wire [7:0] t_r20_c26_3;
  wire [7:0] t_r20_c26_4;
  wire [7:0] t_r20_c26_5;
  wire [7:0] t_r20_c26_6;
  wire [7:0] t_r20_c26_7;
  wire [7:0] t_r20_c26_8;
  wire [7:0] t_r20_c26_9;
  wire [7:0] t_r20_c26_10;
  wire [7:0] t_r20_c26_11;
  wire [7:0] t_r20_c26_12;
  wire [7:0] t_r20_c27_0;
  wire [7:0] t_r20_c27_1;
  wire [7:0] t_r20_c27_2;
  wire [7:0] t_r20_c27_3;
  wire [7:0] t_r20_c27_4;
  wire [7:0] t_r20_c27_5;
  wire [7:0] t_r20_c27_6;
  wire [7:0] t_r20_c27_7;
  wire [7:0] t_r20_c27_8;
  wire [7:0] t_r20_c27_9;
  wire [7:0] t_r20_c27_10;
  wire [7:0] t_r20_c27_11;
  wire [7:0] t_r20_c27_12;
  wire [7:0] t_r20_c28_0;
  wire [7:0] t_r20_c28_1;
  wire [7:0] t_r20_c28_2;
  wire [7:0] t_r20_c28_3;
  wire [7:0] t_r20_c28_4;
  wire [7:0] t_r20_c28_5;
  wire [7:0] t_r20_c28_6;
  wire [7:0] t_r20_c28_7;
  wire [7:0] t_r20_c28_8;
  wire [7:0] t_r20_c28_9;
  wire [7:0] t_r20_c28_10;
  wire [7:0] t_r20_c28_11;
  wire [7:0] t_r20_c28_12;
  wire [7:0] t_r20_c29_0;
  wire [7:0] t_r20_c29_1;
  wire [7:0] t_r20_c29_2;
  wire [7:0] t_r20_c29_3;
  wire [7:0] t_r20_c29_4;
  wire [7:0] t_r20_c29_5;
  wire [7:0] t_r20_c29_6;
  wire [7:0] t_r20_c29_7;
  wire [7:0] t_r20_c29_8;
  wire [7:0] t_r20_c29_9;
  wire [7:0] t_r20_c29_10;
  wire [7:0] t_r20_c29_11;
  wire [7:0] t_r20_c29_12;
  wire [7:0] t_r20_c30_0;
  wire [7:0] t_r20_c30_1;
  wire [7:0] t_r20_c30_2;
  wire [7:0] t_r20_c30_3;
  wire [7:0] t_r20_c30_4;
  wire [7:0] t_r20_c30_5;
  wire [7:0] t_r20_c30_6;
  wire [7:0] t_r20_c30_7;
  wire [7:0] t_r20_c30_8;
  wire [7:0] t_r20_c30_9;
  wire [7:0] t_r20_c30_10;
  wire [7:0] t_r20_c30_11;
  wire [7:0] t_r20_c30_12;
  wire [7:0] t_r20_c31_0;
  wire [7:0] t_r20_c31_1;
  wire [7:0] t_r20_c31_2;
  wire [7:0] t_r20_c31_3;
  wire [7:0] t_r20_c31_4;
  wire [7:0] t_r20_c31_5;
  wire [7:0] t_r20_c31_6;
  wire [7:0] t_r20_c31_7;
  wire [7:0] t_r20_c31_8;
  wire [7:0] t_r20_c31_9;
  wire [7:0] t_r20_c31_10;
  wire [7:0] t_r20_c31_11;
  wire [7:0] t_r20_c31_12;
  wire [7:0] t_r20_c32_0;
  wire [7:0] t_r20_c32_1;
  wire [7:0] t_r20_c32_2;
  wire [7:0] t_r20_c32_3;
  wire [7:0] t_r20_c32_4;
  wire [7:0] t_r20_c32_5;
  wire [7:0] t_r20_c32_6;
  wire [7:0] t_r20_c32_7;
  wire [7:0] t_r20_c32_8;
  wire [7:0] t_r20_c32_9;
  wire [7:0] t_r20_c32_10;
  wire [7:0] t_r20_c32_11;
  wire [7:0] t_r20_c32_12;
  wire [7:0] t_r20_c33_0;
  wire [7:0] t_r20_c33_1;
  wire [7:0] t_r20_c33_2;
  wire [7:0] t_r20_c33_3;
  wire [7:0] t_r20_c33_4;
  wire [7:0] t_r20_c33_5;
  wire [7:0] t_r20_c33_6;
  wire [7:0] t_r20_c33_7;
  wire [7:0] t_r20_c33_8;
  wire [7:0] t_r20_c33_9;
  wire [7:0] t_r20_c33_10;
  wire [7:0] t_r20_c33_11;
  wire [7:0] t_r20_c33_12;
  wire [7:0] t_r20_c34_0;
  wire [7:0] t_r20_c34_1;
  wire [7:0] t_r20_c34_2;
  wire [7:0] t_r20_c34_3;
  wire [7:0] t_r20_c34_4;
  wire [7:0] t_r20_c34_5;
  wire [7:0] t_r20_c34_6;
  wire [7:0] t_r20_c34_7;
  wire [7:0] t_r20_c34_8;
  wire [7:0] t_r20_c34_9;
  wire [7:0] t_r20_c34_10;
  wire [7:0] t_r20_c34_11;
  wire [7:0] t_r20_c34_12;
  wire [7:0] t_r20_c35_0;
  wire [7:0] t_r20_c35_1;
  wire [7:0] t_r20_c35_2;
  wire [7:0] t_r20_c35_3;
  wire [7:0] t_r20_c35_4;
  wire [7:0] t_r20_c35_5;
  wire [7:0] t_r20_c35_6;
  wire [7:0] t_r20_c35_7;
  wire [7:0] t_r20_c35_8;
  wire [7:0] t_r20_c35_9;
  wire [7:0] t_r20_c35_10;
  wire [7:0] t_r20_c35_11;
  wire [7:0] t_r20_c35_12;
  wire [7:0] t_r20_c36_0;
  wire [7:0] t_r20_c36_1;
  wire [7:0] t_r20_c36_2;
  wire [7:0] t_r20_c36_3;
  wire [7:0] t_r20_c36_4;
  wire [7:0] t_r20_c36_5;
  wire [7:0] t_r20_c36_6;
  wire [7:0] t_r20_c36_7;
  wire [7:0] t_r20_c36_8;
  wire [7:0] t_r20_c36_9;
  wire [7:0] t_r20_c36_10;
  wire [7:0] t_r20_c36_11;
  wire [7:0] t_r20_c36_12;
  wire [7:0] t_r20_c37_0;
  wire [7:0] t_r20_c37_1;
  wire [7:0] t_r20_c37_2;
  wire [7:0] t_r20_c37_3;
  wire [7:0] t_r20_c37_4;
  wire [7:0] t_r20_c37_5;
  wire [7:0] t_r20_c37_6;
  wire [7:0] t_r20_c37_7;
  wire [7:0] t_r20_c37_8;
  wire [7:0] t_r20_c37_9;
  wire [7:0] t_r20_c37_10;
  wire [7:0] t_r20_c37_11;
  wire [7:0] t_r20_c37_12;
  wire [7:0] t_r20_c38_0;
  wire [7:0] t_r20_c38_1;
  wire [7:0] t_r20_c38_2;
  wire [7:0] t_r20_c38_3;
  wire [7:0] t_r20_c38_4;
  wire [7:0] t_r20_c38_5;
  wire [7:0] t_r20_c38_6;
  wire [7:0] t_r20_c38_7;
  wire [7:0] t_r20_c38_8;
  wire [7:0] t_r20_c38_9;
  wire [7:0] t_r20_c38_10;
  wire [7:0] t_r20_c38_11;
  wire [7:0] t_r20_c38_12;
  wire [7:0] t_r20_c39_0;
  wire [7:0] t_r20_c39_1;
  wire [7:0] t_r20_c39_2;
  wire [7:0] t_r20_c39_3;
  wire [7:0] t_r20_c39_4;
  wire [7:0] t_r20_c39_5;
  wire [7:0] t_r20_c39_6;
  wire [7:0] t_r20_c39_7;
  wire [7:0] t_r20_c39_8;
  wire [7:0] t_r20_c39_9;
  wire [7:0] t_r20_c39_10;
  wire [7:0] t_r20_c39_11;
  wire [7:0] t_r20_c39_12;
  wire [7:0] t_r20_c40_0;
  wire [7:0] t_r20_c40_1;
  wire [7:0] t_r20_c40_2;
  wire [7:0] t_r20_c40_3;
  wire [7:0] t_r20_c40_4;
  wire [7:0] t_r20_c40_5;
  wire [7:0] t_r20_c40_6;
  wire [7:0] t_r20_c40_7;
  wire [7:0] t_r20_c40_8;
  wire [7:0] t_r20_c40_9;
  wire [7:0] t_r20_c40_10;
  wire [7:0] t_r20_c40_11;
  wire [7:0] t_r20_c40_12;
  wire [7:0] t_r20_c41_0;
  wire [7:0] t_r20_c41_1;
  wire [7:0] t_r20_c41_2;
  wire [7:0] t_r20_c41_3;
  wire [7:0] t_r20_c41_4;
  wire [7:0] t_r20_c41_5;
  wire [7:0] t_r20_c41_6;
  wire [7:0] t_r20_c41_7;
  wire [7:0] t_r20_c41_8;
  wire [7:0] t_r20_c41_9;
  wire [7:0] t_r20_c41_10;
  wire [7:0] t_r20_c41_11;
  wire [7:0] t_r20_c41_12;
  wire [7:0] t_r20_c42_0;
  wire [7:0] t_r20_c42_1;
  wire [7:0] t_r20_c42_2;
  wire [7:0] t_r20_c42_3;
  wire [7:0] t_r20_c42_4;
  wire [7:0] t_r20_c42_5;
  wire [7:0] t_r20_c42_6;
  wire [7:0] t_r20_c42_7;
  wire [7:0] t_r20_c42_8;
  wire [7:0] t_r20_c42_9;
  wire [7:0] t_r20_c42_10;
  wire [7:0] t_r20_c42_11;
  wire [7:0] t_r20_c42_12;
  wire [7:0] t_r20_c43_0;
  wire [7:0] t_r20_c43_1;
  wire [7:0] t_r20_c43_2;
  wire [7:0] t_r20_c43_3;
  wire [7:0] t_r20_c43_4;
  wire [7:0] t_r20_c43_5;
  wire [7:0] t_r20_c43_6;
  wire [7:0] t_r20_c43_7;
  wire [7:0] t_r20_c43_8;
  wire [7:0] t_r20_c43_9;
  wire [7:0] t_r20_c43_10;
  wire [7:0] t_r20_c43_11;
  wire [7:0] t_r20_c43_12;
  wire [7:0] t_r20_c44_0;
  wire [7:0] t_r20_c44_1;
  wire [7:0] t_r20_c44_2;
  wire [7:0] t_r20_c44_3;
  wire [7:0] t_r20_c44_4;
  wire [7:0] t_r20_c44_5;
  wire [7:0] t_r20_c44_6;
  wire [7:0] t_r20_c44_7;
  wire [7:0] t_r20_c44_8;
  wire [7:0] t_r20_c44_9;
  wire [7:0] t_r20_c44_10;
  wire [7:0] t_r20_c44_11;
  wire [7:0] t_r20_c44_12;
  wire [7:0] t_r20_c45_0;
  wire [7:0] t_r20_c45_1;
  wire [7:0] t_r20_c45_2;
  wire [7:0] t_r20_c45_3;
  wire [7:0] t_r20_c45_4;
  wire [7:0] t_r20_c45_5;
  wire [7:0] t_r20_c45_6;
  wire [7:0] t_r20_c45_7;
  wire [7:0] t_r20_c45_8;
  wire [7:0] t_r20_c45_9;
  wire [7:0] t_r20_c45_10;
  wire [7:0] t_r20_c45_11;
  wire [7:0] t_r20_c45_12;
  wire [7:0] t_r20_c46_0;
  wire [7:0] t_r20_c46_1;
  wire [7:0] t_r20_c46_2;
  wire [7:0] t_r20_c46_3;
  wire [7:0] t_r20_c46_4;
  wire [7:0] t_r20_c46_5;
  wire [7:0] t_r20_c46_6;
  wire [7:0] t_r20_c46_7;
  wire [7:0] t_r20_c46_8;
  wire [7:0] t_r20_c46_9;
  wire [7:0] t_r20_c46_10;
  wire [7:0] t_r20_c46_11;
  wire [7:0] t_r20_c46_12;
  wire [7:0] t_r20_c47_0;
  wire [7:0] t_r20_c47_1;
  wire [7:0] t_r20_c47_2;
  wire [7:0] t_r20_c47_3;
  wire [7:0] t_r20_c47_4;
  wire [7:0] t_r20_c47_5;
  wire [7:0] t_r20_c47_6;
  wire [7:0] t_r20_c47_7;
  wire [7:0] t_r20_c47_8;
  wire [7:0] t_r20_c47_9;
  wire [7:0] t_r20_c47_10;
  wire [7:0] t_r20_c47_11;
  wire [7:0] t_r20_c47_12;
  wire [7:0] t_r20_c48_0;
  wire [7:0] t_r20_c48_1;
  wire [7:0] t_r20_c48_2;
  wire [7:0] t_r20_c48_3;
  wire [7:0] t_r20_c48_4;
  wire [7:0] t_r20_c48_5;
  wire [7:0] t_r20_c48_6;
  wire [7:0] t_r20_c48_7;
  wire [7:0] t_r20_c48_8;
  wire [7:0] t_r20_c48_9;
  wire [7:0] t_r20_c48_10;
  wire [7:0] t_r20_c48_11;
  wire [7:0] t_r20_c48_12;
  wire [7:0] t_r20_c49_0;
  wire [7:0] t_r20_c49_1;
  wire [7:0] t_r20_c49_2;
  wire [7:0] t_r20_c49_3;
  wire [7:0] t_r20_c49_4;
  wire [7:0] t_r20_c49_5;
  wire [7:0] t_r20_c49_6;
  wire [7:0] t_r20_c49_7;
  wire [7:0] t_r20_c49_8;
  wire [7:0] t_r20_c49_9;
  wire [7:0] t_r20_c49_10;
  wire [7:0] t_r20_c49_11;
  wire [7:0] t_r20_c49_12;
  wire [7:0] t_r20_c50_0;
  wire [7:0] t_r20_c50_1;
  wire [7:0] t_r20_c50_2;
  wire [7:0] t_r20_c50_3;
  wire [7:0] t_r20_c50_4;
  wire [7:0] t_r20_c50_5;
  wire [7:0] t_r20_c50_6;
  wire [7:0] t_r20_c50_7;
  wire [7:0] t_r20_c50_8;
  wire [7:0] t_r20_c50_9;
  wire [7:0] t_r20_c50_10;
  wire [7:0] t_r20_c50_11;
  wire [7:0] t_r20_c50_12;
  wire [7:0] t_r20_c51_0;
  wire [7:0] t_r20_c51_1;
  wire [7:0] t_r20_c51_2;
  wire [7:0] t_r20_c51_3;
  wire [7:0] t_r20_c51_4;
  wire [7:0] t_r20_c51_5;
  wire [7:0] t_r20_c51_6;
  wire [7:0] t_r20_c51_7;
  wire [7:0] t_r20_c51_8;
  wire [7:0] t_r20_c51_9;
  wire [7:0] t_r20_c51_10;
  wire [7:0] t_r20_c51_11;
  wire [7:0] t_r20_c51_12;
  wire [7:0] t_r20_c52_0;
  wire [7:0] t_r20_c52_1;
  wire [7:0] t_r20_c52_2;
  wire [7:0] t_r20_c52_3;
  wire [7:0] t_r20_c52_4;
  wire [7:0] t_r20_c52_5;
  wire [7:0] t_r20_c52_6;
  wire [7:0] t_r20_c52_7;
  wire [7:0] t_r20_c52_8;
  wire [7:0] t_r20_c52_9;
  wire [7:0] t_r20_c52_10;
  wire [7:0] t_r20_c52_11;
  wire [7:0] t_r20_c52_12;
  wire [7:0] t_r20_c53_0;
  wire [7:0] t_r20_c53_1;
  wire [7:0] t_r20_c53_2;
  wire [7:0] t_r20_c53_3;
  wire [7:0] t_r20_c53_4;
  wire [7:0] t_r20_c53_5;
  wire [7:0] t_r20_c53_6;
  wire [7:0] t_r20_c53_7;
  wire [7:0] t_r20_c53_8;
  wire [7:0] t_r20_c53_9;
  wire [7:0] t_r20_c53_10;
  wire [7:0] t_r20_c53_11;
  wire [7:0] t_r20_c53_12;
  wire [7:0] t_r20_c54_0;
  wire [7:0] t_r20_c54_1;
  wire [7:0] t_r20_c54_2;
  wire [7:0] t_r20_c54_3;
  wire [7:0] t_r20_c54_4;
  wire [7:0] t_r20_c54_5;
  wire [7:0] t_r20_c54_6;
  wire [7:0] t_r20_c54_7;
  wire [7:0] t_r20_c54_8;
  wire [7:0] t_r20_c54_9;
  wire [7:0] t_r20_c54_10;
  wire [7:0] t_r20_c54_11;
  wire [7:0] t_r20_c54_12;
  wire [7:0] t_r20_c55_0;
  wire [7:0] t_r20_c55_1;
  wire [7:0] t_r20_c55_2;
  wire [7:0] t_r20_c55_3;
  wire [7:0] t_r20_c55_4;
  wire [7:0] t_r20_c55_5;
  wire [7:0] t_r20_c55_6;
  wire [7:0] t_r20_c55_7;
  wire [7:0] t_r20_c55_8;
  wire [7:0] t_r20_c55_9;
  wire [7:0] t_r20_c55_10;
  wire [7:0] t_r20_c55_11;
  wire [7:0] t_r20_c55_12;
  wire [7:0] t_r20_c56_0;
  wire [7:0] t_r20_c56_1;
  wire [7:0] t_r20_c56_2;
  wire [7:0] t_r20_c56_3;
  wire [7:0] t_r20_c56_4;
  wire [7:0] t_r20_c56_5;
  wire [7:0] t_r20_c56_6;
  wire [7:0] t_r20_c56_7;
  wire [7:0] t_r20_c56_8;
  wire [7:0] t_r20_c56_9;
  wire [7:0] t_r20_c56_10;
  wire [7:0] t_r20_c56_11;
  wire [7:0] t_r20_c56_12;
  wire [7:0] t_r20_c57_0;
  wire [7:0] t_r20_c57_1;
  wire [7:0] t_r20_c57_2;
  wire [7:0] t_r20_c57_3;
  wire [7:0] t_r20_c57_4;
  wire [7:0] t_r20_c57_5;
  wire [7:0] t_r20_c57_6;
  wire [7:0] t_r20_c57_7;
  wire [7:0] t_r20_c57_8;
  wire [7:0] t_r20_c57_9;
  wire [7:0] t_r20_c57_10;
  wire [7:0] t_r20_c57_11;
  wire [7:0] t_r20_c57_12;
  wire [7:0] t_r20_c58_0;
  wire [7:0] t_r20_c58_1;
  wire [7:0] t_r20_c58_2;
  wire [7:0] t_r20_c58_3;
  wire [7:0] t_r20_c58_4;
  wire [7:0] t_r20_c58_5;
  wire [7:0] t_r20_c58_6;
  wire [7:0] t_r20_c58_7;
  wire [7:0] t_r20_c58_8;
  wire [7:0] t_r20_c58_9;
  wire [7:0] t_r20_c58_10;
  wire [7:0] t_r20_c58_11;
  wire [7:0] t_r20_c58_12;
  wire [7:0] t_r20_c59_0;
  wire [7:0] t_r20_c59_1;
  wire [7:0] t_r20_c59_2;
  wire [7:0] t_r20_c59_3;
  wire [7:0] t_r20_c59_4;
  wire [7:0] t_r20_c59_5;
  wire [7:0] t_r20_c59_6;
  wire [7:0] t_r20_c59_7;
  wire [7:0] t_r20_c59_8;
  wire [7:0] t_r20_c59_9;
  wire [7:0] t_r20_c59_10;
  wire [7:0] t_r20_c59_11;
  wire [7:0] t_r20_c59_12;
  wire [7:0] t_r20_c60_0;
  wire [7:0] t_r20_c60_1;
  wire [7:0] t_r20_c60_2;
  wire [7:0] t_r20_c60_3;
  wire [7:0] t_r20_c60_4;
  wire [7:0] t_r20_c60_5;
  wire [7:0] t_r20_c60_6;
  wire [7:0] t_r20_c60_7;
  wire [7:0] t_r20_c60_8;
  wire [7:0] t_r20_c60_9;
  wire [7:0] t_r20_c60_10;
  wire [7:0] t_r20_c60_11;
  wire [7:0] t_r20_c60_12;
  wire [7:0] t_r20_c61_0;
  wire [7:0] t_r20_c61_1;
  wire [7:0] t_r20_c61_2;
  wire [7:0] t_r20_c61_3;
  wire [7:0] t_r20_c61_4;
  wire [7:0] t_r20_c61_5;
  wire [7:0] t_r20_c61_6;
  wire [7:0] t_r20_c61_7;
  wire [7:0] t_r20_c61_8;
  wire [7:0] t_r20_c61_9;
  wire [7:0] t_r20_c61_10;
  wire [7:0] t_r20_c61_11;
  wire [7:0] t_r20_c61_12;
  wire [7:0] t_r20_c62_0;
  wire [7:0] t_r20_c62_1;
  wire [7:0] t_r20_c62_2;
  wire [7:0] t_r20_c62_3;
  wire [7:0] t_r20_c62_4;
  wire [7:0] t_r20_c62_5;
  wire [7:0] t_r20_c62_6;
  wire [7:0] t_r20_c62_7;
  wire [7:0] t_r20_c62_8;
  wire [7:0] t_r20_c62_9;
  wire [7:0] t_r20_c62_10;
  wire [7:0] t_r20_c62_11;
  wire [7:0] t_r20_c62_12;
  wire [7:0] t_r20_c63_0;
  wire [7:0] t_r20_c63_1;
  wire [7:0] t_r20_c63_2;
  wire [7:0] t_r20_c63_3;
  wire [7:0] t_r20_c63_4;
  wire [7:0] t_r20_c63_5;
  wire [7:0] t_r20_c63_6;
  wire [7:0] t_r20_c63_7;
  wire [7:0] t_r20_c63_8;
  wire [7:0] t_r20_c63_9;
  wire [7:0] t_r20_c63_10;
  wire [7:0] t_r20_c63_11;
  wire [7:0] t_r20_c63_12;
  wire [7:0] t_r20_c64_0;
  wire [7:0] t_r20_c64_1;
  wire [7:0] t_r20_c64_2;
  wire [7:0] t_r20_c64_3;
  wire [7:0] t_r20_c64_4;
  wire [7:0] t_r20_c64_5;
  wire [7:0] t_r20_c64_6;
  wire [7:0] t_r20_c64_7;
  wire [7:0] t_r20_c64_8;
  wire [7:0] t_r20_c64_9;
  wire [7:0] t_r20_c64_10;
  wire [7:0] t_r20_c64_11;
  wire [7:0] t_r20_c64_12;
  wire [7:0] t_r20_c65_0;
  wire [7:0] t_r20_c65_1;
  wire [7:0] t_r20_c65_2;
  wire [7:0] t_r20_c65_3;
  wire [7:0] t_r20_c65_4;
  wire [7:0] t_r20_c65_5;
  wire [7:0] t_r20_c65_6;
  wire [7:0] t_r20_c65_7;
  wire [7:0] t_r20_c65_8;
  wire [7:0] t_r20_c65_9;
  wire [7:0] t_r20_c65_10;
  wire [7:0] t_r20_c65_11;
  wire [7:0] t_r20_c65_12;
  wire [7:0] t_r21_c0_0;
  wire [7:0] t_r21_c0_1;
  wire [7:0] t_r21_c0_2;
  wire [7:0] t_r21_c0_3;
  wire [7:0] t_r21_c0_4;
  wire [7:0] t_r21_c0_5;
  wire [7:0] t_r21_c0_6;
  wire [7:0] t_r21_c0_7;
  wire [7:0] t_r21_c0_8;
  wire [7:0] t_r21_c0_9;
  wire [7:0] t_r21_c0_10;
  wire [7:0] t_r21_c0_11;
  wire [7:0] t_r21_c0_12;
  wire [7:0] t_r21_c1_0;
  wire [7:0] t_r21_c1_1;
  wire [7:0] t_r21_c1_2;
  wire [7:0] t_r21_c1_3;
  wire [7:0] t_r21_c1_4;
  wire [7:0] t_r21_c1_5;
  wire [7:0] t_r21_c1_6;
  wire [7:0] t_r21_c1_7;
  wire [7:0] t_r21_c1_8;
  wire [7:0] t_r21_c1_9;
  wire [7:0] t_r21_c1_10;
  wire [7:0] t_r21_c1_11;
  wire [7:0] t_r21_c1_12;
  wire [7:0] t_r21_c2_0;
  wire [7:0] t_r21_c2_1;
  wire [7:0] t_r21_c2_2;
  wire [7:0] t_r21_c2_3;
  wire [7:0] t_r21_c2_4;
  wire [7:0] t_r21_c2_5;
  wire [7:0] t_r21_c2_6;
  wire [7:0] t_r21_c2_7;
  wire [7:0] t_r21_c2_8;
  wire [7:0] t_r21_c2_9;
  wire [7:0] t_r21_c2_10;
  wire [7:0] t_r21_c2_11;
  wire [7:0] t_r21_c2_12;
  wire [7:0] t_r21_c3_0;
  wire [7:0] t_r21_c3_1;
  wire [7:0] t_r21_c3_2;
  wire [7:0] t_r21_c3_3;
  wire [7:0] t_r21_c3_4;
  wire [7:0] t_r21_c3_5;
  wire [7:0] t_r21_c3_6;
  wire [7:0] t_r21_c3_7;
  wire [7:0] t_r21_c3_8;
  wire [7:0] t_r21_c3_9;
  wire [7:0] t_r21_c3_10;
  wire [7:0] t_r21_c3_11;
  wire [7:0] t_r21_c3_12;
  wire [7:0] t_r21_c4_0;
  wire [7:0] t_r21_c4_1;
  wire [7:0] t_r21_c4_2;
  wire [7:0] t_r21_c4_3;
  wire [7:0] t_r21_c4_4;
  wire [7:0] t_r21_c4_5;
  wire [7:0] t_r21_c4_6;
  wire [7:0] t_r21_c4_7;
  wire [7:0] t_r21_c4_8;
  wire [7:0] t_r21_c4_9;
  wire [7:0] t_r21_c4_10;
  wire [7:0] t_r21_c4_11;
  wire [7:0] t_r21_c4_12;
  wire [7:0] t_r21_c5_0;
  wire [7:0] t_r21_c5_1;
  wire [7:0] t_r21_c5_2;
  wire [7:0] t_r21_c5_3;
  wire [7:0] t_r21_c5_4;
  wire [7:0] t_r21_c5_5;
  wire [7:0] t_r21_c5_6;
  wire [7:0] t_r21_c5_7;
  wire [7:0] t_r21_c5_8;
  wire [7:0] t_r21_c5_9;
  wire [7:0] t_r21_c5_10;
  wire [7:0] t_r21_c5_11;
  wire [7:0] t_r21_c5_12;
  wire [7:0] t_r21_c6_0;
  wire [7:0] t_r21_c6_1;
  wire [7:0] t_r21_c6_2;
  wire [7:0] t_r21_c6_3;
  wire [7:0] t_r21_c6_4;
  wire [7:0] t_r21_c6_5;
  wire [7:0] t_r21_c6_6;
  wire [7:0] t_r21_c6_7;
  wire [7:0] t_r21_c6_8;
  wire [7:0] t_r21_c6_9;
  wire [7:0] t_r21_c6_10;
  wire [7:0] t_r21_c6_11;
  wire [7:0] t_r21_c6_12;
  wire [7:0] t_r21_c7_0;
  wire [7:0] t_r21_c7_1;
  wire [7:0] t_r21_c7_2;
  wire [7:0] t_r21_c7_3;
  wire [7:0] t_r21_c7_4;
  wire [7:0] t_r21_c7_5;
  wire [7:0] t_r21_c7_6;
  wire [7:0] t_r21_c7_7;
  wire [7:0] t_r21_c7_8;
  wire [7:0] t_r21_c7_9;
  wire [7:0] t_r21_c7_10;
  wire [7:0] t_r21_c7_11;
  wire [7:0] t_r21_c7_12;
  wire [7:0] t_r21_c8_0;
  wire [7:0] t_r21_c8_1;
  wire [7:0] t_r21_c8_2;
  wire [7:0] t_r21_c8_3;
  wire [7:0] t_r21_c8_4;
  wire [7:0] t_r21_c8_5;
  wire [7:0] t_r21_c8_6;
  wire [7:0] t_r21_c8_7;
  wire [7:0] t_r21_c8_8;
  wire [7:0] t_r21_c8_9;
  wire [7:0] t_r21_c8_10;
  wire [7:0] t_r21_c8_11;
  wire [7:0] t_r21_c8_12;
  wire [7:0] t_r21_c9_0;
  wire [7:0] t_r21_c9_1;
  wire [7:0] t_r21_c9_2;
  wire [7:0] t_r21_c9_3;
  wire [7:0] t_r21_c9_4;
  wire [7:0] t_r21_c9_5;
  wire [7:0] t_r21_c9_6;
  wire [7:0] t_r21_c9_7;
  wire [7:0] t_r21_c9_8;
  wire [7:0] t_r21_c9_9;
  wire [7:0] t_r21_c9_10;
  wire [7:0] t_r21_c9_11;
  wire [7:0] t_r21_c9_12;
  wire [7:0] t_r21_c10_0;
  wire [7:0] t_r21_c10_1;
  wire [7:0] t_r21_c10_2;
  wire [7:0] t_r21_c10_3;
  wire [7:0] t_r21_c10_4;
  wire [7:0] t_r21_c10_5;
  wire [7:0] t_r21_c10_6;
  wire [7:0] t_r21_c10_7;
  wire [7:0] t_r21_c10_8;
  wire [7:0] t_r21_c10_9;
  wire [7:0] t_r21_c10_10;
  wire [7:0] t_r21_c10_11;
  wire [7:0] t_r21_c10_12;
  wire [7:0] t_r21_c11_0;
  wire [7:0] t_r21_c11_1;
  wire [7:0] t_r21_c11_2;
  wire [7:0] t_r21_c11_3;
  wire [7:0] t_r21_c11_4;
  wire [7:0] t_r21_c11_5;
  wire [7:0] t_r21_c11_6;
  wire [7:0] t_r21_c11_7;
  wire [7:0] t_r21_c11_8;
  wire [7:0] t_r21_c11_9;
  wire [7:0] t_r21_c11_10;
  wire [7:0] t_r21_c11_11;
  wire [7:0] t_r21_c11_12;
  wire [7:0] t_r21_c12_0;
  wire [7:0] t_r21_c12_1;
  wire [7:0] t_r21_c12_2;
  wire [7:0] t_r21_c12_3;
  wire [7:0] t_r21_c12_4;
  wire [7:0] t_r21_c12_5;
  wire [7:0] t_r21_c12_6;
  wire [7:0] t_r21_c12_7;
  wire [7:0] t_r21_c12_8;
  wire [7:0] t_r21_c12_9;
  wire [7:0] t_r21_c12_10;
  wire [7:0] t_r21_c12_11;
  wire [7:0] t_r21_c12_12;
  wire [7:0] t_r21_c13_0;
  wire [7:0] t_r21_c13_1;
  wire [7:0] t_r21_c13_2;
  wire [7:0] t_r21_c13_3;
  wire [7:0] t_r21_c13_4;
  wire [7:0] t_r21_c13_5;
  wire [7:0] t_r21_c13_6;
  wire [7:0] t_r21_c13_7;
  wire [7:0] t_r21_c13_8;
  wire [7:0] t_r21_c13_9;
  wire [7:0] t_r21_c13_10;
  wire [7:0] t_r21_c13_11;
  wire [7:0] t_r21_c13_12;
  wire [7:0] t_r21_c14_0;
  wire [7:0] t_r21_c14_1;
  wire [7:0] t_r21_c14_2;
  wire [7:0] t_r21_c14_3;
  wire [7:0] t_r21_c14_4;
  wire [7:0] t_r21_c14_5;
  wire [7:0] t_r21_c14_6;
  wire [7:0] t_r21_c14_7;
  wire [7:0] t_r21_c14_8;
  wire [7:0] t_r21_c14_9;
  wire [7:0] t_r21_c14_10;
  wire [7:0] t_r21_c14_11;
  wire [7:0] t_r21_c14_12;
  wire [7:0] t_r21_c15_0;
  wire [7:0] t_r21_c15_1;
  wire [7:0] t_r21_c15_2;
  wire [7:0] t_r21_c15_3;
  wire [7:0] t_r21_c15_4;
  wire [7:0] t_r21_c15_5;
  wire [7:0] t_r21_c15_6;
  wire [7:0] t_r21_c15_7;
  wire [7:0] t_r21_c15_8;
  wire [7:0] t_r21_c15_9;
  wire [7:0] t_r21_c15_10;
  wire [7:0] t_r21_c15_11;
  wire [7:0] t_r21_c15_12;
  wire [7:0] t_r21_c16_0;
  wire [7:0] t_r21_c16_1;
  wire [7:0] t_r21_c16_2;
  wire [7:0] t_r21_c16_3;
  wire [7:0] t_r21_c16_4;
  wire [7:0] t_r21_c16_5;
  wire [7:0] t_r21_c16_6;
  wire [7:0] t_r21_c16_7;
  wire [7:0] t_r21_c16_8;
  wire [7:0] t_r21_c16_9;
  wire [7:0] t_r21_c16_10;
  wire [7:0] t_r21_c16_11;
  wire [7:0] t_r21_c16_12;
  wire [7:0] t_r21_c17_0;
  wire [7:0] t_r21_c17_1;
  wire [7:0] t_r21_c17_2;
  wire [7:0] t_r21_c17_3;
  wire [7:0] t_r21_c17_4;
  wire [7:0] t_r21_c17_5;
  wire [7:0] t_r21_c17_6;
  wire [7:0] t_r21_c17_7;
  wire [7:0] t_r21_c17_8;
  wire [7:0] t_r21_c17_9;
  wire [7:0] t_r21_c17_10;
  wire [7:0] t_r21_c17_11;
  wire [7:0] t_r21_c17_12;
  wire [7:0] t_r21_c18_0;
  wire [7:0] t_r21_c18_1;
  wire [7:0] t_r21_c18_2;
  wire [7:0] t_r21_c18_3;
  wire [7:0] t_r21_c18_4;
  wire [7:0] t_r21_c18_5;
  wire [7:0] t_r21_c18_6;
  wire [7:0] t_r21_c18_7;
  wire [7:0] t_r21_c18_8;
  wire [7:0] t_r21_c18_9;
  wire [7:0] t_r21_c18_10;
  wire [7:0] t_r21_c18_11;
  wire [7:0] t_r21_c18_12;
  wire [7:0] t_r21_c19_0;
  wire [7:0] t_r21_c19_1;
  wire [7:0] t_r21_c19_2;
  wire [7:0] t_r21_c19_3;
  wire [7:0] t_r21_c19_4;
  wire [7:0] t_r21_c19_5;
  wire [7:0] t_r21_c19_6;
  wire [7:0] t_r21_c19_7;
  wire [7:0] t_r21_c19_8;
  wire [7:0] t_r21_c19_9;
  wire [7:0] t_r21_c19_10;
  wire [7:0] t_r21_c19_11;
  wire [7:0] t_r21_c19_12;
  wire [7:0] t_r21_c20_0;
  wire [7:0] t_r21_c20_1;
  wire [7:0] t_r21_c20_2;
  wire [7:0] t_r21_c20_3;
  wire [7:0] t_r21_c20_4;
  wire [7:0] t_r21_c20_5;
  wire [7:0] t_r21_c20_6;
  wire [7:0] t_r21_c20_7;
  wire [7:0] t_r21_c20_8;
  wire [7:0] t_r21_c20_9;
  wire [7:0] t_r21_c20_10;
  wire [7:0] t_r21_c20_11;
  wire [7:0] t_r21_c20_12;
  wire [7:0] t_r21_c21_0;
  wire [7:0] t_r21_c21_1;
  wire [7:0] t_r21_c21_2;
  wire [7:0] t_r21_c21_3;
  wire [7:0] t_r21_c21_4;
  wire [7:0] t_r21_c21_5;
  wire [7:0] t_r21_c21_6;
  wire [7:0] t_r21_c21_7;
  wire [7:0] t_r21_c21_8;
  wire [7:0] t_r21_c21_9;
  wire [7:0] t_r21_c21_10;
  wire [7:0] t_r21_c21_11;
  wire [7:0] t_r21_c21_12;
  wire [7:0] t_r21_c22_0;
  wire [7:0] t_r21_c22_1;
  wire [7:0] t_r21_c22_2;
  wire [7:0] t_r21_c22_3;
  wire [7:0] t_r21_c22_4;
  wire [7:0] t_r21_c22_5;
  wire [7:0] t_r21_c22_6;
  wire [7:0] t_r21_c22_7;
  wire [7:0] t_r21_c22_8;
  wire [7:0] t_r21_c22_9;
  wire [7:0] t_r21_c22_10;
  wire [7:0] t_r21_c22_11;
  wire [7:0] t_r21_c22_12;
  wire [7:0] t_r21_c23_0;
  wire [7:0] t_r21_c23_1;
  wire [7:0] t_r21_c23_2;
  wire [7:0] t_r21_c23_3;
  wire [7:0] t_r21_c23_4;
  wire [7:0] t_r21_c23_5;
  wire [7:0] t_r21_c23_6;
  wire [7:0] t_r21_c23_7;
  wire [7:0] t_r21_c23_8;
  wire [7:0] t_r21_c23_9;
  wire [7:0] t_r21_c23_10;
  wire [7:0] t_r21_c23_11;
  wire [7:0] t_r21_c23_12;
  wire [7:0] t_r21_c24_0;
  wire [7:0] t_r21_c24_1;
  wire [7:0] t_r21_c24_2;
  wire [7:0] t_r21_c24_3;
  wire [7:0] t_r21_c24_4;
  wire [7:0] t_r21_c24_5;
  wire [7:0] t_r21_c24_6;
  wire [7:0] t_r21_c24_7;
  wire [7:0] t_r21_c24_8;
  wire [7:0] t_r21_c24_9;
  wire [7:0] t_r21_c24_10;
  wire [7:0] t_r21_c24_11;
  wire [7:0] t_r21_c24_12;
  wire [7:0] t_r21_c25_0;
  wire [7:0] t_r21_c25_1;
  wire [7:0] t_r21_c25_2;
  wire [7:0] t_r21_c25_3;
  wire [7:0] t_r21_c25_4;
  wire [7:0] t_r21_c25_5;
  wire [7:0] t_r21_c25_6;
  wire [7:0] t_r21_c25_7;
  wire [7:0] t_r21_c25_8;
  wire [7:0] t_r21_c25_9;
  wire [7:0] t_r21_c25_10;
  wire [7:0] t_r21_c25_11;
  wire [7:0] t_r21_c25_12;
  wire [7:0] t_r21_c26_0;
  wire [7:0] t_r21_c26_1;
  wire [7:0] t_r21_c26_2;
  wire [7:0] t_r21_c26_3;
  wire [7:0] t_r21_c26_4;
  wire [7:0] t_r21_c26_5;
  wire [7:0] t_r21_c26_6;
  wire [7:0] t_r21_c26_7;
  wire [7:0] t_r21_c26_8;
  wire [7:0] t_r21_c26_9;
  wire [7:0] t_r21_c26_10;
  wire [7:0] t_r21_c26_11;
  wire [7:0] t_r21_c26_12;
  wire [7:0] t_r21_c27_0;
  wire [7:0] t_r21_c27_1;
  wire [7:0] t_r21_c27_2;
  wire [7:0] t_r21_c27_3;
  wire [7:0] t_r21_c27_4;
  wire [7:0] t_r21_c27_5;
  wire [7:0] t_r21_c27_6;
  wire [7:0] t_r21_c27_7;
  wire [7:0] t_r21_c27_8;
  wire [7:0] t_r21_c27_9;
  wire [7:0] t_r21_c27_10;
  wire [7:0] t_r21_c27_11;
  wire [7:0] t_r21_c27_12;
  wire [7:0] t_r21_c28_0;
  wire [7:0] t_r21_c28_1;
  wire [7:0] t_r21_c28_2;
  wire [7:0] t_r21_c28_3;
  wire [7:0] t_r21_c28_4;
  wire [7:0] t_r21_c28_5;
  wire [7:0] t_r21_c28_6;
  wire [7:0] t_r21_c28_7;
  wire [7:0] t_r21_c28_8;
  wire [7:0] t_r21_c28_9;
  wire [7:0] t_r21_c28_10;
  wire [7:0] t_r21_c28_11;
  wire [7:0] t_r21_c28_12;
  wire [7:0] t_r21_c29_0;
  wire [7:0] t_r21_c29_1;
  wire [7:0] t_r21_c29_2;
  wire [7:0] t_r21_c29_3;
  wire [7:0] t_r21_c29_4;
  wire [7:0] t_r21_c29_5;
  wire [7:0] t_r21_c29_6;
  wire [7:0] t_r21_c29_7;
  wire [7:0] t_r21_c29_8;
  wire [7:0] t_r21_c29_9;
  wire [7:0] t_r21_c29_10;
  wire [7:0] t_r21_c29_11;
  wire [7:0] t_r21_c29_12;
  wire [7:0] t_r21_c30_0;
  wire [7:0] t_r21_c30_1;
  wire [7:0] t_r21_c30_2;
  wire [7:0] t_r21_c30_3;
  wire [7:0] t_r21_c30_4;
  wire [7:0] t_r21_c30_5;
  wire [7:0] t_r21_c30_6;
  wire [7:0] t_r21_c30_7;
  wire [7:0] t_r21_c30_8;
  wire [7:0] t_r21_c30_9;
  wire [7:0] t_r21_c30_10;
  wire [7:0] t_r21_c30_11;
  wire [7:0] t_r21_c30_12;
  wire [7:0] t_r21_c31_0;
  wire [7:0] t_r21_c31_1;
  wire [7:0] t_r21_c31_2;
  wire [7:0] t_r21_c31_3;
  wire [7:0] t_r21_c31_4;
  wire [7:0] t_r21_c31_5;
  wire [7:0] t_r21_c31_6;
  wire [7:0] t_r21_c31_7;
  wire [7:0] t_r21_c31_8;
  wire [7:0] t_r21_c31_9;
  wire [7:0] t_r21_c31_10;
  wire [7:0] t_r21_c31_11;
  wire [7:0] t_r21_c31_12;
  wire [7:0] t_r21_c32_0;
  wire [7:0] t_r21_c32_1;
  wire [7:0] t_r21_c32_2;
  wire [7:0] t_r21_c32_3;
  wire [7:0] t_r21_c32_4;
  wire [7:0] t_r21_c32_5;
  wire [7:0] t_r21_c32_6;
  wire [7:0] t_r21_c32_7;
  wire [7:0] t_r21_c32_8;
  wire [7:0] t_r21_c32_9;
  wire [7:0] t_r21_c32_10;
  wire [7:0] t_r21_c32_11;
  wire [7:0] t_r21_c32_12;
  wire [7:0] t_r21_c33_0;
  wire [7:0] t_r21_c33_1;
  wire [7:0] t_r21_c33_2;
  wire [7:0] t_r21_c33_3;
  wire [7:0] t_r21_c33_4;
  wire [7:0] t_r21_c33_5;
  wire [7:0] t_r21_c33_6;
  wire [7:0] t_r21_c33_7;
  wire [7:0] t_r21_c33_8;
  wire [7:0] t_r21_c33_9;
  wire [7:0] t_r21_c33_10;
  wire [7:0] t_r21_c33_11;
  wire [7:0] t_r21_c33_12;
  wire [7:0] t_r21_c34_0;
  wire [7:0] t_r21_c34_1;
  wire [7:0] t_r21_c34_2;
  wire [7:0] t_r21_c34_3;
  wire [7:0] t_r21_c34_4;
  wire [7:0] t_r21_c34_5;
  wire [7:0] t_r21_c34_6;
  wire [7:0] t_r21_c34_7;
  wire [7:0] t_r21_c34_8;
  wire [7:0] t_r21_c34_9;
  wire [7:0] t_r21_c34_10;
  wire [7:0] t_r21_c34_11;
  wire [7:0] t_r21_c34_12;
  wire [7:0] t_r21_c35_0;
  wire [7:0] t_r21_c35_1;
  wire [7:0] t_r21_c35_2;
  wire [7:0] t_r21_c35_3;
  wire [7:0] t_r21_c35_4;
  wire [7:0] t_r21_c35_5;
  wire [7:0] t_r21_c35_6;
  wire [7:0] t_r21_c35_7;
  wire [7:0] t_r21_c35_8;
  wire [7:0] t_r21_c35_9;
  wire [7:0] t_r21_c35_10;
  wire [7:0] t_r21_c35_11;
  wire [7:0] t_r21_c35_12;
  wire [7:0] t_r21_c36_0;
  wire [7:0] t_r21_c36_1;
  wire [7:0] t_r21_c36_2;
  wire [7:0] t_r21_c36_3;
  wire [7:0] t_r21_c36_4;
  wire [7:0] t_r21_c36_5;
  wire [7:0] t_r21_c36_6;
  wire [7:0] t_r21_c36_7;
  wire [7:0] t_r21_c36_8;
  wire [7:0] t_r21_c36_9;
  wire [7:0] t_r21_c36_10;
  wire [7:0] t_r21_c36_11;
  wire [7:0] t_r21_c36_12;
  wire [7:0] t_r21_c37_0;
  wire [7:0] t_r21_c37_1;
  wire [7:0] t_r21_c37_2;
  wire [7:0] t_r21_c37_3;
  wire [7:0] t_r21_c37_4;
  wire [7:0] t_r21_c37_5;
  wire [7:0] t_r21_c37_6;
  wire [7:0] t_r21_c37_7;
  wire [7:0] t_r21_c37_8;
  wire [7:0] t_r21_c37_9;
  wire [7:0] t_r21_c37_10;
  wire [7:0] t_r21_c37_11;
  wire [7:0] t_r21_c37_12;
  wire [7:0] t_r21_c38_0;
  wire [7:0] t_r21_c38_1;
  wire [7:0] t_r21_c38_2;
  wire [7:0] t_r21_c38_3;
  wire [7:0] t_r21_c38_4;
  wire [7:0] t_r21_c38_5;
  wire [7:0] t_r21_c38_6;
  wire [7:0] t_r21_c38_7;
  wire [7:0] t_r21_c38_8;
  wire [7:0] t_r21_c38_9;
  wire [7:0] t_r21_c38_10;
  wire [7:0] t_r21_c38_11;
  wire [7:0] t_r21_c38_12;
  wire [7:0] t_r21_c39_0;
  wire [7:0] t_r21_c39_1;
  wire [7:0] t_r21_c39_2;
  wire [7:0] t_r21_c39_3;
  wire [7:0] t_r21_c39_4;
  wire [7:0] t_r21_c39_5;
  wire [7:0] t_r21_c39_6;
  wire [7:0] t_r21_c39_7;
  wire [7:0] t_r21_c39_8;
  wire [7:0] t_r21_c39_9;
  wire [7:0] t_r21_c39_10;
  wire [7:0] t_r21_c39_11;
  wire [7:0] t_r21_c39_12;
  wire [7:0] t_r21_c40_0;
  wire [7:0] t_r21_c40_1;
  wire [7:0] t_r21_c40_2;
  wire [7:0] t_r21_c40_3;
  wire [7:0] t_r21_c40_4;
  wire [7:0] t_r21_c40_5;
  wire [7:0] t_r21_c40_6;
  wire [7:0] t_r21_c40_7;
  wire [7:0] t_r21_c40_8;
  wire [7:0] t_r21_c40_9;
  wire [7:0] t_r21_c40_10;
  wire [7:0] t_r21_c40_11;
  wire [7:0] t_r21_c40_12;
  wire [7:0] t_r21_c41_0;
  wire [7:0] t_r21_c41_1;
  wire [7:0] t_r21_c41_2;
  wire [7:0] t_r21_c41_3;
  wire [7:0] t_r21_c41_4;
  wire [7:0] t_r21_c41_5;
  wire [7:0] t_r21_c41_6;
  wire [7:0] t_r21_c41_7;
  wire [7:0] t_r21_c41_8;
  wire [7:0] t_r21_c41_9;
  wire [7:0] t_r21_c41_10;
  wire [7:0] t_r21_c41_11;
  wire [7:0] t_r21_c41_12;
  wire [7:0] t_r21_c42_0;
  wire [7:0] t_r21_c42_1;
  wire [7:0] t_r21_c42_2;
  wire [7:0] t_r21_c42_3;
  wire [7:0] t_r21_c42_4;
  wire [7:0] t_r21_c42_5;
  wire [7:0] t_r21_c42_6;
  wire [7:0] t_r21_c42_7;
  wire [7:0] t_r21_c42_8;
  wire [7:0] t_r21_c42_9;
  wire [7:0] t_r21_c42_10;
  wire [7:0] t_r21_c42_11;
  wire [7:0] t_r21_c42_12;
  wire [7:0] t_r21_c43_0;
  wire [7:0] t_r21_c43_1;
  wire [7:0] t_r21_c43_2;
  wire [7:0] t_r21_c43_3;
  wire [7:0] t_r21_c43_4;
  wire [7:0] t_r21_c43_5;
  wire [7:0] t_r21_c43_6;
  wire [7:0] t_r21_c43_7;
  wire [7:0] t_r21_c43_8;
  wire [7:0] t_r21_c43_9;
  wire [7:0] t_r21_c43_10;
  wire [7:0] t_r21_c43_11;
  wire [7:0] t_r21_c43_12;
  wire [7:0] t_r21_c44_0;
  wire [7:0] t_r21_c44_1;
  wire [7:0] t_r21_c44_2;
  wire [7:0] t_r21_c44_3;
  wire [7:0] t_r21_c44_4;
  wire [7:0] t_r21_c44_5;
  wire [7:0] t_r21_c44_6;
  wire [7:0] t_r21_c44_7;
  wire [7:0] t_r21_c44_8;
  wire [7:0] t_r21_c44_9;
  wire [7:0] t_r21_c44_10;
  wire [7:0] t_r21_c44_11;
  wire [7:0] t_r21_c44_12;
  wire [7:0] t_r21_c45_0;
  wire [7:0] t_r21_c45_1;
  wire [7:0] t_r21_c45_2;
  wire [7:0] t_r21_c45_3;
  wire [7:0] t_r21_c45_4;
  wire [7:0] t_r21_c45_5;
  wire [7:0] t_r21_c45_6;
  wire [7:0] t_r21_c45_7;
  wire [7:0] t_r21_c45_8;
  wire [7:0] t_r21_c45_9;
  wire [7:0] t_r21_c45_10;
  wire [7:0] t_r21_c45_11;
  wire [7:0] t_r21_c45_12;
  wire [7:0] t_r21_c46_0;
  wire [7:0] t_r21_c46_1;
  wire [7:0] t_r21_c46_2;
  wire [7:0] t_r21_c46_3;
  wire [7:0] t_r21_c46_4;
  wire [7:0] t_r21_c46_5;
  wire [7:0] t_r21_c46_6;
  wire [7:0] t_r21_c46_7;
  wire [7:0] t_r21_c46_8;
  wire [7:0] t_r21_c46_9;
  wire [7:0] t_r21_c46_10;
  wire [7:0] t_r21_c46_11;
  wire [7:0] t_r21_c46_12;
  wire [7:0] t_r21_c47_0;
  wire [7:0] t_r21_c47_1;
  wire [7:0] t_r21_c47_2;
  wire [7:0] t_r21_c47_3;
  wire [7:0] t_r21_c47_4;
  wire [7:0] t_r21_c47_5;
  wire [7:0] t_r21_c47_6;
  wire [7:0] t_r21_c47_7;
  wire [7:0] t_r21_c47_8;
  wire [7:0] t_r21_c47_9;
  wire [7:0] t_r21_c47_10;
  wire [7:0] t_r21_c47_11;
  wire [7:0] t_r21_c47_12;
  wire [7:0] t_r21_c48_0;
  wire [7:0] t_r21_c48_1;
  wire [7:0] t_r21_c48_2;
  wire [7:0] t_r21_c48_3;
  wire [7:0] t_r21_c48_4;
  wire [7:0] t_r21_c48_5;
  wire [7:0] t_r21_c48_6;
  wire [7:0] t_r21_c48_7;
  wire [7:0] t_r21_c48_8;
  wire [7:0] t_r21_c48_9;
  wire [7:0] t_r21_c48_10;
  wire [7:0] t_r21_c48_11;
  wire [7:0] t_r21_c48_12;
  wire [7:0] t_r21_c49_0;
  wire [7:0] t_r21_c49_1;
  wire [7:0] t_r21_c49_2;
  wire [7:0] t_r21_c49_3;
  wire [7:0] t_r21_c49_4;
  wire [7:0] t_r21_c49_5;
  wire [7:0] t_r21_c49_6;
  wire [7:0] t_r21_c49_7;
  wire [7:0] t_r21_c49_8;
  wire [7:0] t_r21_c49_9;
  wire [7:0] t_r21_c49_10;
  wire [7:0] t_r21_c49_11;
  wire [7:0] t_r21_c49_12;
  wire [7:0] t_r21_c50_0;
  wire [7:0] t_r21_c50_1;
  wire [7:0] t_r21_c50_2;
  wire [7:0] t_r21_c50_3;
  wire [7:0] t_r21_c50_4;
  wire [7:0] t_r21_c50_5;
  wire [7:0] t_r21_c50_6;
  wire [7:0] t_r21_c50_7;
  wire [7:0] t_r21_c50_8;
  wire [7:0] t_r21_c50_9;
  wire [7:0] t_r21_c50_10;
  wire [7:0] t_r21_c50_11;
  wire [7:0] t_r21_c50_12;
  wire [7:0] t_r21_c51_0;
  wire [7:0] t_r21_c51_1;
  wire [7:0] t_r21_c51_2;
  wire [7:0] t_r21_c51_3;
  wire [7:0] t_r21_c51_4;
  wire [7:0] t_r21_c51_5;
  wire [7:0] t_r21_c51_6;
  wire [7:0] t_r21_c51_7;
  wire [7:0] t_r21_c51_8;
  wire [7:0] t_r21_c51_9;
  wire [7:0] t_r21_c51_10;
  wire [7:0] t_r21_c51_11;
  wire [7:0] t_r21_c51_12;
  wire [7:0] t_r21_c52_0;
  wire [7:0] t_r21_c52_1;
  wire [7:0] t_r21_c52_2;
  wire [7:0] t_r21_c52_3;
  wire [7:0] t_r21_c52_4;
  wire [7:0] t_r21_c52_5;
  wire [7:0] t_r21_c52_6;
  wire [7:0] t_r21_c52_7;
  wire [7:0] t_r21_c52_8;
  wire [7:0] t_r21_c52_9;
  wire [7:0] t_r21_c52_10;
  wire [7:0] t_r21_c52_11;
  wire [7:0] t_r21_c52_12;
  wire [7:0] t_r21_c53_0;
  wire [7:0] t_r21_c53_1;
  wire [7:0] t_r21_c53_2;
  wire [7:0] t_r21_c53_3;
  wire [7:0] t_r21_c53_4;
  wire [7:0] t_r21_c53_5;
  wire [7:0] t_r21_c53_6;
  wire [7:0] t_r21_c53_7;
  wire [7:0] t_r21_c53_8;
  wire [7:0] t_r21_c53_9;
  wire [7:0] t_r21_c53_10;
  wire [7:0] t_r21_c53_11;
  wire [7:0] t_r21_c53_12;
  wire [7:0] t_r21_c54_0;
  wire [7:0] t_r21_c54_1;
  wire [7:0] t_r21_c54_2;
  wire [7:0] t_r21_c54_3;
  wire [7:0] t_r21_c54_4;
  wire [7:0] t_r21_c54_5;
  wire [7:0] t_r21_c54_6;
  wire [7:0] t_r21_c54_7;
  wire [7:0] t_r21_c54_8;
  wire [7:0] t_r21_c54_9;
  wire [7:0] t_r21_c54_10;
  wire [7:0] t_r21_c54_11;
  wire [7:0] t_r21_c54_12;
  wire [7:0] t_r21_c55_0;
  wire [7:0] t_r21_c55_1;
  wire [7:0] t_r21_c55_2;
  wire [7:0] t_r21_c55_3;
  wire [7:0] t_r21_c55_4;
  wire [7:0] t_r21_c55_5;
  wire [7:0] t_r21_c55_6;
  wire [7:0] t_r21_c55_7;
  wire [7:0] t_r21_c55_8;
  wire [7:0] t_r21_c55_9;
  wire [7:0] t_r21_c55_10;
  wire [7:0] t_r21_c55_11;
  wire [7:0] t_r21_c55_12;
  wire [7:0] t_r21_c56_0;
  wire [7:0] t_r21_c56_1;
  wire [7:0] t_r21_c56_2;
  wire [7:0] t_r21_c56_3;
  wire [7:0] t_r21_c56_4;
  wire [7:0] t_r21_c56_5;
  wire [7:0] t_r21_c56_6;
  wire [7:0] t_r21_c56_7;
  wire [7:0] t_r21_c56_8;
  wire [7:0] t_r21_c56_9;
  wire [7:0] t_r21_c56_10;
  wire [7:0] t_r21_c56_11;
  wire [7:0] t_r21_c56_12;
  wire [7:0] t_r21_c57_0;
  wire [7:0] t_r21_c57_1;
  wire [7:0] t_r21_c57_2;
  wire [7:0] t_r21_c57_3;
  wire [7:0] t_r21_c57_4;
  wire [7:0] t_r21_c57_5;
  wire [7:0] t_r21_c57_6;
  wire [7:0] t_r21_c57_7;
  wire [7:0] t_r21_c57_8;
  wire [7:0] t_r21_c57_9;
  wire [7:0] t_r21_c57_10;
  wire [7:0] t_r21_c57_11;
  wire [7:0] t_r21_c57_12;
  wire [7:0] t_r21_c58_0;
  wire [7:0] t_r21_c58_1;
  wire [7:0] t_r21_c58_2;
  wire [7:0] t_r21_c58_3;
  wire [7:0] t_r21_c58_4;
  wire [7:0] t_r21_c58_5;
  wire [7:0] t_r21_c58_6;
  wire [7:0] t_r21_c58_7;
  wire [7:0] t_r21_c58_8;
  wire [7:0] t_r21_c58_9;
  wire [7:0] t_r21_c58_10;
  wire [7:0] t_r21_c58_11;
  wire [7:0] t_r21_c58_12;
  wire [7:0] t_r21_c59_0;
  wire [7:0] t_r21_c59_1;
  wire [7:0] t_r21_c59_2;
  wire [7:0] t_r21_c59_3;
  wire [7:0] t_r21_c59_4;
  wire [7:0] t_r21_c59_5;
  wire [7:0] t_r21_c59_6;
  wire [7:0] t_r21_c59_7;
  wire [7:0] t_r21_c59_8;
  wire [7:0] t_r21_c59_9;
  wire [7:0] t_r21_c59_10;
  wire [7:0] t_r21_c59_11;
  wire [7:0] t_r21_c59_12;
  wire [7:0] t_r21_c60_0;
  wire [7:0] t_r21_c60_1;
  wire [7:0] t_r21_c60_2;
  wire [7:0] t_r21_c60_3;
  wire [7:0] t_r21_c60_4;
  wire [7:0] t_r21_c60_5;
  wire [7:0] t_r21_c60_6;
  wire [7:0] t_r21_c60_7;
  wire [7:0] t_r21_c60_8;
  wire [7:0] t_r21_c60_9;
  wire [7:0] t_r21_c60_10;
  wire [7:0] t_r21_c60_11;
  wire [7:0] t_r21_c60_12;
  wire [7:0] t_r21_c61_0;
  wire [7:0] t_r21_c61_1;
  wire [7:0] t_r21_c61_2;
  wire [7:0] t_r21_c61_3;
  wire [7:0] t_r21_c61_4;
  wire [7:0] t_r21_c61_5;
  wire [7:0] t_r21_c61_6;
  wire [7:0] t_r21_c61_7;
  wire [7:0] t_r21_c61_8;
  wire [7:0] t_r21_c61_9;
  wire [7:0] t_r21_c61_10;
  wire [7:0] t_r21_c61_11;
  wire [7:0] t_r21_c61_12;
  wire [7:0] t_r21_c62_0;
  wire [7:0] t_r21_c62_1;
  wire [7:0] t_r21_c62_2;
  wire [7:0] t_r21_c62_3;
  wire [7:0] t_r21_c62_4;
  wire [7:0] t_r21_c62_5;
  wire [7:0] t_r21_c62_6;
  wire [7:0] t_r21_c62_7;
  wire [7:0] t_r21_c62_8;
  wire [7:0] t_r21_c62_9;
  wire [7:0] t_r21_c62_10;
  wire [7:0] t_r21_c62_11;
  wire [7:0] t_r21_c62_12;
  wire [7:0] t_r21_c63_0;
  wire [7:0] t_r21_c63_1;
  wire [7:0] t_r21_c63_2;
  wire [7:0] t_r21_c63_3;
  wire [7:0] t_r21_c63_4;
  wire [7:0] t_r21_c63_5;
  wire [7:0] t_r21_c63_6;
  wire [7:0] t_r21_c63_7;
  wire [7:0] t_r21_c63_8;
  wire [7:0] t_r21_c63_9;
  wire [7:0] t_r21_c63_10;
  wire [7:0] t_r21_c63_11;
  wire [7:0] t_r21_c63_12;
  wire [7:0] t_r21_c64_0;
  wire [7:0] t_r21_c64_1;
  wire [7:0] t_r21_c64_2;
  wire [7:0] t_r21_c64_3;
  wire [7:0] t_r21_c64_4;
  wire [7:0] t_r21_c64_5;
  wire [7:0] t_r21_c64_6;
  wire [7:0] t_r21_c64_7;
  wire [7:0] t_r21_c64_8;
  wire [7:0] t_r21_c64_9;
  wire [7:0] t_r21_c64_10;
  wire [7:0] t_r21_c64_11;
  wire [7:0] t_r21_c64_12;
  wire [7:0] t_r21_c65_0;
  wire [7:0] t_r21_c65_1;
  wire [7:0] t_r21_c65_2;
  wire [7:0] t_r21_c65_3;
  wire [7:0] t_r21_c65_4;
  wire [7:0] t_r21_c65_5;
  wire [7:0] t_r21_c65_6;
  wire [7:0] t_r21_c65_7;
  wire [7:0] t_r21_c65_8;
  wire [7:0] t_r21_c65_9;
  wire [7:0] t_r21_c65_10;
  wire [7:0] t_r21_c65_11;
  wire [7:0] t_r21_c65_12;
  wire [7:0] t_r22_c0_0;
  wire [7:0] t_r22_c0_1;
  wire [7:0] t_r22_c0_2;
  wire [7:0] t_r22_c0_3;
  wire [7:0] t_r22_c0_4;
  wire [7:0] t_r22_c0_5;
  wire [7:0] t_r22_c0_6;
  wire [7:0] t_r22_c0_7;
  wire [7:0] t_r22_c0_8;
  wire [7:0] t_r22_c0_9;
  wire [7:0] t_r22_c0_10;
  wire [7:0] t_r22_c0_11;
  wire [7:0] t_r22_c0_12;
  wire [7:0] t_r22_c1_0;
  wire [7:0] t_r22_c1_1;
  wire [7:0] t_r22_c1_2;
  wire [7:0] t_r22_c1_3;
  wire [7:0] t_r22_c1_4;
  wire [7:0] t_r22_c1_5;
  wire [7:0] t_r22_c1_6;
  wire [7:0] t_r22_c1_7;
  wire [7:0] t_r22_c1_8;
  wire [7:0] t_r22_c1_9;
  wire [7:0] t_r22_c1_10;
  wire [7:0] t_r22_c1_11;
  wire [7:0] t_r22_c1_12;
  wire [7:0] t_r22_c2_0;
  wire [7:0] t_r22_c2_1;
  wire [7:0] t_r22_c2_2;
  wire [7:0] t_r22_c2_3;
  wire [7:0] t_r22_c2_4;
  wire [7:0] t_r22_c2_5;
  wire [7:0] t_r22_c2_6;
  wire [7:0] t_r22_c2_7;
  wire [7:0] t_r22_c2_8;
  wire [7:0] t_r22_c2_9;
  wire [7:0] t_r22_c2_10;
  wire [7:0] t_r22_c2_11;
  wire [7:0] t_r22_c2_12;
  wire [7:0] t_r22_c3_0;
  wire [7:0] t_r22_c3_1;
  wire [7:0] t_r22_c3_2;
  wire [7:0] t_r22_c3_3;
  wire [7:0] t_r22_c3_4;
  wire [7:0] t_r22_c3_5;
  wire [7:0] t_r22_c3_6;
  wire [7:0] t_r22_c3_7;
  wire [7:0] t_r22_c3_8;
  wire [7:0] t_r22_c3_9;
  wire [7:0] t_r22_c3_10;
  wire [7:0] t_r22_c3_11;
  wire [7:0] t_r22_c3_12;
  wire [7:0] t_r22_c4_0;
  wire [7:0] t_r22_c4_1;
  wire [7:0] t_r22_c4_2;
  wire [7:0] t_r22_c4_3;
  wire [7:0] t_r22_c4_4;
  wire [7:0] t_r22_c4_5;
  wire [7:0] t_r22_c4_6;
  wire [7:0] t_r22_c4_7;
  wire [7:0] t_r22_c4_8;
  wire [7:0] t_r22_c4_9;
  wire [7:0] t_r22_c4_10;
  wire [7:0] t_r22_c4_11;
  wire [7:0] t_r22_c4_12;
  wire [7:0] t_r22_c5_0;
  wire [7:0] t_r22_c5_1;
  wire [7:0] t_r22_c5_2;
  wire [7:0] t_r22_c5_3;
  wire [7:0] t_r22_c5_4;
  wire [7:0] t_r22_c5_5;
  wire [7:0] t_r22_c5_6;
  wire [7:0] t_r22_c5_7;
  wire [7:0] t_r22_c5_8;
  wire [7:0] t_r22_c5_9;
  wire [7:0] t_r22_c5_10;
  wire [7:0] t_r22_c5_11;
  wire [7:0] t_r22_c5_12;
  wire [7:0] t_r22_c6_0;
  wire [7:0] t_r22_c6_1;
  wire [7:0] t_r22_c6_2;
  wire [7:0] t_r22_c6_3;
  wire [7:0] t_r22_c6_4;
  wire [7:0] t_r22_c6_5;
  wire [7:0] t_r22_c6_6;
  wire [7:0] t_r22_c6_7;
  wire [7:0] t_r22_c6_8;
  wire [7:0] t_r22_c6_9;
  wire [7:0] t_r22_c6_10;
  wire [7:0] t_r22_c6_11;
  wire [7:0] t_r22_c6_12;
  wire [7:0] t_r22_c7_0;
  wire [7:0] t_r22_c7_1;
  wire [7:0] t_r22_c7_2;
  wire [7:0] t_r22_c7_3;
  wire [7:0] t_r22_c7_4;
  wire [7:0] t_r22_c7_5;
  wire [7:0] t_r22_c7_6;
  wire [7:0] t_r22_c7_7;
  wire [7:0] t_r22_c7_8;
  wire [7:0] t_r22_c7_9;
  wire [7:0] t_r22_c7_10;
  wire [7:0] t_r22_c7_11;
  wire [7:0] t_r22_c7_12;
  wire [7:0] t_r22_c8_0;
  wire [7:0] t_r22_c8_1;
  wire [7:0] t_r22_c8_2;
  wire [7:0] t_r22_c8_3;
  wire [7:0] t_r22_c8_4;
  wire [7:0] t_r22_c8_5;
  wire [7:0] t_r22_c8_6;
  wire [7:0] t_r22_c8_7;
  wire [7:0] t_r22_c8_8;
  wire [7:0] t_r22_c8_9;
  wire [7:0] t_r22_c8_10;
  wire [7:0] t_r22_c8_11;
  wire [7:0] t_r22_c8_12;
  wire [7:0] t_r22_c9_0;
  wire [7:0] t_r22_c9_1;
  wire [7:0] t_r22_c9_2;
  wire [7:0] t_r22_c9_3;
  wire [7:0] t_r22_c9_4;
  wire [7:0] t_r22_c9_5;
  wire [7:0] t_r22_c9_6;
  wire [7:0] t_r22_c9_7;
  wire [7:0] t_r22_c9_8;
  wire [7:0] t_r22_c9_9;
  wire [7:0] t_r22_c9_10;
  wire [7:0] t_r22_c9_11;
  wire [7:0] t_r22_c9_12;
  wire [7:0] t_r22_c10_0;
  wire [7:0] t_r22_c10_1;
  wire [7:0] t_r22_c10_2;
  wire [7:0] t_r22_c10_3;
  wire [7:0] t_r22_c10_4;
  wire [7:0] t_r22_c10_5;
  wire [7:0] t_r22_c10_6;
  wire [7:0] t_r22_c10_7;
  wire [7:0] t_r22_c10_8;
  wire [7:0] t_r22_c10_9;
  wire [7:0] t_r22_c10_10;
  wire [7:0] t_r22_c10_11;
  wire [7:0] t_r22_c10_12;
  wire [7:0] t_r22_c11_0;
  wire [7:0] t_r22_c11_1;
  wire [7:0] t_r22_c11_2;
  wire [7:0] t_r22_c11_3;
  wire [7:0] t_r22_c11_4;
  wire [7:0] t_r22_c11_5;
  wire [7:0] t_r22_c11_6;
  wire [7:0] t_r22_c11_7;
  wire [7:0] t_r22_c11_8;
  wire [7:0] t_r22_c11_9;
  wire [7:0] t_r22_c11_10;
  wire [7:0] t_r22_c11_11;
  wire [7:0] t_r22_c11_12;
  wire [7:0] t_r22_c12_0;
  wire [7:0] t_r22_c12_1;
  wire [7:0] t_r22_c12_2;
  wire [7:0] t_r22_c12_3;
  wire [7:0] t_r22_c12_4;
  wire [7:0] t_r22_c12_5;
  wire [7:0] t_r22_c12_6;
  wire [7:0] t_r22_c12_7;
  wire [7:0] t_r22_c12_8;
  wire [7:0] t_r22_c12_9;
  wire [7:0] t_r22_c12_10;
  wire [7:0] t_r22_c12_11;
  wire [7:0] t_r22_c12_12;
  wire [7:0] t_r22_c13_0;
  wire [7:0] t_r22_c13_1;
  wire [7:0] t_r22_c13_2;
  wire [7:0] t_r22_c13_3;
  wire [7:0] t_r22_c13_4;
  wire [7:0] t_r22_c13_5;
  wire [7:0] t_r22_c13_6;
  wire [7:0] t_r22_c13_7;
  wire [7:0] t_r22_c13_8;
  wire [7:0] t_r22_c13_9;
  wire [7:0] t_r22_c13_10;
  wire [7:0] t_r22_c13_11;
  wire [7:0] t_r22_c13_12;
  wire [7:0] t_r22_c14_0;
  wire [7:0] t_r22_c14_1;
  wire [7:0] t_r22_c14_2;
  wire [7:0] t_r22_c14_3;
  wire [7:0] t_r22_c14_4;
  wire [7:0] t_r22_c14_5;
  wire [7:0] t_r22_c14_6;
  wire [7:0] t_r22_c14_7;
  wire [7:0] t_r22_c14_8;
  wire [7:0] t_r22_c14_9;
  wire [7:0] t_r22_c14_10;
  wire [7:0] t_r22_c14_11;
  wire [7:0] t_r22_c14_12;
  wire [7:0] t_r22_c15_0;
  wire [7:0] t_r22_c15_1;
  wire [7:0] t_r22_c15_2;
  wire [7:0] t_r22_c15_3;
  wire [7:0] t_r22_c15_4;
  wire [7:0] t_r22_c15_5;
  wire [7:0] t_r22_c15_6;
  wire [7:0] t_r22_c15_7;
  wire [7:0] t_r22_c15_8;
  wire [7:0] t_r22_c15_9;
  wire [7:0] t_r22_c15_10;
  wire [7:0] t_r22_c15_11;
  wire [7:0] t_r22_c15_12;
  wire [7:0] t_r22_c16_0;
  wire [7:0] t_r22_c16_1;
  wire [7:0] t_r22_c16_2;
  wire [7:0] t_r22_c16_3;
  wire [7:0] t_r22_c16_4;
  wire [7:0] t_r22_c16_5;
  wire [7:0] t_r22_c16_6;
  wire [7:0] t_r22_c16_7;
  wire [7:0] t_r22_c16_8;
  wire [7:0] t_r22_c16_9;
  wire [7:0] t_r22_c16_10;
  wire [7:0] t_r22_c16_11;
  wire [7:0] t_r22_c16_12;
  wire [7:0] t_r22_c17_0;
  wire [7:0] t_r22_c17_1;
  wire [7:0] t_r22_c17_2;
  wire [7:0] t_r22_c17_3;
  wire [7:0] t_r22_c17_4;
  wire [7:0] t_r22_c17_5;
  wire [7:0] t_r22_c17_6;
  wire [7:0] t_r22_c17_7;
  wire [7:0] t_r22_c17_8;
  wire [7:0] t_r22_c17_9;
  wire [7:0] t_r22_c17_10;
  wire [7:0] t_r22_c17_11;
  wire [7:0] t_r22_c17_12;
  wire [7:0] t_r22_c18_0;
  wire [7:0] t_r22_c18_1;
  wire [7:0] t_r22_c18_2;
  wire [7:0] t_r22_c18_3;
  wire [7:0] t_r22_c18_4;
  wire [7:0] t_r22_c18_5;
  wire [7:0] t_r22_c18_6;
  wire [7:0] t_r22_c18_7;
  wire [7:0] t_r22_c18_8;
  wire [7:0] t_r22_c18_9;
  wire [7:0] t_r22_c18_10;
  wire [7:0] t_r22_c18_11;
  wire [7:0] t_r22_c18_12;
  wire [7:0] t_r22_c19_0;
  wire [7:0] t_r22_c19_1;
  wire [7:0] t_r22_c19_2;
  wire [7:0] t_r22_c19_3;
  wire [7:0] t_r22_c19_4;
  wire [7:0] t_r22_c19_5;
  wire [7:0] t_r22_c19_6;
  wire [7:0] t_r22_c19_7;
  wire [7:0] t_r22_c19_8;
  wire [7:0] t_r22_c19_9;
  wire [7:0] t_r22_c19_10;
  wire [7:0] t_r22_c19_11;
  wire [7:0] t_r22_c19_12;
  wire [7:0] t_r22_c20_0;
  wire [7:0] t_r22_c20_1;
  wire [7:0] t_r22_c20_2;
  wire [7:0] t_r22_c20_3;
  wire [7:0] t_r22_c20_4;
  wire [7:0] t_r22_c20_5;
  wire [7:0] t_r22_c20_6;
  wire [7:0] t_r22_c20_7;
  wire [7:0] t_r22_c20_8;
  wire [7:0] t_r22_c20_9;
  wire [7:0] t_r22_c20_10;
  wire [7:0] t_r22_c20_11;
  wire [7:0] t_r22_c20_12;
  wire [7:0] t_r22_c21_0;
  wire [7:0] t_r22_c21_1;
  wire [7:0] t_r22_c21_2;
  wire [7:0] t_r22_c21_3;
  wire [7:0] t_r22_c21_4;
  wire [7:0] t_r22_c21_5;
  wire [7:0] t_r22_c21_6;
  wire [7:0] t_r22_c21_7;
  wire [7:0] t_r22_c21_8;
  wire [7:0] t_r22_c21_9;
  wire [7:0] t_r22_c21_10;
  wire [7:0] t_r22_c21_11;
  wire [7:0] t_r22_c21_12;
  wire [7:0] t_r22_c22_0;
  wire [7:0] t_r22_c22_1;
  wire [7:0] t_r22_c22_2;
  wire [7:0] t_r22_c22_3;
  wire [7:0] t_r22_c22_4;
  wire [7:0] t_r22_c22_5;
  wire [7:0] t_r22_c22_6;
  wire [7:0] t_r22_c22_7;
  wire [7:0] t_r22_c22_8;
  wire [7:0] t_r22_c22_9;
  wire [7:0] t_r22_c22_10;
  wire [7:0] t_r22_c22_11;
  wire [7:0] t_r22_c22_12;
  wire [7:0] t_r22_c23_0;
  wire [7:0] t_r22_c23_1;
  wire [7:0] t_r22_c23_2;
  wire [7:0] t_r22_c23_3;
  wire [7:0] t_r22_c23_4;
  wire [7:0] t_r22_c23_5;
  wire [7:0] t_r22_c23_6;
  wire [7:0] t_r22_c23_7;
  wire [7:0] t_r22_c23_8;
  wire [7:0] t_r22_c23_9;
  wire [7:0] t_r22_c23_10;
  wire [7:0] t_r22_c23_11;
  wire [7:0] t_r22_c23_12;
  wire [7:0] t_r22_c24_0;
  wire [7:0] t_r22_c24_1;
  wire [7:0] t_r22_c24_2;
  wire [7:0] t_r22_c24_3;
  wire [7:0] t_r22_c24_4;
  wire [7:0] t_r22_c24_5;
  wire [7:0] t_r22_c24_6;
  wire [7:0] t_r22_c24_7;
  wire [7:0] t_r22_c24_8;
  wire [7:0] t_r22_c24_9;
  wire [7:0] t_r22_c24_10;
  wire [7:0] t_r22_c24_11;
  wire [7:0] t_r22_c24_12;
  wire [7:0] t_r22_c25_0;
  wire [7:0] t_r22_c25_1;
  wire [7:0] t_r22_c25_2;
  wire [7:0] t_r22_c25_3;
  wire [7:0] t_r22_c25_4;
  wire [7:0] t_r22_c25_5;
  wire [7:0] t_r22_c25_6;
  wire [7:0] t_r22_c25_7;
  wire [7:0] t_r22_c25_8;
  wire [7:0] t_r22_c25_9;
  wire [7:0] t_r22_c25_10;
  wire [7:0] t_r22_c25_11;
  wire [7:0] t_r22_c25_12;
  wire [7:0] t_r22_c26_0;
  wire [7:0] t_r22_c26_1;
  wire [7:0] t_r22_c26_2;
  wire [7:0] t_r22_c26_3;
  wire [7:0] t_r22_c26_4;
  wire [7:0] t_r22_c26_5;
  wire [7:0] t_r22_c26_6;
  wire [7:0] t_r22_c26_7;
  wire [7:0] t_r22_c26_8;
  wire [7:0] t_r22_c26_9;
  wire [7:0] t_r22_c26_10;
  wire [7:0] t_r22_c26_11;
  wire [7:0] t_r22_c26_12;
  wire [7:0] t_r22_c27_0;
  wire [7:0] t_r22_c27_1;
  wire [7:0] t_r22_c27_2;
  wire [7:0] t_r22_c27_3;
  wire [7:0] t_r22_c27_4;
  wire [7:0] t_r22_c27_5;
  wire [7:0] t_r22_c27_6;
  wire [7:0] t_r22_c27_7;
  wire [7:0] t_r22_c27_8;
  wire [7:0] t_r22_c27_9;
  wire [7:0] t_r22_c27_10;
  wire [7:0] t_r22_c27_11;
  wire [7:0] t_r22_c27_12;
  wire [7:0] t_r22_c28_0;
  wire [7:0] t_r22_c28_1;
  wire [7:0] t_r22_c28_2;
  wire [7:0] t_r22_c28_3;
  wire [7:0] t_r22_c28_4;
  wire [7:0] t_r22_c28_5;
  wire [7:0] t_r22_c28_6;
  wire [7:0] t_r22_c28_7;
  wire [7:0] t_r22_c28_8;
  wire [7:0] t_r22_c28_9;
  wire [7:0] t_r22_c28_10;
  wire [7:0] t_r22_c28_11;
  wire [7:0] t_r22_c28_12;
  wire [7:0] t_r22_c29_0;
  wire [7:0] t_r22_c29_1;
  wire [7:0] t_r22_c29_2;
  wire [7:0] t_r22_c29_3;
  wire [7:0] t_r22_c29_4;
  wire [7:0] t_r22_c29_5;
  wire [7:0] t_r22_c29_6;
  wire [7:0] t_r22_c29_7;
  wire [7:0] t_r22_c29_8;
  wire [7:0] t_r22_c29_9;
  wire [7:0] t_r22_c29_10;
  wire [7:0] t_r22_c29_11;
  wire [7:0] t_r22_c29_12;
  wire [7:0] t_r22_c30_0;
  wire [7:0] t_r22_c30_1;
  wire [7:0] t_r22_c30_2;
  wire [7:0] t_r22_c30_3;
  wire [7:0] t_r22_c30_4;
  wire [7:0] t_r22_c30_5;
  wire [7:0] t_r22_c30_6;
  wire [7:0] t_r22_c30_7;
  wire [7:0] t_r22_c30_8;
  wire [7:0] t_r22_c30_9;
  wire [7:0] t_r22_c30_10;
  wire [7:0] t_r22_c30_11;
  wire [7:0] t_r22_c30_12;
  wire [7:0] t_r22_c31_0;
  wire [7:0] t_r22_c31_1;
  wire [7:0] t_r22_c31_2;
  wire [7:0] t_r22_c31_3;
  wire [7:0] t_r22_c31_4;
  wire [7:0] t_r22_c31_5;
  wire [7:0] t_r22_c31_6;
  wire [7:0] t_r22_c31_7;
  wire [7:0] t_r22_c31_8;
  wire [7:0] t_r22_c31_9;
  wire [7:0] t_r22_c31_10;
  wire [7:0] t_r22_c31_11;
  wire [7:0] t_r22_c31_12;
  wire [7:0] t_r22_c32_0;
  wire [7:0] t_r22_c32_1;
  wire [7:0] t_r22_c32_2;
  wire [7:0] t_r22_c32_3;
  wire [7:0] t_r22_c32_4;
  wire [7:0] t_r22_c32_5;
  wire [7:0] t_r22_c32_6;
  wire [7:0] t_r22_c32_7;
  wire [7:0] t_r22_c32_8;
  wire [7:0] t_r22_c32_9;
  wire [7:0] t_r22_c32_10;
  wire [7:0] t_r22_c32_11;
  wire [7:0] t_r22_c32_12;
  wire [7:0] t_r22_c33_0;
  wire [7:0] t_r22_c33_1;
  wire [7:0] t_r22_c33_2;
  wire [7:0] t_r22_c33_3;
  wire [7:0] t_r22_c33_4;
  wire [7:0] t_r22_c33_5;
  wire [7:0] t_r22_c33_6;
  wire [7:0] t_r22_c33_7;
  wire [7:0] t_r22_c33_8;
  wire [7:0] t_r22_c33_9;
  wire [7:0] t_r22_c33_10;
  wire [7:0] t_r22_c33_11;
  wire [7:0] t_r22_c33_12;
  wire [7:0] t_r22_c34_0;
  wire [7:0] t_r22_c34_1;
  wire [7:0] t_r22_c34_2;
  wire [7:0] t_r22_c34_3;
  wire [7:0] t_r22_c34_4;
  wire [7:0] t_r22_c34_5;
  wire [7:0] t_r22_c34_6;
  wire [7:0] t_r22_c34_7;
  wire [7:0] t_r22_c34_8;
  wire [7:0] t_r22_c34_9;
  wire [7:0] t_r22_c34_10;
  wire [7:0] t_r22_c34_11;
  wire [7:0] t_r22_c34_12;
  wire [7:0] t_r22_c35_0;
  wire [7:0] t_r22_c35_1;
  wire [7:0] t_r22_c35_2;
  wire [7:0] t_r22_c35_3;
  wire [7:0] t_r22_c35_4;
  wire [7:0] t_r22_c35_5;
  wire [7:0] t_r22_c35_6;
  wire [7:0] t_r22_c35_7;
  wire [7:0] t_r22_c35_8;
  wire [7:0] t_r22_c35_9;
  wire [7:0] t_r22_c35_10;
  wire [7:0] t_r22_c35_11;
  wire [7:0] t_r22_c35_12;
  wire [7:0] t_r22_c36_0;
  wire [7:0] t_r22_c36_1;
  wire [7:0] t_r22_c36_2;
  wire [7:0] t_r22_c36_3;
  wire [7:0] t_r22_c36_4;
  wire [7:0] t_r22_c36_5;
  wire [7:0] t_r22_c36_6;
  wire [7:0] t_r22_c36_7;
  wire [7:0] t_r22_c36_8;
  wire [7:0] t_r22_c36_9;
  wire [7:0] t_r22_c36_10;
  wire [7:0] t_r22_c36_11;
  wire [7:0] t_r22_c36_12;
  wire [7:0] t_r22_c37_0;
  wire [7:0] t_r22_c37_1;
  wire [7:0] t_r22_c37_2;
  wire [7:0] t_r22_c37_3;
  wire [7:0] t_r22_c37_4;
  wire [7:0] t_r22_c37_5;
  wire [7:0] t_r22_c37_6;
  wire [7:0] t_r22_c37_7;
  wire [7:0] t_r22_c37_8;
  wire [7:0] t_r22_c37_9;
  wire [7:0] t_r22_c37_10;
  wire [7:0] t_r22_c37_11;
  wire [7:0] t_r22_c37_12;
  wire [7:0] t_r22_c38_0;
  wire [7:0] t_r22_c38_1;
  wire [7:0] t_r22_c38_2;
  wire [7:0] t_r22_c38_3;
  wire [7:0] t_r22_c38_4;
  wire [7:0] t_r22_c38_5;
  wire [7:0] t_r22_c38_6;
  wire [7:0] t_r22_c38_7;
  wire [7:0] t_r22_c38_8;
  wire [7:0] t_r22_c38_9;
  wire [7:0] t_r22_c38_10;
  wire [7:0] t_r22_c38_11;
  wire [7:0] t_r22_c38_12;
  wire [7:0] t_r22_c39_0;
  wire [7:0] t_r22_c39_1;
  wire [7:0] t_r22_c39_2;
  wire [7:0] t_r22_c39_3;
  wire [7:0] t_r22_c39_4;
  wire [7:0] t_r22_c39_5;
  wire [7:0] t_r22_c39_6;
  wire [7:0] t_r22_c39_7;
  wire [7:0] t_r22_c39_8;
  wire [7:0] t_r22_c39_9;
  wire [7:0] t_r22_c39_10;
  wire [7:0] t_r22_c39_11;
  wire [7:0] t_r22_c39_12;
  wire [7:0] t_r22_c40_0;
  wire [7:0] t_r22_c40_1;
  wire [7:0] t_r22_c40_2;
  wire [7:0] t_r22_c40_3;
  wire [7:0] t_r22_c40_4;
  wire [7:0] t_r22_c40_5;
  wire [7:0] t_r22_c40_6;
  wire [7:0] t_r22_c40_7;
  wire [7:0] t_r22_c40_8;
  wire [7:0] t_r22_c40_9;
  wire [7:0] t_r22_c40_10;
  wire [7:0] t_r22_c40_11;
  wire [7:0] t_r22_c40_12;
  wire [7:0] t_r22_c41_0;
  wire [7:0] t_r22_c41_1;
  wire [7:0] t_r22_c41_2;
  wire [7:0] t_r22_c41_3;
  wire [7:0] t_r22_c41_4;
  wire [7:0] t_r22_c41_5;
  wire [7:0] t_r22_c41_6;
  wire [7:0] t_r22_c41_7;
  wire [7:0] t_r22_c41_8;
  wire [7:0] t_r22_c41_9;
  wire [7:0] t_r22_c41_10;
  wire [7:0] t_r22_c41_11;
  wire [7:0] t_r22_c41_12;
  wire [7:0] t_r22_c42_0;
  wire [7:0] t_r22_c42_1;
  wire [7:0] t_r22_c42_2;
  wire [7:0] t_r22_c42_3;
  wire [7:0] t_r22_c42_4;
  wire [7:0] t_r22_c42_5;
  wire [7:0] t_r22_c42_6;
  wire [7:0] t_r22_c42_7;
  wire [7:0] t_r22_c42_8;
  wire [7:0] t_r22_c42_9;
  wire [7:0] t_r22_c42_10;
  wire [7:0] t_r22_c42_11;
  wire [7:0] t_r22_c42_12;
  wire [7:0] t_r22_c43_0;
  wire [7:0] t_r22_c43_1;
  wire [7:0] t_r22_c43_2;
  wire [7:0] t_r22_c43_3;
  wire [7:0] t_r22_c43_4;
  wire [7:0] t_r22_c43_5;
  wire [7:0] t_r22_c43_6;
  wire [7:0] t_r22_c43_7;
  wire [7:0] t_r22_c43_8;
  wire [7:0] t_r22_c43_9;
  wire [7:0] t_r22_c43_10;
  wire [7:0] t_r22_c43_11;
  wire [7:0] t_r22_c43_12;
  wire [7:0] t_r22_c44_0;
  wire [7:0] t_r22_c44_1;
  wire [7:0] t_r22_c44_2;
  wire [7:0] t_r22_c44_3;
  wire [7:0] t_r22_c44_4;
  wire [7:0] t_r22_c44_5;
  wire [7:0] t_r22_c44_6;
  wire [7:0] t_r22_c44_7;
  wire [7:0] t_r22_c44_8;
  wire [7:0] t_r22_c44_9;
  wire [7:0] t_r22_c44_10;
  wire [7:0] t_r22_c44_11;
  wire [7:0] t_r22_c44_12;
  wire [7:0] t_r22_c45_0;
  wire [7:0] t_r22_c45_1;
  wire [7:0] t_r22_c45_2;
  wire [7:0] t_r22_c45_3;
  wire [7:0] t_r22_c45_4;
  wire [7:0] t_r22_c45_5;
  wire [7:0] t_r22_c45_6;
  wire [7:0] t_r22_c45_7;
  wire [7:0] t_r22_c45_8;
  wire [7:0] t_r22_c45_9;
  wire [7:0] t_r22_c45_10;
  wire [7:0] t_r22_c45_11;
  wire [7:0] t_r22_c45_12;
  wire [7:0] t_r22_c46_0;
  wire [7:0] t_r22_c46_1;
  wire [7:0] t_r22_c46_2;
  wire [7:0] t_r22_c46_3;
  wire [7:0] t_r22_c46_4;
  wire [7:0] t_r22_c46_5;
  wire [7:0] t_r22_c46_6;
  wire [7:0] t_r22_c46_7;
  wire [7:0] t_r22_c46_8;
  wire [7:0] t_r22_c46_9;
  wire [7:0] t_r22_c46_10;
  wire [7:0] t_r22_c46_11;
  wire [7:0] t_r22_c46_12;
  wire [7:0] t_r22_c47_0;
  wire [7:0] t_r22_c47_1;
  wire [7:0] t_r22_c47_2;
  wire [7:0] t_r22_c47_3;
  wire [7:0] t_r22_c47_4;
  wire [7:0] t_r22_c47_5;
  wire [7:0] t_r22_c47_6;
  wire [7:0] t_r22_c47_7;
  wire [7:0] t_r22_c47_8;
  wire [7:0] t_r22_c47_9;
  wire [7:0] t_r22_c47_10;
  wire [7:0] t_r22_c47_11;
  wire [7:0] t_r22_c47_12;
  wire [7:0] t_r22_c48_0;
  wire [7:0] t_r22_c48_1;
  wire [7:0] t_r22_c48_2;
  wire [7:0] t_r22_c48_3;
  wire [7:0] t_r22_c48_4;
  wire [7:0] t_r22_c48_5;
  wire [7:0] t_r22_c48_6;
  wire [7:0] t_r22_c48_7;
  wire [7:0] t_r22_c48_8;
  wire [7:0] t_r22_c48_9;
  wire [7:0] t_r22_c48_10;
  wire [7:0] t_r22_c48_11;
  wire [7:0] t_r22_c48_12;
  wire [7:0] t_r22_c49_0;
  wire [7:0] t_r22_c49_1;
  wire [7:0] t_r22_c49_2;
  wire [7:0] t_r22_c49_3;
  wire [7:0] t_r22_c49_4;
  wire [7:0] t_r22_c49_5;
  wire [7:0] t_r22_c49_6;
  wire [7:0] t_r22_c49_7;
  wire [7:0] t_r22_c49_8;
  wire [7:0] t_r22_c49_9;
  wire [7:0] t_r22_c49_10;
  wire [7:0] t_r22_c49_11;
  wire [7:0] t_r22_c49_12;
  wire [7:0] t_r22_c50_0;
  wire [7:0] t_r22_c50_1;
  wire [7:0] t_r22_c50_2;
  wire [7:0] t_r22_c50_3;
  wire [7:0] t_r22_c50_4;
  wire [7:0] t_r22_c50_5;
  wire [7:0] t_r22_c50_6;
  wire [7:0] t_r22_c50_7;
  wire [7:0] t_r22_c50_8;
  wire [7:0] t_r22_c50_9;
  wire [7:0] t_r22_c50_10;
  wire [7:0] t_r22_c50_11;
  wire [7:0] t_r22_c50_12;
  wire [7:0] t_r22_c51_0;
  wire [7:0] t_r22_c51_1;
  wire [7:0] t_r22_c51_2;
  wire [7:0] t_r22_c51_3;
  wire [7:0] t_r22_c51_4;
  wire [7:0] t_r22_c51_5;
  wire [7:0] t_r22_c51_6;
  wire [7:0] t_r22_c51_7;
  wire [7:0] t_r22_c51_8;
  wire [7:0] t_r22_c51_9;
  wire [7:0] t_r22_c51_10;
  wire [7:0] t_r22_c51_11;
  wire [7:0] t_r22_c51_12;
  wire [7:0] t_r22_c52_0;
  wire [7:0] t_r22_c52_1;
  wire [7:0] t_r22_c52_2;
  wire [7:0] t_r22_c52_3;
  wire [7:0] t_r22_c52_4;
  wire [7:0] t_r22_c52_5;
  wire [7:0] t_r22_c52_6;
  wire [7:0] t_r22_c52_7;
  wire [7:0] t_r22_c52_8;
  wire [7:0] t_r22_c52_9;
  wire [7:0] t_r22_c52_10;
  wire [7:0] t_r22_c52_11;
  wire [7:0] t_r22_c52_12;
  wire [7:0] t_r22_c53_0;
  wire [7:0] t_r22_c53_1;
  wire [7:0] t_r22_c53_2;
  wire [7:0] t_r22_c53_3;
  wire [7:0] t_r22_c53_4;
  wire [7:0] t_r22_c53_5;
  wire [7:0] t_r22_c53_6;
  wire [7:0] t_r22_c53_7;
  wire [7:0] t_r22_c53_8;
  wire [7:0] t_r22_c53_9;
  wire [7:0] t_r22_c53_10;
  wire [7:0] t_r22_c53_11;
  wire [7:0] t_r22_c53_12;
  wire [7:0] t_r22_c54_0;
  wire [7:0] t_r22_c54_1;
  wire [7:0] t_r22_c54_2;
  wire [7:0] t_r22_c54_3;
  wire [7:0] t_r22_c54_4;
  wire [7:0] t_r22_c54_5;
  wire [7:0] t_r22_c54_6;
  wire [7:0] t_r22_c54_7;
  wire [7:0] t_r22_c54_8;
  wire [7:0] t_r22_c54_9;
  wire [7:0] t_r22_c54_10;
  wire [7:0] t_r22_c54_11;
  wire [7:0] t_r22_c54_12;
  wire [7:0] t_r22_c55_0;
  wire [7:0] t_r22_c55_1;
  wire [7:0] t_r22_c55_2;
  wire [7:0] t_r22_c55_3;
  wire [7:0] t_r22_c55_4;
  wire [7:0] t_r22_c55_5;
  wire [7:0] t_r22_c55_6;
  wire [7:0] t_r22_c55_7;
  wire [7:0] t_r22_c55_8;
  wire [7:0] t_r22_c55_9;
  wire [7:0] t_r22_c55_10;
  wire [7:0] t_r22_c55_11;
  wire [7:0] t_r22_c55_12;
  wire [7:0] t_r22_c56_0;
  wire [7:0] t_r22_c56_1;
  wire [7:0] t_r22_c56_2;
  wire [7:0] t_r22_c56_3;
  wire [7:0] t_r22_c56_4;
  wire [7:0] t_r22_c56_5;
  wire [7:0] t_r22_c56_6;
  wire [7:0] t_r22_c56_7;
  wire [7:0] t_r22_c56_8;
  wire [7:0] t_r22_c56_9;
  wire [7:0] t_r22_c56_10;
  wire [7:0] t_r22_c56_11;
  wire [7:0] t_r22_c56_12;
  wire [7:0] t_r22_c57_0;
  wire [7:0] t_r22_c57_1;
  wire [7:0] t_r22_c57_2;
  wire [7:0] t_r22_c57_3;
  wire [7:0] t_r22_c57_4;
  wire [7:0] t_r22_c57_5;
  wire [7:0] t_r22_c57_6;
  wire [7:0] t_r22_c57_7;
  wire [7:0] t_r22_c57_8;
  wire [7:0] t_r22_c57_9;
  wire [7:0] t_r22_c57_10;
  wire [7:0] t_r22_c57_11;
  wire [7:0] t_r22_c57_12;
  wire [7:0] t_r22_c58_0;
  wire [7:0] t_r22_c58_1;
  wire [7:0] t_r22_c58_2;
  wire [7:0] t_r22_c58_3;
  wire [7:0] t_r22_c58_4;
  wire [7:0] t_r22_c58_5;
  wire [7:0] t_r22_c58_6;
  wire [7:0] t_r22_c58_7;
  wire [7:0] t_r22_c58_8;
  wire [7:0] t_r22_c58_9;
  wire [7:0] t_r22_c58_10;
  wire [7:0] t_r22_c58_11;
  wire [7:0] t_r22_c58_12;
  wire [7:0] t_r22_c59_0;
  wire [7:0] t_r22_c59_1;
  wire [7:0] t_r22_c59_2;
  wire [7:0] t_r22_c59_3;
  wire [7:0] t_r22_c59_4;
  wire [7:0] t_r22_c59_5;
  wire [7:0] t_r22_c59_6;
  wire [7:0] t_r22_c59_7;
  wire [7:0] t_r22_c59_8;
  wire [7:0] t_r22_c59_9;
  wire [7:0] t_r22_c59_10;
  wire [7:0] t_r22_c59_11;
  wire [7:0] t_r22_c59_12;
  wire [7:0] t_r22_c60_0;
  wire [7:0] t_r22_c60_1;
  wire [7:0] t_r22_c60_2;
  wire [7:0] t_r22_c60_3;
  wire [7:0] t_r22_c60_4;
  wire [7:0] t_r22_c60_5;
  wire [7:0] t_r22_c60_6;
  wire [7:0] t_r22_c60_7;
  wire [7:0] t_r22_c60_8;
  wire [7:0] t_r22_c60_9;
  wire [7:0] t_r22_c60_10;
  wire [7:0] t_r22_c60_11;
  wire [7:0] t_r22_c60_12;
  wire [7:0] t_r22_c61_0;
  wire [7:0] t_r22_c61_1;
  wire [7:0] t_r22_c61_2;
  wire [7:0] t_r22_c61_3;
  wire [7:0] t_r22_c61_4;
  wire [7:0] t_r22_c61_5;
  wire [7:0] t_r22_c61_6;
  wire [7:0] t_r22_c61_7;
  wire [7:0] t_r22_c61_8;
  wire [7:0] t_r22_c61_9;
  wire [7:0] t_r22_c61_10;
  wire [7:0] t_r22_c61_11;
  wire [7:0] t_r22_c61_12;
  wire [7:0] t_r22_c62_0;
  wire [7:0] t_r22_c62_1;
  wire [7:0] t_r22_c62_2;
  wire [7:0] t_r22_c62_3;
  wire [7:0] t_r22_c62_4;
  wire [7:0] t_r22_c62_5;
  wire [7:0] t_r22_c62_6;
  wire [7:0] t_r22_c62_7;
  wire [7:0] t_r22_c62_8;
  wire [7:0] t_r22_c62_9;
  wire [7:0] t_r22_c62_10;
  wire [7:0] t_r22_c62_11;
  wire [7:0] t_r22_c62_12;
  wire [7:0] t_r22_c63_0;
  wire [7:0] t_r22_c63_1;
  wire [7:0] t_r22_c63_2;
  wire [7:0] t_r22_c63_3;
  wire [7:0] t_r22_c63_4;
  wire [7:0] t_r22_c63_5;
  wire [7:0] t_r22_c63_6;
  wire [7:0] t_r22_c63_7;
  wire [7:0] t_r22_c63_8;
  wire [7:0] t_r22_c63_9;
  wire [7:0] t_r22_c63_10;
  wire [7:0] t_r22_c63_11;
  wire [7:0] t_r22_c63_12;
  wire [7:0] t_r22_c64_0;
  wire [7:0] t_r22_c64_1;
  wire [7:0] t_r22_c64_2;
  wire [7:0] t_r22_c64_3;
  wire [7:0] t_r22_c64_4;
  wire [7:0] t_r22_c64_5;
  wire [7:0] t_r22_c64_6;
  wire [7:0] t_r22_c64_7;
  wire [7:0] t_r22_c64_8;
  wire [7:0] t_r22_c64_9;
  wire [7:0] t_r22_c64_10;
  wire [7:0] t_r22_c64_11;
  wire [7:0] t_r22_c64_12;
  wire [7:0] t_r22_c65_0;
  wire [7:0] t_r22_c65_1;
  wire [7:0] t_r22_c65_2;
  wire [7:0] t_r22_c65_3;
  wire [7:0] t_r22_c65_4;
  wire [7:0] t_r22_c65_5;
  wire [7:0] t_r22_c65_6;
  wire [7:0] t_r22_c65_7;
  wire [7:0] t_r22_c65_8;
  wire [7:0] t_r22_c65_9;
  wire [7:0] t_r22_c65_10;
  wire [7:0] t_r22_c65_11;
  wire [7:0] t_r22_c65_12;
  wire [7:0] t_r23_c0_0;
  wire [7:0] t_r23_c0_1;
  wire [7:0] t_r23_c0_2;
  wire [7:0] t_r23_c0_3;
  wire [7:0] t_r23_c0_4;
  wire [7:0] t_r23_c0_5;
  wire [7:0] t_r23_c0_6;
  wire [7:0] t_r23_c0_7;
  wire [7:0] t_r23_c0_8;
  wire [7:0] t_r23_c0_9;
  wire [7:0] t_r23_c0_10;
  wire [7:0] t_r23_c0_11;
  wire [7:0] t_r23_c0_12;
  wire [7:0] t_r23_c1_0;
  wire [7:0] t_r23_c1_1;
  wire [7:0] t_r23_c1_2;
  wire [7:0] t_r23_c1_3;
  wire [7:0] t_r23_c1_4;
  wire [7:0] t_r23_c1_5;
  wire [7:0] t_r23_c1_6;
  wire [7:0] t_r23_c1_7;
  wire [7:0] t_r23_c1_8;
  wire [7:0] t_r23_c1_9;
  wire [7:0] t_r23_c1_10;
  wire [7:0] t_r23_c1_11;
  wire [7:0] t_r23_c1_12;
  wire [7:0] t_r23_c2_0;
  wire [7:0] t_r23_c2_1;
  wire [7:0] t_r23_c2_2;
  wire [7:0] t_r23_c2_3;
  wire [7:0] t_r23_c2_4;
  wire [7:0] t_r23_c2_5;
  wire [7:0] t_r23_c2_6;
  wire [7:0] t_r23_c2_7;
  wire [7:0] t_r23_c2_8;
  wire [7:0] t_r23_c2_9;
  wire [7:0] t_r23_c2_10;
  wire [7:0] t_r23_c2_11;
  wire [7:0] t_r23_c2_12;
  wire [7:0] t_r23_c3_0;
  wire [7:0] t_r23_c3_1;
  wire [7:0] t_r23_c3_2;
  wire [7:0] t_r23_c3_3;
  wire [7:0] t_r23_c3_4;
  wire [7:0] t_r23_c3_5;
  wire [7:0] t_r23_c3_6;
  wire [7:0] t_r23_c3_7;
  wire [7:0] t_r23_c3_8;
  wire [7:0] t_r23_c3_9;
  wire [7:0] t_r23_c3_10;
  wire [7:0] t_r23_c3_11;
  wire [7:0] t_r23_c3_12;
  wire [7:0] t_r23_c4_0;
  wire [7:0] t_r23_c4_1;
  wire [7:0] t_r23_c4_2;
  wire [7:0] t_r23_c4_3;
  wire [7:0] t_r23_c4_4;
  wire [7:0] t_r23_c4_5;
  wire [7:0] t_r23_c4_6;
  wire [7:0] t_r23_c4_7;
  wire [7:0] t_r23_c4_8;
  wire [7:0] t_r23_c4_9;
  wire [7:0] t_r23_c4_10;
  wire [7:0] t_r23_c4_11;
  wire [7:0] t_r23_c4_12;
  wire [7:0] t_r23_c5_0;
  wire [7:0] t_r23_c5_1;
  wire [7:0] t_r23_c5_2;
  wire [7:0] t_r23_c5_3;
  wire [7:0] t_r23_c5_4;
  wire [7:0] t_r23_c5_5;
  wire [7:0] t_r23_c5_6;
  wire [7:0] t_r23_c5_7;
  wire [7:0] t_r23_c5_8;
  wire [7:0] t_r23_c5_9;
  wire [7:0] t_r23_c5_10;
  wire [7:0] t_r23_c5_11;
  wire [7:0] t_r23_c5_12;
  wire [7:0] t_r23_c6_0;
  wire [7:0] t_r23_c6_1;
  wire [7:0] t_r23_c6_2;
  wire [7:0] t_r23_c6_3;
  wire [7:0] t_r23_c6_4;
  wire [7:0] t_r23_c6_5;
  wire [7:0] t_r23_c6_6;
  wire [7:0] t_r23_c6_7;
  wire [7:0] t_r23_c6_8;
  wire [7:0] t_r23_c6_9;
  wire [7:0] t_r23_c6_10;
  wire [7:0] t_r23_c6_11;
  wire [7:0] t_r23_c6_12;
  wire [7:0] t_r23_c7_0;
  wire [7:0] t_r23_c7_1;
  wire [7:0] t_r23_c7_2;
  wire [7:0] t_r23_c7_3;
  wire [7:0] t_r23_c7_4;
  wire [7:0] t_r23_c7_5;
  wire [7:0] t_r23_c7_6;
  wire [7:0] t_r23_c7_7;
  wire [7:0] t_r23_c7_8;
  wire [7:0] t_r23_c7_9;
  wire [7:0] t_r23_c7_10;
  wire [7:0] t_r23_c7_11;
  wire [7:0] t_r23_c7_12;
  wire [7:0] t_r23_c8_0;
  wire [7:0] t_r23_c8_1;
  wire [7:0] t_r23_c8_2;
  wire [7:0] t_r23_c8_3;
  wire [7:0] t_r23_c8_4;
  wire [7:0] t_r23_c8_5;
  wire [7:0] t_r23_c8_6;
  wire [7:0] t_r23_c8_7;
  wire [7:0] t_r23_c8_8;
  wire [7:0] t_r23_c8_9;
  wire [7:0] t_r23_c8_10;
  wire [7:0] t_r23_c8_11;
  wire [7:0] t_r23_c8_12;
  wire [7:0] t_r23_c9_0;
  wire [7:0] t_r23_c9_1;
  wire [7:0] t_r23_c9_2;
  wire [7:0] t_r23_c9_3;
  wire [7:0] t_r23_c9_4;
  wire [7:0] t_r23_c9_5;
  wire [7:0] t_r23_c9_6;
  wire [7:0] t_r23_c9_7;
  wire [7:0] t_r23_c9_8;
  wire [7:0] t_r23_c9_9;
  wire [7:0] t_r23_c9_10;
  wire [7:0] t_r23_c9_11;
  wire [7:0] t_r23_c9_12;
  wire [7:0] t_r23_c10_0;
  wire [7:0] t_r23_c10_1;
  wire [7:0] t_r23_c10_2;
  wire [7:0] t_r23_c10_3;
  wire [7:0] t_r23_c10_4;
  wire [7:0] t_r23_c10_5;
  wire [7:0] t_r23_c10_6;
  wire [7:0] t_r23_c10_7;
  wire [7:0] t_r23_c10_8;
  wire [7:0] t_r23_c10_9;
  wire [7:0] t_r23_c10_10;
  wire [7:0] t_r23_c10_11;
  wire [7:0] t_r23_c10_12;
  wire [7:0] t_r23_c11_0;
  wire [7:0] t_r23_c11_1;
  wire [7:0] t_r23_c11_2;
  wire [7:0] t_r23_c11_3;
  wire [7:0] t_r23_c11_4;
  wire [7:0] t_r23_c11_5;
  wire [7:0] t_r23_c11_6;
  wire [7:0] t_r23_c11_7;
  wire [7:0] t_r23_c11_8;
  wire [7:0] t_r23_c11_9;
  wire [7:0] t_r23_c11_10;
  wire [7:0] t_r23_c11_11;
  wire [7:0] t_r23_c11_12;
  wire [7:0] t_r23_c12_0;
  wire [7:0] t_r23_c12_1;
  wire [7:0] t_r23_c12_2;
  wire [7:0] t_r23_c12_3;
  wire [7:0] t_r23_c12_4;
  wire [7:0] t_r23_c12_5;
  wire [7:0] t_r23_c12_6;
  wire [7:0] t_r23_c12_7;
  wire [7:0] t_r23_c12_8;
  wire [7:0] t_r23_c12_9;
  wire [7:0] t_r23_c12_10;
  wire [7:0] t_r23_c12_11;
  wire [7:0] t_r23_c12_12;
  wire [7:0] t_r23_c13_0;
  wire [7:0] t_r23_c13_1;
  wire [7:0] t_r23_c13_2;
  wire [7:0] t_r23_c13_3;
  wire [7:0] t_r23_c13_4;
  wire [7:0] t_r23_c13_5;
  wire [7:0] t_r23_c13_6;
  wire [7:0] t_r23_c13_7;
  wire [7:0] t_r23_c13_8;
  wire [7:0] t_r23_c13_9;
  wire [7:0] t_r23_c13_10;
  wire [7:0] t_r23_c13_11;
  wire [7:0] t_r23_c13_12;
  wire [7:0] t_r23_c14_0;
  wire [7:0] t_r23_c14_1;
  wire [7:0] t_r23_c14_2;
  wire [7:0] t_r23_c14_3;
  wire [7:0] t_r23_c14_4;
  wire [7:0] t_r23_c14_5;
  wire [7:0] t_r23_c14_6;
  wire [7:0] t_r23_c14_7;
  wire [7:0] t_r23_c14_8;
  wire [7:0] t_r23_c14_9;
  wire [7:0] t_r23_c14_10;
  wire [7:0] t_r23_c14_11;
  wire [7:0] t_r23_c14_12;
  wire [7:0] t_r23_c15_0;
  wire [7:0] t_r23_c15_1;
  wire [7:0] t_r23_c15_2;
  wire [7:0] t_r23_c15_3;
  wire [7:0] t_r23_c15_4;
  wire [7:0] t_r23_c15_5;
  wire [7:0] t_r23_c15_6;
  wire [7:0] t_r23_c15_7;
  wire [7:0] t_r23_c15_8;
  wire [7:0] t_r23_c15_9;
  wire [7:0] t_r23_c15_10;
  wire [7:0] t_r23_c15_11;
  wire [7:0] t_r23_c15_12;
  wire [7:0] t_r23_c16_0;
  wire [7:0] t_r23_c16_1;
  wire [7:0] t_r23_c16_2;
  wire [7:0] t_r23_c16_3;
  wire [7:0] t_r23_c16_4;
  wire [7:0] t_r23_c16_5;
  wire [7:0] t_r23_c16_6;
  wire [7:0] t_r23_c16_7;
  wire [7:0] t_r23_c16_8;
  wire [7:0] t_r23_c16_9;
  wire [7:0] t_r23_c16_10;
  wire [7:0] t_r23_c16_11;
  wire [7:0] t_r23_c16_12;
  wire [7:0] t_r23_c17_0;
  wire [7:0] t_r23_c17_1;
  wire [7:0] t_r23_c17_2;
  wire [7:0] t_r23_c17_3;
  wire [7:0] t_r23_c17_4;
  wire [7:0] t_r23_c17_5;
  wire [7:0] t_r23_c17_6;
  wire [7:0] t_r23_c17_7;
  wire [7:0] t_r23_c17_8;
  wire [7:0] t_r23_c17_9;
  wire [7:0] t_r23_c17_10;
  wire [7:0] t_r23_c17_11;
  wire [7:0] t_r23_c17_12;
  wire [7:0] t_r23_c18_0;
  wire [7:0] t_r23_c18_1;
  wire [7:0] t_r23_c18_2;
  wire [7:0] t_r23_c18_3;
  wire [7:0] t_r23_c18_4;
  wire [7:0] t_r23_c18_5;
  wire [7:0] t_r23_c18_6;
  wire [7:0] t_r23_c18_7;
  wire [7:0] t_r23_c18_8;
  wire [7:0] t_r23_c18_9;
  wire [7:0] t_r23_c18_10;
  wire [7:0] t_r23_c18_11;
  wire [7:0] t_r23_c18_12;
  wire [7:0] t_r23_c19_0;
  wire [7:0] t_r23_c19_1;
  wire [7:0] t_r23_c19_2;
  wire [7:0] t_r23_c19_3;
  wire [7:0] t_r23_c19_4;
  wire [7:0] t_r23_c19_5;
  wire [7:0] t_r23_c19_6;
  wire [7:0] t_r23_c19_7;
  wire [7:0] t_r23_c19_8;
  wire [7:0] t_r23_c19_9;
  wire [7:0] t_r23_c19_10;
  wire [7:0] t_r23_c19_11;
  wire [7:0] t_r23_c19_12;
  wire [7:0] t_r23_c20_0;
  wire [7:0] t_r23_c20_1;
  wire [7:0] t_r23_c20_2;
  wire [7:0] t_r23_c20_3;
  wire [7:0] t_r23_c20_4;
  wire [7:0] t_r23_c20_5;
  wire [7:0] t_r23_c20_6;
  wire [7:0] t_r23_c20_7;
  wire [7:0] t_r23_c20_8;
  wire [7:0] t_r23_c20_9;
  wire [7:0] t_r23_c20_10;
  wire [7:0] t_r23_c20_11;
  wire [7:0] t_r23_c20_12;
  wire [7:0] t_r23_c21_0;
  wire [7:0] t_r23_c21_1;
  wire [7:0] t_r23_c21_2;
  wire [7:0] t_r23_c21_3;
  wire [7:0] t_r23_c21_4;
  wire [7:0] t_r23_c21_5;
  wire [7:0] t_r23_c21_6;
  wire [7:0] t_r23_c21_7;
  wire [7:0] t_r23_c21_8;
  wire [7:0] t_r23_c21_9;
  wire [7:0] t_r23_c21_10;
  wire [7:0] t_r23_c21_11;
  wire [7:0] t_r23_c21_12;
  wire [7:0] t_r23_c22_0;
  wire [7:0] t_r23_c22_1;
  wire [7:0] t_r23_c22_2;
  wire [7:0] t_r23_c22_3;
  wire [7:0] t_r23_c22_4;
  wire [7:0] t_r23_c22_5;
  wire [7:0] t_r23_c22_6;
  wire [7:0] t_r23_c22_7;
  wire [7:0] t_r23_c22_8;
  wire [7:0] t_r23_c22_9;
  wire [7:0] t_r23_c22_10;
  wire [7:0] t_r23_c22_11;
  wire [7:0] t_r23_c22_12;
  wire [7:0] t_r23_c23_0;
  wire [7:0] t_r23_c23_1;
  wire [7:0] t_r23_c23_2;
  wire [7:0] t_r23_c23_3;
  wire [7:0] t_r23_c23_4;
  wire [7:0] t_r23_c23_5;
  wire [7:0] t_r23_c23_6;
  wire [7:0] t_r23_c23_7;
  wire [7:0] t_r23_c23_8;
  wire [7:0] t_r23_c23_9;
  wire [7:0] t_r23_c23_10;
  wire [7:0] t_r23_c23_11;
  wire [7:0] t_r23_c23_12;
  wire [7:0] t_r23_c24_0;
  wire [7:0] t_r23_c24_1;
  wire [7:0] t_r23_c24_2;
  wire [7:0] t_r23_c24_3;
  wire [7:0] t_r23_c24_4;
  wire [7:0] t_r23_c24_5;
  wire [7:0] t_r23_c24_6;
  wire [7:0] t_r23_c24_7;
  wire [7:0] t_r23_c24_8;
  wire [7:0] t_r23_c24_9;
  wire [7:0] t_r23_c24_10;
  wire [7:0] t_r23_c24_11;
  wire [7:0] t_r23_c24_12;
  wire [7:0] t_r23_c25_0;
  wire [7:0] t_r23_c25_1;
  wire [7:0] t_r23_c25_2;
  wire [7:0] t_r23_c25_3;
  wire [7:0] t_r23_c25_4;
  wire [7:0] t_r23_c25_5;
  wire [7:0] t_r23_c25_6;
  wire [7:0] t_r23_c25_7;
  wire [7:0] t_r23_c25_8;
  wire [7:0] t_r23_c25_9;
  wire [7:0] t_r23_c25_10;
  wire [7:0] t_r23_c25_11;
  wire [7:0] t_r23_c25_12;
  wire [7:0] t_r23_c26_0;
  wire [7:0] t_r23_c26_1;
  wire [7:0] t_r23_c26_2;
  wire [7:0] t_r23_c26_3;
  wire [7:0] t_r23_c26_4;
  wire [7:0] t_r23_c26_5;
  wire [7:0] t_r23_c26_6;
  wire [7:0] t_r23_c26_7;
  wire [7:0] t_r23_c26_8;
  wire [7:0] t_r23_c26_9;
  wire [7:0] t_r23_c26_10;
  wire [7:0] t_r23_c26_11;
  wire [7:0] t_r23_c26_12;
  wire [7:0] t_r23_c27_0;
  wire [7:0] t_r23_c27_1;
  wire [7:0] t_r23_c27_2;
  wire [7:0] t_r23_c27_3;
  wire [7:0] t_r23_c27_4;
  wire [7:0] t_r23_c27_5;
  wire [7:0] t_r23_c27_6;
  wire [7:0] t_r23_c27_7;
  wire [7:0] t_r23_c27_8;
  wire [7:0] t_r23_c27_9;
  wire [7:0] t_r23_c27_10;
  wire [7:0] t_r23_c27_11;
  wire [7:0] t_r23_c27_12;
  wire [7:0] t_r23_c28_0;
  wire [7:0] t_r23_c28_1;
  wire [7:0] t_r23_c28_2;
  wire [7:0] t_r23_c28_3;
  wire [7:0] t_r23_c28_4;
  wire [7:0] t_r23_c28_5;
  wire [7:0] t_r23_c28_6;
  wire [7:0] t_r23_c28_7;
  wire [7:0] t_r23_c28_8;
  wire [7:0] t_r23_c28_9;
  wire [7:0] t_r23_c28_10;
  wire [7:0] t_r23_c28_11;
  wire [7:0] t_r23_c28_12;
  wire [7:0] t_r23_c29_0;
  wire [7:0] t_r23_c29_1;
  wire [7:0] t_r23_c29_2;
  wire [7:0] t_r23_c29_3;
  wire [7:0] t_r23_c29_4;
  wire [7:0] t_r23_c29_5;
  wire [7:0] t_r23_c29_6;
  wire [7:0] t_r23_c29_7;
  wire [7:0] t_r23_c29_8;
  wire [7:0] t_r23_c29_9;
  wire [7:0] t_r23_c29_10;
  wire [7:0] t_r23_c29_11;
  wire [7:0] t_r23_c29_12;
  wire [7:0] t_r23_c30_0;
  wire [7:0] t_r23_c30_1;
  wire [7:0] t_r23_c30_2;
  wire [7:0] t_r23_c30_3;
  wire [7:0] t_r23_c30_4;
  wire [7:0] t_r23_c30_5;
  wire [7:0] t_r23_c30_6;
  wire [7:0] t_r23_c30_7;
  wire [7:0] t_r23_c30_8;
  wire [7:0] t_r23_c30_9;
  wire [7:0] t_r23_c30_10;
  wire [7:0] t_r23_c30_11;
  wire [7:0] t_r23_c30_12;
  wire [7:0] t_r23_c31_0;
  wire [7:0] t_r23_c31_1;
  wire [7:0] t_r23_c31_2;
  wire [7:0] t_r23_c31_3;
  wire [7:0] t_r23_c31_4;
  wire [7:0] t_r23_c31_5;
  wire [7:0] t_r23_c31_6;
  wire [7:0] t_r23_c31_7;
  wire [7:0] t_r23_c31_8;
  wire [7:0] t_r23_c31_9;
  wire [7:0] t_r23_c31_10;
  wire [7:0] t_r23_c31_11;
  wire [7:0] t_r23_c31_12;
  wire [7:0] t_r23_c32_0;
  wire [7:0] t_r23_c32_1;
  wire [7:0] t_r23_c32_2;
  wire [7:0] t_r23_c32_3;
  wire [7:0] t_r23_c32_4;
  wire [7:0] t_r23_c32_5;
  wire [7:0] t_r23_c32_6;
  wire [7:0] t_r23_c32_7;
  wire [7:0] t_r23_c32_8;
  wire [7:0] t_r23_c32_9;
  wire [7:0] t_r23_c32_10;
  wire [7:0] t_r23_c32_11;
  wire [7:0] t_r23_c32_12;
  wire [7:0] t_r23_c33_0;
  wire [7:0] t_r23_c33_1;
  wire [7:0] t_r23_c33_2;
  wire [7:0] t_r23_c33_3;
  wire [7:0] t_r23_c33_4;
  wire [7:0] t_r23_c33_5;
  wire [7:0] t_r23_c33_6;
  wire [7:0] t_r23_c33_7;
  wire [7:0] t_r23_c33_8;
  wire [7:0] t_r23_c33_9;
  wire [7:0] t_r23_c33_10;
  wire [7:0] t_r23_c33_11;
  wire [7:0] t_r23_c33_12;
  wire [7:0] t_r23_c34_0;
  wire [7:0] t_r23_c34_1;
  wire [7:0] t_r23_c34_2;
  wire [7:0] t_r23_c34_3;
  wire [7:0] t_r23_c34_4;
  wire [7:0] t_r23_c34_5;
  wire [7:0] t_r23_c34_6;
  wire [7:0] t_r23_c34_7;
  wire [7:0] t_r23_c34_8;
  wire [7:0] t_r23_c34_9;
  wire [7:0] t_r23_c34_10;
  wire [7:0] t_r23_c34_11;
  wire [7:0] t_r23_c34_12;
  wire [7:0] t_r23_c35_0;
  wire [7:0] t_r23_c35_1;
  wire [7:0] t_r23_c35_2;
  wire [7:0] t_r23_c35_3;
  wire [7:0] t_r23_c35_4;
  wire [7:0] t_r23_c35_5;
  wire [7:0] t_r23_c35_6;
  wire [7:0] t_r23_c35_7;
  wire [7:0] t_r23_c35_8;
  wire [7:0] t_r23_c35_9;
  wire [7:0] t_r23_c35_10;
  wire [7:0] t_r23_c35_11;
  wire [7:0] t_r23_c35_12;
  wire [7:0] t_r23_c36_0;
  wire [7:0] t_r23_c36_1;
  wire [7:0] t_r23_c36_2;
  wire [7:0] t_r23_c36_3;
  wire [7:0] t_r23_c36_4;
  wire [7:0] t_r23_c36_5;
  wire [7:0] t_r23_c36_6;
  wire [7:0] t_r23_c36_7;
  wire [7:0] t_r23_c36_8;
  wire [7:0] t_r23_c36_9;
  wire [7:0] t_r23_c36_10;
  wire [7:0] t_r23_c36_11;
  wire [7:0] t_r23_c36_12;
  wire [7:0] t_r23_c37_0;
  wire [7:0] t_r23_c37_1;
  wire [7:0] t_r23_c37_2;
  wire [7:0] t_r23_c37_3;
  wire [7:0] t_r23_c37_4;
  wire [7:0] t_r23_c37_5;
  wire [7:0] t_r23_c37_6;
  wire [7:0] t_r23_c37_7;
  wire [7:0] t_r23_c37_8;
  wire [7:0] t_r23_c37_9;
  wire [7:0] t_r23_c37_10;
  wire [7:0] t_r23_c37_11;
  wire [7:0] t_r23_c37_12;
  wire [7:0] t_r23_c38_0;
  wire [7:0] t_r23_c38_1;
  wire [7:0] t_r23_c38_2;
  wire [7:0] t_r23_c38_3;
  wire [7:0] t_r23_c38_4;
  wire [7:0] t_r23_c38_5;
  wire [7:0] t_r23_c38_6;
  wire [7:0] t_r23_c38_7;
  wire [7:0] t_r23_c38_8;
  wire [7:0] t_r23_c38_9;
  wire [7:0] t_r23_c38_10;
  wire [7:0] t_r23_c38_11;
  wire [7:0] t_r23_c38_12;
  wire [7:0] t_r23_c39_0;
  wire [7:0] t_r23_c39_1;
  wire [7:0] t_r23_c39_2;
  wire [7:0] t_r23_c39_3;
  wire [7:0] t_r23_c39_4;
  wire [7:0] t_r23_c39_5;
  wire [7:0] t_r23_c39_6;
  wire [7:0] t_r23_c39_7;
  wire [7:0] t_r23_c39_8;
  wire [7:0] t_r23_c39_9;
  wire [7:0] t_r23_c39_10;
  wire [7:0] t_r23_c39_11;
  wire [7:0] t_r23_c39_12;
  wire [7:0] t_r23_c40_0;
  wire [7:0] t_r23_c40_1;
  wire [7:0] t_r23_c40_2;
  wire [7:0] t_r23_c40_3;
  wire [7:0] t_r23_c40_4;
  wire [7:0] t_r23_c40_5;
  wire [7:0] t_r23_c40_6;
  wire [7:0] t_r23_c40_7;
  wire [7:0] t_r23_c40_8;
  wire [7:0] t_r23_c40_9;
  wire [7:0] t_r23_c40_10;
  wire [7:0] t_r23_c40_11;
  wire [7:0] t_r23_c40_12;
  wire [7:0] t_r23_c41_0;
  wire [7:0] t_r23_c41_1;
  wire [7:0] t_r23_c41_2;
  wire [7:0] t_r23_c41_3;
  wire [7:0] t_r23_c41_4;
  wire [7:0] t_r23_c41_5;
  wire [7:0] t_r23_c41_6;
  wire [7:0] t_r23_c41_7;
  wire [7:0] t_r23_c41_8;
  wire [7:0] t_r23_c41_9;
  wire [7:0] t_r23_c41_10;
  wire [7:0] t_r23_c41_11;
  wire [7:0] t_r23_c41_12;
  wire [7:0] t_r23_c42_0;
  wire [7:0] t_r23_c42_1;
  wire [7:0] t_r23_c42_2;
  wire [7:0] t_r23_c42_3;
  wire [7:0] t_r23_c42_4;
  wire [7:0] t_r23_c42_5;
  wire [7:0] t_r23_c42_6;
  wire [7:0] t_r23_c42_7;
  wire [7:0] t_r23_c42_8;
  wire [7:0] t_r23_c42_9;
  wire [7:0] t_r23_c42_10;
  wire [7:0] t_r23_c42_11;
  wire [7:0] t_r23_c42_12;
  wire [7:0] t_r23_c43_0;
  wire [7:0] t_r23_c43_1;
  wire [7:0] t_r23_c43_2;
  wire [7:0] t_r23_c43_3;
  wire [7:0] t_r23_c43_4;
  wire [7:0] t_r23_c43_5;
  wire [7:0] t_r23_c43_6;
  wire [7:0] t_r23_c43_7;
  wire [7:0] t_r23_c43_8;
  wire [7:0] t_r23_c43_9;
  wire [7:0] t_r23_c43_10;
  wire [7:0] t_r23_c43_11;
  wire [7:0] t_r23_c43_12;
  wire [7:0] t_r23_c44_0;
  wire [7:0] t_r23_c44_1;
  wire [7:0] t_r23_c44_2;
  wire [7:0] t_r23_c44_3;
  wire [7:0] t_r23_c44_4;
  wire [7:0] t_r23_c44_5;
  wire [7:0] t_r23_c44_6;
  wire [7:0] t_r23_c44_7;
  wire [7:0] t_r23_c44_8;
  wire [7:0] t_r23_c44_9;
  wire [7:0] t_r23_c44_10;
  wire [7:0] t_r23_c44_11;
  wire [7:0] t_r23_c44_12;
  wire [7:0] t_r23_c45_0;
  wire [7:0] t_r23_c45_1;
  wire [7:0] t_r23_c45_2;
  wire [7:0] t_r23_c45_3;
  wire [7:0] t_r23_c45_4;
  wire [7:0] t_r23_c45_5;
  wire [7:0] t_r23_c45_6;
  wire [7:0] t_r23_c45_7;
  wire [7:0] t_r23_c45_8;
  wire [7:0] t_r23_c45_9;
  wire [7:0] t_r23_c45_10;
  wire [7:0] t_r23_c45_11;
  wire [7:0] t_r23_c45_12;
  wire [7:0] t_r23_c46_0;
  wire [7:0] t_r23_c46_1;
  wire [7:0] t_r23_c46_2;
  wire [7:0] t_r23_c46_3;
  wire [7:0] t_r23_c46_4;
  wire [7:0] t_r23_c46_5;
  wire [7:0] t_r23_c46_6;
  wire [7:0] t_r23_c46_7;
  wire [7:0] t_r23_c46_8;
  wire [7:0] t_r23_c46_9;
  wire [7:0] t_r23_c46_10;
  wire [7:0] t_r23_c46_11;
  wire [7:0] t_r23_c46_12;
  wire [7:0] t_r23_c47_0;
  wire [7:0] t_r23_c47_1;
  wire [7:0] t_r23_c47_2;
  wire [7:0] t_r23_c47_3;
  wire [7:0] t_r23_c47_4;
  wire [7:0] t_r23_c47_5;
  wire [7:0] t_r23_c47_6;
  wire [7:0] t_r23_c47_7;
  wire [7:0] t_r23_c47_8;
  wire [7:0] t_r23_c47_9;
  wire [7:0] t_r23_c47_10;
  wire [7:0] t_r23_c47_11;
  wire [7:0] t_r23_c47_12;
  wire [7:0] t_r23_c48_0;
  wire [7:0] t_r23_c48_1;
  wire [7:0] t_r23_c48_2;
  wire [7:0] t_r23_c48_3;
  wire [7:0] t_r23_c48_4;
  wire [7:0] t_r23_c48_5;
  wire [7:0] t_r23_c48_6;
  wire [7:0] t_r23_c48_7;
  wire [7:0] t_r23_c48_8;
  wire [7:0] t_r23_c48_9;
  wire [7:0] t_r23_c48_10;
  wire [7:0] t_r23_c48_11;
  wire [7:0] t_r23_c48_12;
  wire [7:0] t_r23_c49_0;
  wire [7:0] t_r23_c49_1;
  wire [7:0] t_r23_c49_2;
  wire [7:0] t_r23_c49_3;
  wire [7:0] t_r23_c49_4;
  wire [7:0] t_r23_c49_5;
  wire [7:0] t_r23_c49_6;
  wire [7:0] t_r23_c49_7;
  wire [7:0] t_r23_c49_8;
  wire [7:0] t_r23_c49_9;
  wire [7:0] t_r23_c49_10;
  wire [7:0] t_r23_c49_11;
  wire [7:0] t_r23_c49_12;
  wire [7:0] t_r23_c50_0;
  wire [7:0] t_r23_c50_1;
  wire [7:0] t_r23_c50_2;
  wire [7:0] t_r23_c50_3;
  wire [7:0] t_r23_c50_4;
  wire [7:0] t_r23_c50_5;
  wire [7:0] t_r23_c50_6;
  wire [7:0] t_r23_c50_7;
  wire [7:0] t_r23_c50_8;
  wire [7:0] t_r23_c50_9;
  wire [7:0] t_r23_c50_10;
  wire [7:0] t_r23_c50_11;
  wire [7:0] t_r23_c50_12;
  wire [7:0] t_r23_c51_0;
  wire [7:0] t_r23_c51_1;
  wire [7:0] t_r23_c51_2;
  wire [7:0] t_r23_c51_3;
  wire [7:0] t_r23_c51_4;
  wire [7:0] t_r23_c51_5;
  wire [7:0] t_r23_c51_6;
  wire [7:0] t_r23_c51_7;
  wire [7:0] t_r23_c51_8;
  wire [7:0] t_r23_c51_9;
  wire [7:0] t_r23_c51_10;
  wire [7:0] t_r23_c51_11;
  wire [7:0] t_r23_c51_12;
  wire [7:0] t_r23_c52_0;
  wire [7:0] t_r23_c52_1;
  wire [7:0] t_r23_c52_2;
  wire [7:0] t_r23_c52_3;
  wire [7:0] t_r23_c52_4;
  wire [7:0] t_r23_c52_5;
  wire [7:0] t_r23_c52_6;
  wire [7:0] t_r23_c52_7;
  wire [7:0] t_r23_c52_8;
  wire [7:0] t_r23_c52_9;
  wire [7:0] t_r23_c52_10;
  wire [7:0] t_r23_c52_11;
  wire [7:0] t_r23_c52_12;
  wire [7:0] t_r23_c53_0;
  wire [7:0] t_r23_c53_1;
  wire [7:0] t_r23_c53_2;
  wire [7:0] t_r23_c53_3;
  wire [7:0] t_r23_c53_4;
  wire [7:0] t_r23_c53_5;
  wire [7:0] t_r23_c53_6;
  wire [7:0] t_r23_c53_7;
  wire [7:0] t_r23_c53_8;
  wire [7:0] t_r23_c53_9;
  wire [7:0] t_r23_c53_10;
  wire [7:0] t_r23_c53_11;
  wire [7:0] t_r23_c53_12;
  wire [7:0] t_r23_c54_0;
  wire [7:0] t_r23_c54_1;
  wire [7:0] t_r23_c54_2;
  wire [7:0] t_r23_c54_3;
  wire [7:0] t_r23_c54_4;
  wire [7:0] t_r23_c54_5;
  wire [7:0] t_r23_c54_6;
  wire [7:0] t_r23_c54_7;
  wire [7:0] t_r23_c54_8;
  wire [7:0] t_r23_c54_9;
  wire [7:0] t_r23_c54_10;
  wire [7:0] t_r23_c54_11;
  wire [7:0] t_r23_c54_12;
  wire [7:0] t_r23_c55_0;
  wire [7:0] t_r23_c55_1;
  wire [7:0] t_r23_c55_2;
  wire [7:0] t_r23_c55_3;
  wire [7:0] t_r23_c55_4;
  wire [7:0] t_r23_c55_5;
  wire [7:0] t_r23_c55_6;
  wire [7:0] t_r23_c55_7;
  wire [7:0] t_r23_c55_8;
  wire [7:0] t_r23_c55_9;
  wire [7:0] t_r23_c55_10;
  wire [7:0] t_r23_c55_11;
  wire [7:0] t_r23_c55_12;
  wire [7:0] t_r23_c56_0;
  wire [7:0] t_r23_c56_1;
  wire [7:0] t_r23_c56_2;
  wire [7:0] t_r23_c56_3;
  wire [7:0] t_r23_c56_4;
  wire [7:0] t_r23_c56_5;
  wire [7:0] t_r23_c56_6;
  wire [7:0] t_r23_c56_7;
  wire [7:0] t_r23_c56_8;
  wire [7:0] t_r23_c56_9;
  wire [7:0] t_r23_c56_10;
  wire [7:0] t_r23_c56_11;
  wire [7:0] t_r23_c56_12;
  wire [7:0] t_r23_c57_0;
  wire [7:0] t_r23_c57_1;
  wire [7:0] t_r23_c57_2;
  wire [7:0] t_r23_c57_3;
  wire [7:0] t_r23_c57_4;
  wire [7:0] t_r23_c57_5;
  wire [7:0] t_r23_c57_6;
  wire [7:0] t_r23_c57_7;
  wire [7:0] t_r23_c57_8;
  wire [7:0] t_r23_c57_9;
  wire [7:0] t_r23_c57_10;
  wire [7:0] t_r23_c57_11;
  wire [7:0] t_r23_c57_12;
  wire [7:0] t_r23_c58_0;
  wire [7:0] t_r23_c58_1;
  wire [7:0] t_r23_c58_2;
  wire [7:0] t_r23_c58_3;
  wire [7:0] t_r23_c58_4;
  wire [7:0] t_r23_c58_5;
  wire [7:0] t_r23_c58_6;
  wire [7:0] t_r23_c58_7;
  wire [7:0] t_r23_c58_8;
  wire [7:0] t_r23_c58_9;
  wire [7:0] t_r23_c58_10;
  wire [7:0] t_r23_c58_11;
  wire [7:0] t_r23_c58_12;
  wire [7:0] t_r23_c59_0;
  wire [7:0] t_r23_c59_1;
  wire [7:0] t_r23_c59_2;
  wire [7:0] t_r23_c59_3;
  wire [7:0] t_r23_c59_4;
  wire [7:0] t_r23_c59_5;
  wire [7:0] t_r23_c59_6;
  wire [7:0] t_r23_c59_7;
  wire [7:0] t_r23_c59_8;
  wire [7:0] t_r23_c59_9;
  wire [7:0] t_r23_c59_10;
  wire [7:0] t_r23_c59_11;
  wire [7:0] t_r23_c59_12;
  wire [7:0] t_r23_c60_0;
  wire [7:0] t_r23_c60_1;
  wire [7:0] t_r23_c60_2;
  wire [7:0] t_r23_c60_3;
  wire [7:0] t_r23_c60_4;
  wire [7:0] t_r23_c60_5;
  wire [7:0] t_r23_c60_6;
  wire [7:0] t_r23_c60_7;
  wire [7:0] t_r23_c60_8;
  wire [7:0] t_r23_c60_9;
  wire [7:0] t_r23_c60_10;
  wire [7:0] t_r23_c60_11;
  wire [7:0] t_r23_c60_12;
  wire [7:0] t_r23_c61_0;
  wire [7:0] t_r23_c61_1;
  wire [7:0] t_r23_c61_2;
  wire [7:0] t_r23_c61_3;
  wire [7:0] t_r23_c61_4;
  wire [7:0] t_r23_c61_5;
  wire [7:0] t_r23_c61_6;
  wire [7:0] t_r23_c61_7;
  wire [7:0] t_r23_c61_8;
  wire [7:0] t_r23_c61_9;
  wire [7:0] t_r23_c61_10;
  wire [7:0] t_r23_c61_11;
  wire [7:0] t_r23_c61_12;
  wire [7:0] t_r23_c62_0;
  wire [7:0] t_r23_c62_1;
  wire [7:0] t_r23_c62_2;
  wire [7:0] t_r23_c62_3;
  wire [7:0] t_r23_c62_4;
  wire [7:0] t_r23_c62_5;
  wire [7:0] t_r23_c62_6;
  wire [7:0] t_r23_c62_7;
  wire [7:0] t_r23_c62_8;
  wire [7:0] t_r23_c62_9;
  wire [7:0] t_r23_c62_10;
  wire [7:0] t_r23_c62_11;
  wire [7:0] t_r23_c62_12;
  wire [7:0] t_r23_c63_0;
  wire [7:0] t_r23_c63_1;
  wire [7:0] t_r23_c63_2;
  wire [7:0] t_r23_c63_3;
  wire [7:0] t_r23_c63_4;
  wire [7:0] t_r23_c63_5;
  wire [7:0] t_r23_c63_6;
  wire [7:0] t_r23_c63_7;
  wire [7:0] t_r23_c63_8;
  wire [7:0] t_r23_c63_9;
  wire [7:0] t_r23_c63_10;
  wire [7:0] t_r23_c63_11;
  wire [7:0] t_r23_c63_12;
  wire [7:0] t_r23_c64_0;
  wire [7:0] t_r23_c64_1;
  wire [7:0] t_r23_c64_2;
  wire [7:0] t_r23_c64_3;
  wire [7:0] t_r23_c64_4;
  wire [7:0] t_r23_c64_5;
  wire [7:0] t_r23_c64_6;
  wire [7:0] t_r23_c64_7;
  wire [7:0] t_r23_c64_8;
  wire [7:0] t_r23_c64_9;
  wire [7:0] t_r23_c64_10;
  wire [7:0] t_r23_c64_11;
  wire [7:0] t_r23_c64_12;
  wire [7:0] t_r23_c65_0;
  wire [7:0] t_r23_c65_1;
  wire [7:0] t_r23_c65_2;
  wire [7:0] t_r23_c65_3;
  wire [7:0] t_r23_c65_4;
  wire [7:0] t_r23_c65_5;
  wire [7:0] t_r23_c65_6;
  wire [7:0] t_r23_c65_7;
  wire [7:0] t_r23_c65_8;
  wire [7:0] t_r23_c65_9;
  wire [7:0] t_r23_c65_10;
  wire [7:0] t_r23_c65_11;
  wire [7:0] t_r23_c65_12;
  wire [7:0] t_r24_c0_0;
  wire [7:0] t_r24_c0_1;
  wire [7:0] t_r24_c0_2;
  wire [7:0] t_r24_c0_3;
  wire [7:0] t_r24_c0_4;
  wire [7:0] t_r24_c0_5;
  wire [7:0] t_r24_c0_6;
  wire [7:0] t_r24_c0_7;
  wire [7:0] t_r24_c0_8;
  wire [7:0] t_r24_c0_9;
  wire [7:0] t_r24_c0_10;
  wire [7:0] t_r24_c0_11;
  wire [7:0] t_r24_c0_12;
  wire [7:0] t_r24_c1_0;
  wire [7:0] t_r24_c1_1;
  wire [7:0] t_r24_c1_2;
  wire [7:0] t_r24_c1_3;
  wire [7:0] t_r24_c1_4;
  wire [7:0] t_r24_c1_5;
  wire [7:0] t_r24_c1_6;
  wire [7:0] t_r24_c1_7;
  wire [7:0] t_r24_c1_8;
  wire [7:0] t_r24_c1_9;
  wire [7:0] t_r24_c1_10;
  wire [7:0] t_r24_c1_11;
  wire [7:0] t_r24_c1_12;
  wire [7:0] t_r24_c2_0;
  wire [7:0] t_r24_c2_1;
  wire [7:0] t_r24_c2_2;
  wire [7:0] t_r24_c2_3;
  wire [7:0] t_r24_c2_4;
  wire [7:0] t_r24_c2_5;
  wire [7:0] t_r24_c2_6;
  wire [7:0] t_r24_c2_7;
  wire [7:0] t_r24_c2_8;
  wire [7:0] t_r24_c2_9;
  wire [7:0] t_r24_c2_10;
  wire [7:0] t_r24_c2_11;
  wire [7:0] t_r24_c2_12;
  wire [7:0] t_r24_c3_0;
  wire [7:0] t_r24_c3_1;
  wire [7:0] t_r24_c3_2;
  wire [7:0] t_r24_c3_3;
  wire [7:0] t_r24_c3_4;
  wire [7:0] t_r24_c3_5;
  wire [7:0] t_r24_c3_6;
  wire [7:0] t_r24_c3_7;
  wire [7:0] t_r24_c3_8;
  wire [7:0] t_r24_c3_9;
  wire [7:0] t_r24_c3_10;
  wire [7:0] t_r24_c3_11;
  wire [7:0] t_r24_c3_12;
  wire [7:0] t_r24_c4_0;
  wire [7:0] t_r24_c4_1;
  wire [7:0] t_r24_c4_2;
  wire [7:0] t_r24_c4_3;
  wire [7:0] t_r24_c4_4;
  wire [7:0] t_r24_c4_5;
  wire [7:0] t_r24_c4_6;
  wire [7:0] t_r24_c4_7;
  wire [7:0] t_r24_c4_8;
  wire [7:0] t_r24_c4_9;
  wire [7:0] t_r24_c4_10;
  wire [7:0] t_r24_c4_11;
  wire [7:0] t_r24_c4_12;
  wire [7:0] t_r24_c5_0;
  wire [7:0] t_r24_c5_1;
  wire [7:0] t_r24_c5_2;
  wire [7:0] t_r24_c5_3;
  wire [7:0] t_r24_c5_4;
  wire [7:0] t_r24_c5_5;
  wire [7:0] t_r24_c5_6;
  wire [7:0] t_r24_c5_7;
  wire [7:0] t_r24_c5_8;
  wire [7:0] t_r24_c5_9;
  wire [7:0] t_r24_c5_10;
  wire [7:0] t_r24_c5_11;
  wire [7:0] t_r24_c5_12;
  wire [7:0] t_r24_c6_0;
  wire [7:0] t_r24_c6_1;
  wire [7:0] t_r24_c6_2;
  wire [7:0] t_r24_c6_3;
  wire [7:0] t_r24_c6_4;
  wire [7:0] t_r24_c6_5;
  wire [7:0] t_r24_c6_6;
  wire [7:0] t_r24_c6_7;
  wire [7:0] t_r24_c6_8;
  wire [7:0] t_r24_c6_9;
  wire [7:0] t_r24_c6_10;
  wire [7:0] t_r24_c6_11;
  wire [7:0] t_r24_c6_12;
  wire [7:0] t_r24_c7_0;
  wire [7:0] t_r24_c7_1;
  wire [7:0] t_r24_c7_2;
  wire [7:0] t_r24_c7_3;
  wire [7:0] t_r24_c7_4;
  wire [7:0] t_r24_c7_5;
  wire [7:0] t_r24_c7_6;
  wire [7:0] t_r24_c7_7;
  wire [7:0] t_r24_c7_8;
  wire [7:0] t_r24_c7_9;
  wire [7:0] t_r24_c7_10;
  wire [7:0] t_r24_c7_11;
  wire [7:0] t_r24_c7_12;
  wire [7:0] t_r24_c8_0;
  wire [7:0] t_r24_c8_1;
  wire [7:0] t_r24_c8_2;
  wire [7:0] t_r24_c8_3;
  wire [7:0] t_r24_c8_4;
  wire [7:0] t_r24_c8_5;
  wire [7:0] t_r24_c8_6;
  wire [7:0] t_r24_c8_7;
  wire [7:0] t_r24_c8_8;
  wire [7:0] t_r24_c8_9;
  wire [7:0] t_r24_c8_10;
  wire [7:0] t_r24_c8_11;
  wire [7:0] t_r24_c8_12;
  wire [7:0] t_r24_c9_0;
  wire [7:0] t_r24_c9_1;
  wire [7:0] t_r24_c9_2;
  wire [7:0] t_r24_c9_3;
  wire [7:0] t_r24_c9_4;
  wire [7:0] t_r24_c9_5;
  wire [7:0] t_r24_c9_6;
  wire [7:0] t_r24_c9_7;
  wire [7:0] t_r24_c9_8;
  wire [7:0] t_r24_c9_9;
  wire [7:0] t_r24_c9_10;
  wire [7:0] t_r24_c9_11;
  wire [7:0] t_r24_c9_12;
  wire [7:0] t_r24_c10_0;
  wire [7:0] t_r24_c10_1;
  wire [7:0] t_r24_c10_2;
  wire [7:0] t_r24_c10_3;
  wire [7:0] t_r24_c10_4;
  wire [7:0] t_r24_c10_5;
  wire [7:0] t_r24_c10_6;
  wire [7:0] t_r24_c10_7;
  wire [7:0] t_r24_c10_8;
  wire [7:0] t_r24_c10_9;
  wire [7:0] t_r24_c10_10;
  wire [7:0] t_r24_c10_11;
  wire [7:0] t_r24_c10_12;
  wire [7:0] t_r24_c11_0;
  wire [7:0] t_r24_c11_1;
  wire [7:0] t_r24_c11_2;
  wire [7:0] t_r24_c11_3;
  wire [7:0] t_r24_c11_4;
  wire [7:0] t_r24_c11_5;
  wire [7:0] t_r24_c11_6;
  wire [7:0] t_r24_c11_7;
  wire [7:0] t_r24_c11_8;
  wire [7:0] t_r24_c11_9;
  wire [7:0] t_r24_c11_10;
  wire [7:0] t_r24_c11_11;
  wire [7:0] t_r24_c11_12;
  wire [7:0] t_r24_c12_0;
  wire [7:0] t_r24_c12_1;
  wire [7:0] t_r24_c12_2;
  wire [7:0] t_r24_c12_3;
  wire [7:0] t_r24_c12_4;
  wire [7:0] t_r24_c12_5;
  wire [7:0] t_r24_c12_6;
  wire [7:0] t_r24_c12_7;
  wire [7:0] t_r24_c12_8;
  wire [7:0] t_r24_c12_9;
  wire [7:0] t_r24_c12_10;
  wire [7:0] t_r24_c12_11;
  wire [7:0] t_r24_c12_12;
  wire [7:0] t_r24_c13_0;
  wire [7:0] t_r24_c13_1;
  wire [7:0] t_r24_c13_2;
  wire [7:0] t_r24_c13_3;
  wire [7:0] t_r24_c13_4;
  wire [7:0] t_r24_c13_5;
  wire [7:0] t_r24_c13_6;
  wire [7:0] t_r24_c13_7;
  wire [7:0] t_r24_c13_8;
  wire [7:0] t_r24_c13_9;
  wire [7:0] t_r24_c13_10;
  wire [7:0] t_r24_c13_11;
  wire [7:0] t_r24_c13_12;
  wire [7:0] t_r24_c14_0;
  wire [7:0] t_r24_c14_1;
  wire [7:0] t_r24_c14_2;
  wire [7:0] t_r24_c14_3;
  wire [7:0] t_r24_c14_4;
  wire [7:0] t_r24_c14_5;
  wire [7:0] t_r24_c14_6;
  wire [7:0] t_r24_c14_7;
  wire [7:0] t_r24_c14_8;
  wire [7:0] t_r24_c14_9;
  wire [7:0] t_r24_c14_10;
  wire [7:0] t_r24_c14_11;
  wire [7:0] t_r24_c14_12;
  wire [7:0] t_r24_c15_0;
  wire [7:0] t_r24_c15_1;
  wire [7:0] t_r24_c15_2;
  wire [7:0] t_r24_c15_3;
  wire [7:0] t_r24_c15_4;
  wire [7:0] t_r24_c15_5;
  wire [7:0] t_r24_c15_6;
  wire [7:0] t_r24_c15_7;
  wire [7:0] t_r24_c15_8;
  wire [7:0] t_r24_c15_9;
  wire [7:0] t_r24_c15_10;
  wire [7:0] t_r24_c15_11;
  wire [7:0] t_r24_c15_12;
  wire [7:0] t_r24_c16_0;
  wire [7:0] t_r24_c16_1;
  wire [7:0] t_r24_c16_2;
  wire [7:0] t_r24_c16_3;
  wire [7:0] t_r24_c16_4;
  wire [7:0] t_r24_c16_5;
  wire [7:0] t_r24_c16_6;
  wire [7:0] t_r24_c16_7;
  wire [7:0] t_r24_c16_8;
  wire [7:0] t_r24_c16_9;
  wire [7:0] t_r24_c16_10;
  wire [7:0] t_r24_c16_11;
  wire [7:0] t_r24_c16_12;
  wire [7:0] t_r24_c17_0;
  wire [7:0] t_r24_c17_1;
  wire [7:0] t_r24_c17_2;
  wire [7:0] t_r24_c17_3;
  wire [7:0] t_r24_c17_4;
  wire [7:0] t_r24_c17_5;
  wire [7:0] t_r24_c17_6;
  wire [7:0] t_r24_c17_7;
  wire [7:0] t_r24_c17_8;
  wire [7:0] t_r24_c17_9;
  wire [7:0] t_r24_c17_10;
  wire [7:0] t_r24_c17_11;
  wire [7:0] t_r24_c17_12;
  wire [7:0] t_r24_c18_0;
  wire [7:0] t_r24_c18_1;
  wire [7:0] t_r24_c18_2;
  wire [7:0] t_r24_c18_3;
  wire [7:0] t_r24_c18_4;
  wire [7:0] t_r24_c18_5;
  wire [7:0] t_r24_c18_6;
  wire [7:0] t_r24_c18_7;
  wire [7:0] t_r24_c18_8;
  wire [7:0] t_r24_c18_9;
  wire [7:0] t_r24_c18_10;
  wire [7:0] t_r24_c18_11;
  wire [7:0] t_r24_c18_12;
  wire [7:0] t_r24_c19_0;
  wire [7:0] t_r24_c19_1;
  wire [7:0] t_r24_c19_2;
  wire [7:0] t_r24_c19_3;
  wire [7:0] t_r24_c19_4;
  wire [7:0] t_r24_c19_5;
  wire [7:0] t_r24_c19_6;
  wire [7:0] t_r24_c19_7;
  wire [7:0] t_r24_c19_8;
  wire [7:0] t_r24_c19_9;
  wire [7:0] t_r24_c19_10;
  wire [7:0] t_r24_c19_11;
  wire [7:0] t_r24_c19_12;
  wire [7:0] t_r24_c20_0;
  wire [7:0] t_r24_c20_1;
  wire [7:0] t_r24_c20_2;
  wire [7:0] t_r24_c20_3;
  wire [7:0] t_r24_c20_4;
  wire [7:0] t_r24_c20_5;
  wire [7:0] t_r24_c20_6;
  wire [7:0] t_r24_c20_7;
  wire [7:0] t_r24_c20_8;
  wire [7:0] t_r24_c20_9;
  wire [7:0] t_r24_c20_10;
  wire [7:0] t_r24_c20_11;
  wire [7:0] t_r24_c20_12;
  wire [7:0] t_r24_c21_0;
  wire [7:0] t_r24_c21_1;
  wire [7:0] t_r24_c21_2;
  wire [7:0] t_r24_c21_3;
  wire [7:0] t_r24_c21_4;
  wire [7:0] t_r24_c21_5;
  wire [7:0] t_r24_c21_6;
  wire [7:0] t_r24_c21_7;
  wire [7:0] t_r24_c21_8;
  wire [7:0] t_r24_c21_9;
  wire [7:0] t_r24_c21_10;
  wire [7:0] t_r24_c21_11;
  wire [7:0] t_r24_c21_12;
  wire [7:0] t_r24_c22_0;
  wire [7:0] t_r24_c22_1;
  wire [7:0] t_r24_c22_2;
  wire [7:0] t_r24_c22_3;
  wire [7:0] t_r24_c22_4;
  wire [7:0] t_r24_c22_5;
  wire [7:0] t_r24_c22_6;
  wire [7:0] t_r24_c22_7;
  wire [7:0] t_r24_c22_8;
  wire [7:0] t_r24_c22_9;
  wire [7:0] t_r24_c22_10;
  wire [7:0] t_r24_c22_11;
  wire [7:0] t_r24_c22_12;
  wire [7:0] t_r24_c23_0;
  wire [7:0] t_r24_c23_1;
  wire [7:0] t_r24_c23_2;
  wire [7:0] t_r24_c23_3;
  wire [7:0] t_r24_c23_4;
  wire [7:0] t_r24_c23_5;
  wire [7:0] t_r24_c23_6;
  wire [7:0] t_r24_c23_7;
  wire [7:0] t_r24_c23_8;
  wire [7:0] t_r24_c23_9;
  wire [7:0] t_r24_c23_10;
  wire [7:0] t_r24_c23_11;
  wire [7:0] t_r24_c23_12;
  wire [7:0] t_r24_c24_0;
  wire [7:0] t_r24_c24_1;
  wire [7:0] t_r24_c24_2;
  wire [7:0] t_r24_c24_3;
  wire [7:0] t_r24_c24_4;
  wire [7:0] t_r24_c24_5;
  wire [7:0] t_r24_c24_6;
  wire [7:0] t_r24_c24_7;
  wire [7:0] t_r24_c24_8;
  wire [7:0] t_r24_c24_9;
  wire [7:0] t_r24_c24_10;
  wire [7:0] t_r24_c24_11;
  wire [7:0] t_r24_c24_12;
  wire [7:0] t_r24_c25_0;
  wire [7:0] t_r24_c25_1;
  wire [7:0] t_r24_c25_2;
  wire [7:0] t_r24_c25_3;
  wire [7:0] t_r24_c25_4;
  wire [7:0] t_r24_c25_5;
  wire [7:0] t_r24_c25_6;
  wire [7:0] t_r24_c25_7;
  wire [7:0] t_r24_c25_8;
  wire [7:0] t_r24_c25_9;
  wire [7:0] t_r24_c25_10;
  wire [7:0] t_r24_c25_11;
  wire [7:0] t_r24_c25_12;
  wire [7:0] t_r24_c26_0;
  wire [7:0] t_r24_c26_1;
  wire [7:0] t_r24_c26_2;
  wire [7:0] t_r24_c26_3;
  wire [7:0] t_r24_c26_4;
  wire [7:0] t_r24_c26_5;
  wire [7:0] t_r24_c26_6;
  wire [7:0] t_r24_c26_7;
  wire [7:0] t_r24_c26_8;
  wire [7:0] t_r24_c26_9;
  wire [7:0] t_r24_c26_10;
  wire [7:0] t_r24_c26_11;
  wire [7:0] t_r24_c26_12;
  wire [7:0] t_r24_c27_0;
  wire [7:0] t_r24_c27_1;
  wire [7:0] t_r24_c27_2;
  wire [7:0] t_r24_c27_3;
  wire [7:0] t_r24_c27_4;
  wire [7:0] t_r24_c27_5;
  wire [7:0] t_r24_c27_6;
  wire [7:0] t_r24_c27_7;
  wire [7:0] t_r24_c27_8;
  wire [7:0] t_r24_c27_9;
  wire [7:0] t_r24_c27_10;
  wire [7:0] t_r24_c27_11;
  wire [7:0] t_r24_c27_12;
  wire [7:0] t_r24_c28_0;
  wire [7:0] t_r24_c28_1;
  wire [7:0] t_r24_c28_2;
  wire [7:0] t_r24_c28_3;
  wire [7:0] t_r24_c28_4;
  wire [7:0] t_r24_c28_5;
  wire [7:0] t_r24_c28_6;
  wire [7:0] t_r24_c28_7;
  wire [7:0] t_r24_c28_8;
  wire [7:0] t_r24_c28_9;
  wire [7:0] t_r24_c28_10;
  wire [7:0] t_r24_c28_11;
  wire [7:0] t_r24_c28_12;
  wire [7:0] t_r24_c29_0;
  wire [7:0] t_r24_c29_1;
  wire [7:0] t_r24_c29_2;
  wire [7:0] t_r24_c29_3;
  wire [7:0] t_r24_c29_4;
  wire [7:0] t_r24_c29_5;
  wire [7:0] t_r24_c29_6;
  wire [7:0] t_r24_c29_7;
  wire [7:0] t_r24_c29_8;
  wire [7:0] t_r24_c29_9;
  wire [7:0] t_r24_c29_10;
  wire [7:0] t_r24_c29_11;
  wire [7:0] t_r24_c29_12;
  wire [7:0] t_r24_c30_0;
  wire [7:0] t_r24_c30_1;
  wire [7:0] t_r24_c30_2;
  wire [7:0] t_r24_c30_3;
  wire [7:0] t_r24_c30_4;
  wire [7:0] t_r24_c30_5;
  wire [7:0] t_r24_c30_6;
  wire [7:0] t_r24_c30_7;
  wire [7:0] t_r24_c30_8;
  wire [7:0] t_r24_c30_9;
  wire [7:0] t_r24_c30_10;
  wire [7:0] t_r24_c30_11;
  wire [7:0] t_r24_c30_12;
  wire [7:0] t_r24_c31_0;
  wire [7:0] t_r24_c31_1;
  wire [7:0] t_r24_c31_2;
  wire [7:0] t_r24_c31_3;
  wire [7:0] t_r24_c31_4;
  wire [7:0] t_r24_c31_5;
  wire [7:0] t_r24_c31_6;
  wire [7:0] t_r24_c31_7;
  wire [7:0] t_r24_c31_8;
  wire [7:0] t_r24_c31_9;
  wire [7:0] t_r24_c31_10;
  wire [7:0] t_r24_c31_11;
  wire [7:0] t_r24_c31_12;
  wire [7:0] t_r24_c32_0;
  wire [7:0] t_r24_c32_1;
  wire [7:0] t_r24_c32_2;
  wire [7:0] t_r24_c32_3;
  wire [7:0] t_r24_c32_4;
  wire [7:0] t_r24_c32_5;
  wire [7:0] t_r24_c32_6;
  wire [7:0] t_r24_c32_7;
  wire [7:0] t_r24_c32_8;
  wire [7:0] t_r24_c32_9;
  wire [7:0] t_r24_c32_10;
  wire [7:0] t_r24_c32_11;
  wire [7:0] t_r24_c32_12;
  wire [7:0] t_r24_c33_0;
  wire [7:0] t_r24_c33_1;
  wire [7:0] t_r24_c33_2;
  wire [7:0] t_r24_c33_3;
  wire [7:0] t_r24_c33_4;
  wire [7:0] t_r24_c33_5;
  wire [7:0] t_r24_c33_6;
  wire [7:0] t_r24_c33_7;
  wire [7:0] t_r24_c33_8;
  wire [7:0] t_r24_c33_9;
  wire [7:0] t_r24_c33_10;
  wire [7:0] t_r24_c33_11;
  wire [7:0] t_r24_c33_12;
  wire [7:0] t_r24_c34_0;
  wire [7:0] t_r24_c34_1;
  wire [7:0] t_r24_c34_2;
  wire [7:0] t_r24_c34_3;
  wire [7:0] t_r24_c34_4;
  wire [7:0] t_r24_c34_5;
  wire [7:0] t_r24_c34_6;
  wire [7:0] t_r24_c34_7;
  wire [7:0] t_r24_c34_8;
  wire [7:0] t_r24_c34_9;
  wire [7:0] t_r24_c34_10;
  wire [7:0] t_r24_c34_11;
  wire [7:0] t_r24_c34_12;
  wire [7:0] t_r24_c35_0;
  wire [7:0] t_r24_c35_1;
  wire [7:0] t_r24_c35_2;
  wire [7:0] t_r24_c35_3;
  wire [7:0] t_r24_c35_4;
  wire [7:0] t_r24_c35_5;
  wire [7:0] t_r24_c35_6;
  wire [7:0] t_r24_c35_7;
  wire [7:0] t_r24_c35_8;
  wire [7:0] t_r24_c35_9;
  wire [7:0] t_r24_c35_10;
  wire [7:0] t_r24_c35_11;
  wire [7:0] t_r24_c35_12;
  wire [7:0] t_r24_c36_0;
  wire [7:0] t_r24_c36_1;
  wire [7:0] t_r24_c36_2;
  wire [7:0] t_r24_c36_3;
  wire [7:0] t_r24_c36_4;
  wire [7:0] t_r24_c36_5;
  wire [7:0] t_r24_c36_6;
  wire [7:0] t_r24_c36_7;
  wire [7:0] t_r24_c36_8;
  wire [7:0] t_r24_c36_9;
  wire [7:0] t_r24_c36_10;
  wire [7:0] t_r24_c36_11;
  wire [7:0] t_r24_c36_12;
  wire [7:0] t_r24_c37_0;
  wire [7:0] t_r24_c37_1;
  wire [7:0] t_r24_c37_2;
  wire [7:0] t_r24_c37_3;
  wire [7:0] t_r24_c37_4;
  wire [7:0] t_r24_c37_5;
  wire [7:0] t_r24_c37_6;
  wire [7:0] t_r24_c37_7;
  wire [7:0] t_r24_c37_8;
  wire [7:0] t_r24_c37_9;
  wire [7:0] t_r24_c37_10;
  wire [7:0] t_r24_c37_11;
  wire [7:0] t_r24_c37_12;
  wire [7:0] t_r24_c38_0;
  wire [7:0] t_r24_c38_1;
  wire [7:0] t_r24_c38_2;
  wire [7:0] t_r24_c38_3;
  wire [7:0] t_r24_c38_4;
  wire [7:0] t_r24_c38_5;
  wire [7:0] t_r24_c38_6;
  wire [7:0] t_r24_c38_7;
  wire [7:0] t_r24_c38_8;
  wire [7:0] t_r24_c38_9;
  wire [7:0] t_r24_c38_10;
  wire [7:0] t_r24_c38_11;
  wire [7:0] t_r24_c38_12;
  wire [7:0] t_r24_c39_0;
  wire [7:0] t_r24_c39_1;
  wire [7:0] t_r24_c39_2;
  wire [7:0] t_r24_c39_3;
  wire [7:0] t_r24_c39_4;
  wire [7:0] t_r24_c39_5;
  wire [7:0] t_r24_c39_6;
  wire [7:0] t_r24_c39_7;
  wire [7:0] t_r24_c39_8;
  wire [7:0] t_r24_c39_9;
  wire [7:0] t_r24_c39_10;
  wire [7:0] t_r24_c39_11;
  wire [7:0] t_r24_c39_12;
  wire [7:0] t_r24_c40_0;
  wire [7:0] t_r24_c40_1;
  wire [7:0] t_r24_c40_2;
  wire [7:0] t_r24_c40_3;
  wire [7:0] t_r24_c40_4;
  wire [7:0] t_r24_c40_5;
  wire [7:0] t_r24_c40_6;
  wire [7:0] t_r24_c40_7;
  wire [7:0] t_r24_c40_8;
  wire [7:0] t_r24_c40_9;
  wire [7:0] t_r24_c40_10;
  wire [7:0] t_r24_c40_11;
  wire [7:0] t_r24_c40_12;
  wire [7:0] t_r24_c41_0;
  wire [7:0] t_r24_c41_1;
  wire [7:0] t_r24_c41_2;
  wire [7:0] t_r24_c41_3;
  wire [7:0] t_r24_c41_4;
  wire [7:0] t_r24_c41_5;
  wire [7:0] t_r24_c41_6;
  wire [7:0] t_r24_c41_7;
  wire [7:0] t_r24_c41_8;
  wire [7:0] t_r24_c41_9;
  wire [7:0] t_r24_c41_10;
  wire [7:0] t_r24_c41_11;
  wire [7:0] t_r24_c41_12;
  wire [7:0] t_r24_c42_0;
  wire [7:0] t_r24_c42_1;
  wire [7:0] t_r24_c42_2;
  wire [7:0] t_r24_c42_3;
  wire [7:0] t_r24_c42_4;
  wire [7:0] t_r24_c42_5;
  wire [7:0] t_r24_c42_6;
  wire [7:0] t_r24_c42_7;
  wire [7:0] t_r24_c42_8;
  wire [7:0] t_r24_c42_9;
  wire [7:0] t_r24_c42_10;
  wire [7:0] t_r24_c42_11;
  wire [7:0] t_r24_c42_12;
  wire [7:0] t_r24_c43_0;
  wire [7:0] t_r24_c43_1;
  wire [7:0] t_r24_c43_2;
  wire [7:0] t_r24_c43_3;
  wire [7:0] t_r24_c43_4;
  wire [7:0] t_r24_c43_5;
  wire [7:0] t_r24_c43_6;
  wire [7:0] t_r24_c43_7;
  wire [7:0] t_r24_c43_8;
  wire [7:0] t_r24_c43_9;
  wire [7:0] t_r24_c43_10;
  wire [7:0] t_r24_c43_11;
  wire [7:0] t_r24_c43_12;
  wire [7:0] t_r24_c44_0;
  wire [7:0] t_r24_c44_1;
  wire [7:0] t_r24_c44_2;
  wire [7:0] t_r24_c44_3;
  wire [7:0] t_r24_c44_4;
  wire [7:0] t_r24_c44_5;
  wire [7:0] t_r24_c44_6;
  wire [7:0] t_r24_c44_7;
  wire [7:0] t_r24_c44_8;
  wire [7:0] t_r24_c44_9;
  wire [7:0] t_r24_c44_10;
  wire [7:0] t_r24_c44_11;
  wire [7:0] t_r24_c44_12;
  wire [7:0] t_r24_c45_0;
  wire [7:0] t_r24_c45_1;
  wire [7:0] t_r24_c45_2;
  wire [7:0] t_r24_c45_3;
  wire [7:0] t_r24_c45_4;
  wire [7:0] t_r24_c45_5;
  wire [7:0] t_r24_c45_6;
  wire [7:0] t_r24_c45_7;
  wire [7:0] t_r24_c45_8;
  wire [7:0] t_r24_c45_9;
  wire [7:0] t_r24_c45_10;
  wire [7:0] t_r24_c45_11;
  wire [7:0] t_r24_c45_12;
  wire [7:0] t_r24_c46_0;
  wire [7:0] t_r24_c46_1;
  wire [7:0] t_r24_c46_2;
  wire [7:0] t_r24_c46_3;
  wire [7:0] t_r24_c46_4;
  wire [7:0] t_r24_c46_5;
  wire [7:0] t_r24_c46_6;
  wire [7:0] t_r24_c46_7;
  wire [7:0] t_r24_c46_8;
  wire [7:0] t_r24_c46_9;
  wire [7:0] t_r24_c46_10;
  wire [7:0] t_r24_c46_11;
  wire [7:0] t_r24_c46_12;
  wire [7:0] t_r24_c47_0;
  wire [7:0] t_r24_c47_1;
  wire [7:0] t_r24_c47_2;
  wire [7:0] t_r24_c47_3;
  wire [7:0] t_r24_c47_4;
  wire [7:0] t_r24_c47_5;
  wire [7:0] t_r24_c47_6;
  wire [7:0] t_r24_c47_7;
  wire [7:0] t_r24_c47_8;
  wire [7:0] t_r24_c47_9;
  wire [7:0] t_r24_c47_10;
  wire [7:0] t_r24_c47_11;
  wire [7:0] t_r24_c47_12;
  wire [7:0] t_r24_c48_0;
  wire [7:0] t_r24_c48_1;
  wire [7:0] t_r24_c48_2;
  wire [7:0] t_r24_c48_3;
  wire [7:0] t_r24_c48_4;
  wire [7:0] t_r24_c48_5;
  wire [7:0] t_r24_c48_6;
  wire [7:0] t_r24_c48_7;
  wire [7:0] t_r24_c48_8;
  wire [7:0] t_r24_c48_9;
  wire [7:0] t_r24_c48_10;
  wire [7:0] t_r24_c48_11;
  wire [7:0] t_r24_c48_12;
  wire [7:0] t_r24_c49_0;
  wire [7:0] t_r24_c49_1;
  wire [7:0] t_r24_c49_2;
  wire [7:0] t_r24_c49_3;
  wire [7:0] t_r24_c49_4;
  wire [7:0] t_r24_c49_5;
  wire [7:0] t_r24_c49_6;
  wire [7:0] t_r24_c49_7;
  wire [7:0] t_r24_c49_8;
  wire [7:0] t_r24_c49_9;
  wire [7:0] t_r24_c49_10;
  wire [7:0] t_r24_c49_11;
  wire [7:0] t_r24_c49_12;
  wire [7:0] t_r24_c50_0;
  wire [7:0] t_r24_c50_1;
  wire [7:0] t_r24_c50_2;
  wire [7:0] t_r24_c50_3;
  wire [7:0] t_r24_c50_4;
  wire [7:0] t_r24_c50_5;
  wire [7:0] t_r24_c50_6;
  wire [7:0] t_r24_c50_7;
  wire [7:0] t_r24_c50_8;
  wire [7:0] t_r24_c50_9;
  wire [7:0] t_r24_c50_10;
  wire [7:0] t_r24_c50_11;
  wire [7:0] t_r24_c50_12;
  wire [7:0] t_r24_c51_0;
  wire [7:0] t_r24_c51_1;
  wire [7:0] t_r24_c51_2;
  wire [7:0] t_r24_c51_3;
  wire [7:0] t_r24_c51_4;
  wire [7:0] t_r24_c51_5;
  wire [7:0] t_r24_c51_6;
  wire [7:0] t_r24_c51_7;
  wire [7:0] t_r24_c51_8;
  wire [7:0] t_r24_c51_9;
  wire [7:0] t_r24_c51_10;
  wire [7:0] t_r24_c51_11;
  wire [7:0] t_r24_c51_12;
  wire [7:0] t_r24_c52_0;
  wire [7:0] t_r24_c52_1;
  wire [7:0] t_r24_c52_2;
  wire [7:0] t_r24_c52_3;
  wire [7:0] t_r24_c52_4;
  wire [7:0] t_r24_c52_5;
  wire [7:0] t_r24_c52_6;
  wire [7:0] t_r24_c52_7;
  wire [7:0] t_r24_c52_8;
  wire [7:0] t_r24_c52_9;
  wire [7:0] t_r24_c52_10;
  wire [7:0] t_r24_c52_11;
  wire [7:0] t_r24_c52_12;
  wire [7:0] t_r24_c53_0;
  wire [7:0] t_r24_c53_1;
  wire [7:0] t_r24_c53_2;
  wire [7:0] t_r24_c53_3;
  wire [7:0] t_r24_c53_4;
  wire [7:0] t_r24_c53_5;
  wire [7:0] t_r24_c53_6;
  wire [7:0] t_r24_c53_7;
  wire [7:0] t_r24_c53_8;
  wire [7:0] t_r24_c53_9;
  wire [7:0] t_r24_c53_10;
  wire [7:0] t_r24_c53_11;
  wire [7:0] t_r24_c53_12;
  wire [7:0] t_r24_c54_0;
  wire [7:0] t_r24_c54_1;
  wire [7:0] t_r24_c54_2;
  wire [7:0] t_r24_c54_3;
  wire [7:0] t_r24_c54_4;
  wire [7:0] t_r24_c54_5;
  wire [7:0] t_r24_c54_6;
  wire [7:0] t_r24_c54_7;
  wire [7:0] t_r24_c54_8;
  wire [7:0] t_r24_c54_9;
  wire [7:0] t_r24_c54_10;
  wire [7:0] t_r24_c54_11;
  wire [7:0] t_r24_c54_12;
  wire [7:0] t_r24_c55_0;
  wire [7:0] t_r24_c55_1;
  wire [7:0] t_r24_c55_2;
  wire [7:0] t_r24_c55_3;
  wire [7:0] t_r24_c55_4;
  wire [7:0] t_r24_c55_5;
  wire [7:0] t_r24_c55_6;
  wire [7:0] t_r24_c55_7;
  wire [7:0] t_r24_c55_8;
  wire [7:0] t_r24_c55_9;
  wire [7:0] t_r24_c55_10;
  wire [7:0] t_r24_c55_11;
  wire [7:0] t_r24_c55_12;
  wire [7:0] t_r24_c56_0;
  wire [7:0] t_r24_c56_1;
  wire [7:0] t_r24_c56_2;
  wire [7:0] t_r24_c56_3;
  wire [7:0] t_r24_c56_4;
  wire [7:0] t_r24_c56_5;
  wire [7:0] t_r24_c56_6;
  wire [7:0] t_r24_c56_7;
  wire [7:0] t_r24_c56_8;
  wire [7:0] t_r24_c56_9;
  wire [7:0] t_r24_c56_10;
  wire [7:0] t_r24_c56_11;
  wire [7:0] t_r24_c56_12;
  wire [7:0] t_r24_c57_0;
  wire [7:0] t_r24_c57_1;
  wire [7:0] t_r24_c57_2;
  wire [7:0] t_r24_c57_3;
  wire [7:0] t_r24_c57_4;
  wire [7:0] t_r24_c57_5;
  wire [7:0] t_r24_c57_6;
  wire [7:0] t_r24_c57_7;
  wire [7:0] t_r24_c57_8;
  wire [7:0] t_r24_c57_9;
  wire [7:0] t_r24_c57_10;
  wire [7:0] t_r24_c57_11;
  wire [7:0] t_r24_c57_12;
  wire [7:0] t_r24_c58_0;
  wire [7:0] t_r24_c58_1;
  wire [7:0] t_r24_c58_2;
  wire [7:0] t_r24_c58_3;
  wire [7:0] t_r24_c58_4;
  wire [7:0] t_r24_c58_5;
  wire [7:0] t_r24_c58_6;
  wire [7:0] t_r24_c58_7;
  wire [7:0] t_r24_c58_8;
  wire [7:0] t_r24_c58_9;
  wire [7:0] t_r24_c58_10;
  wire [7:0] t_r24_c58_11;
  wire [7:0] t_r24_c58_12;
  wire [7:0] t_r24_c59_0;
  wire [7:0] t_r24_c59_1;
  wire [7:0] t_r24_c59_2;
  wire [7:0] t_r24_c59_3;
  wire [7:0] t_r24_c59_4;
  wire [7:0] t_r24_c59_5;
  wire [7:0] t_r24_c59_6;
  wire [7:0] t_r24_c59_7;
  wire [7:0] t_r24_c59_8;
  wire [7:0] t_r24_c59_9;
  wire [7:0] t_r24_c59_10;
  wire [7:0] t_r24_c59_11;
  wire [7:0] t_r24_c59_12;
  wire [7:0] t_r24_c60_0;
  wire [7:0] t_r24_c60_1;
  wire [7:0] t_r24_c60_2;
  wire [7:0] t_r24_c60_3;
  wire [7:0] t_r24_c60_4;
  wire [7:0] t_r24_c60_5;
  wire [7:0] t_r24_c60_6;
  wire [7:0] t_r24_c60_7;
  wire [7:0] t_r24_c60_8;
  wire [7:0] t_r24_c60_9;
  wire [7:0] t_r24_c60_10;
  wire [7:0] t_r24_c60_11;
  wire [7:0] t_r24_c60_12;
  wire [7:0] t_r24_c61_0;
  wire [7:0] t_r24_c61_1;
  wire [7:0] t_r24_c61_2;
  wire [7:0] t_r24_c61_3;
  wire [7:0] t_r24_c61_4;
  wire [7:0] t_r24_c61_5;
  wire [7:0] t_r24_c61_6;
  wire [7:0] t_r24_c61_7;
  wire [7:0] t_r24_c61_8;
  wire [7:0] t_r24_c61_9;
  wire [7:0] t_r24_c61_10;
  wire [7:0] t_r24_c61_11;
  wire [7:0] t_r24_c61_12;
  wire [7:0] t_r24_c62_0;
  wire [7:0] t_r24_c62_1;
  wire [7:0] t_r24_c62_2;
  wire [7:0] t_r24_c62_3;
  wire [7:0] t_r24_c62_4;
  wire [7:0] t_r24_c62_5;
  wire [7:0] t_r24_c62_6;
  wire [7:0] t_r24_c62_7;
  wire [7:0] t_r24_c62_8;
  wire [7:0] t_r24_c62_9;
  wire [7:0] t_r24_c62_10;
  wire [7:0] t_r24_c62_11;
  wire [7:0] t_r24_c62_12;
  wire [7:0] t_r24_c63_0;
  wire [7:0] t_r24_c63_1;
  wire [7:0] t_r24_c63_2;
  wire [7:0] t_r24_c63_3;
  wire [7:0] t_r24_c63_4;
  wire [7:0] t_r24_c63_5;
  wire [7:0] t_r24_c63_6;
  wire [7:0] t_r24_c63_7;
  wire [7:0] t_r24_c63_8;
  wire [7:0] t_r24_c63_9;
  wire [7:0] t_r24_c63_10;
  wire [7:0] t_r24_c63_11;
  wire [7:0] t_r24_c63_12;
  wire [7:0] t_r24_c64_0;
  wire [7:0] t_r24_c64_1;
  wire [7:0] t_r24_c64_2;
  wire [7:0] t_r24_c64_3;
  wire [7:0] t_r24_c64_4;
  wire [7:0] t_r24_c64_5;
  wire [7:0] t_r24_c64_6;
  wire [7:0] t_r24_c64_7;
  wire [7:0] t_r24_c64_8;
  wire [7:0] t_r24_c64_9;
  wire [7:0] t_r24_c64_10;
  wire [7:0] t_r24_c64_11;
  wire [7:0] t_r24_c64_12;
  wire [7:0] t_r24_c65_0;
  wire [7:0] t_r24_c65_1;
  wire [7:0] t_r24_c65_2;
  wire [7:0] t_r24_c65_3;
  wire [7:0] t_r24_c65_4;
  wire [7:0] t_r24_c65_5;
  wire [7:0] t_r24_c65_6;
  wire [7:0] t_r24_c65_7;
  wire [7:0] t_r24_c65_8;
  wire [7:0] t_r24_c65_9;
  wire [7:0] t_r24_c65_10;
  wire [7:0] t_r24_c65_11;
  wire [7:0] t_r24_c65_12;
  wire [7:0] t_r25_c0_0;
  wire [7:0] t_r25_c0_1;
  wire [7:0] t_r25_c0_2;
  wire [7:0] t_r25_c0_3;
  wire [7:0] t_r25_c0_4;
  wire [7:0] t_r25_c0_5;
  wire [7:0] t_r25_c0_6;
  wire [7:0] t_r25_c0_7;
  wire [7:0] t_r25_c0_8;
  wire [7:0] t_r25_c0_9;
  wire [7:0] t_r25_c0_10;
  wire [7:0] t_r25_c0_11;
  wire [7:0] t_r25_c0_12;
  wire [7:0] t_r25_c1_0;
  wire [7:0] t_r25_c1_1;
  wire [7:0] t_r25_c1_2;
  wire [7:0] t_r25_c1_3;
  wire [7:0] t_r25_c1_4;
  wire [7:0] t_r25_c1_5;
  wire [7:0] t_r25_c1_6;
  wire [7:0] t_r25_c1_7;
  wire [7:0] t_r25_c1_8;
  wire [7:0] t_r25_c1_9;
  wire [7:0] t_r25_c1_10;
  wire [7:0] t_r25_c1_11;
  wire [7:0] t_r25_c1_12;
  wire [7:0] t_r25_c2_0;
  wire [7:0] t_r25_c2_1;
  wire [7:0] t_r25_c2_2;
  wire [7:0] t_r25_c2_3;
  wire [7:0] t_r25_c2_4;
  wire [7:0] t_r25_c2_5;
  wire [7:0] t_r25_c2_6;
  wire [7:0] t_r25_c2_7;
  wire [7:0] t_r25_c2_8;
  wire [7:0] t_r25_c2_9;
  wire [7:0] t_r25_c2_10;
  wire [7:0] t_r25_c2_11;
  wire [7:0] t_r25_c2_12;
  wire [7:0] t_r25_c3_0;
  wire [7:0] t_r25_c3_1;
  wire [7:0] t_r25_c3_2;
  wire [7:0] t_r25_c3_3;
  wire [7:0] t_r25_c3_4;
  wire [7:0] t_r25_c3_5;
  wire [7:0] t_r25_c3_6;
  wire [7:0] t_r25_c3_7;
  wire [7:0] t_r25_c3_8;
  wire [7:0] t_r25_c3_9;
  wire [7:0] t_r25_c3_10;
  wire [7:0] t_r25_c3_11;
  wire [7:0] t_r25_c3_12;
  wire [7:0] t_r25_c4_0;
  wire [7:0] t_r25_c4_1;
  wire [7:0] t_r25_c4_2;
  wire [7:0] t_r25_c4_3;
  wire [7:0] t_r25_c4_4;
  wire [7:0] t_r25_c4_5;
  wire [7:0] t_r25_c4_6;
  wire [7:0] t_r25_c4_7;
  wire [7:0] t_r25_c4_8;
  wire [7:0] t_r25_c4_9;
  wire [7:0] t_r25_c4_10;
  wire [7:0] t_r25_c4_11;
  wire [7:0] t_r25_c4_12;
  wire [7:0] t_r25_c5_0;
  wire [7:0] t_r25_c5_1;
  wire [7:0] t_r25_c5_2;
  wire [7:0] t_r25_c5_3;
  wire [7:0] t_r25_c5_4;
  wire [7:0] t_r25_c5_5;
  wire [7:0] t_r25_c5_6;
  wire [7:0] t_r25_c5_7;
  wire [7:0] t_r25_c5_8;
  wire [7:0] t_r25_c5_9;
  wire [7:0] t_r25_c5_10;
  wire [7:0] t_r25_c5_11;
  wire [7:0] t_r25_c5_12;
  wire [7:0] t_r25_c6_0;
  wire [7:0] t_r25_c6_1;
  wire [7:0] t_r25_c6_2;
  wire [7:0] t_r25_c6_3;
  wire [7:0] t_r25_c6_4;
  wire [7:0] t_r25_c6_5;
  wire [7:0] t_r25_c6_6;
  wire [7:0] t_r25_c6_7;
  wire [7:0] t_r25_c6_8;
  wire [7:0] t_r25_c6_9;
  wire [7:0] t_r25_c6_10;
  wire [7:0] t_r25_c6_11;
  wire [7:0] t_r25_c6_12;
  wire [7:0] t_r25_c7_0;
  wire [7:0] t_r25_c7_1;
  wire [7:0] t_r25_c7_2;
  wire [7:0] t_r25_c7_3;
  wire [7:0] t_r25_c7_4;
  wire [7:0] t_r25_c7_5;
  wire [7:0] t_r25_c7_6;
  wire [7:0] t_r25_c7_7;
  wire [7:0] t_r25_c7_8;
  wire [7:0] t_r25_c7_9;
  wire [7:0] t_r25_c7_10;
  wire [7:0] t_r25_c7_11;
  wire [7:0] t_r25_c7_12;
  wire [7:0] t_r25_c8_0;
  wire [7:0] t_r25_c8_1;
  wire [7:0] t_r25_c8_2;
  wire [7:0] t_r25_c8_3;
  wire [7:0] t_r25_c8_4;
  wire [7:0] t_r25_c8_5;
  wire [7:0] t_r25_c8_6;
  wire [7:0] t_r25_c8_7;
  wire [7:0] t_r25_c8_8;
  wire [7:0] t_r25_c8_9;
  wire [7:0] t_r25_c8_10;
  wire [7:0] t_r25_c8_11;
  wire [7:0] t_r25_c8_12;
  wire [7:0] t_r25_c9_0;
  wire [7:0] t_r25_c9_1;
  wire [7:0] t_r25_c9_2;
  wire [7:0] t_r25_c9_3;
  wire [7:0] t_r25_c9_4;
  wire [7:0] t_r25_c9_5;
  wire [7:0] t_r25_c9_6;
  wire [7:0] t_r25_c9_7;
  wire [7:0] t_r25_c9_8;
  wire [7:0] t_r25_c9_9;
  wire [7:0] t_r25_c9_10;
  wire [7:0] t_r25_c9_11;
  wire [7:0] t_r25_c9_12;
  wire [7:0] t_r25_c10_0;
  wire [7:0] t_r25_c10_1;
  wire [7:0] t_r25_c10_2;
  wire [7:0] t_r25_c10_3;
  wire [7:0] t_r25_c10_4;
  wire [7:0] t_r25_c10_5;
  wire [7:0] t_r25_c10_6;
  wire [7:0] t_r25_c10_7;
  wire [7:0] t_r25_c10_8;
  wire [7:0] t_r25_c10_9;
  wire [7:0] t_r25_c10_10;
  wire [7:0] t_r25_c10_11;
  wire [7:0] t_r25_c10_12;
  wire [7:0] t_r25_c11_0;
  wire [7:0] t_r25_c11_1;
  wire [7:0] t_r25_c11_2;
  wire [7:0] t_r25_c11_3;
  wire [7:0] t_r25_c11_4;
  wire [7:0] t_r25_c11_5;
  wire [7:0] t_r25_c11_6;
  wire [7:0] t_r25_c11_7;
  wire [7:0] t_r25_c11_8;
  wire [7:0] t_r25_c11_9;
  wire [7:0] t_r25_c11_10;
  wire [7:0] t_r25_c11_11;
  wire [7:0] t_r25_c11_12;
  wire [7:0] t_r25_c12_0;
  wire [7:0] t_r25_c12_1;
  wire [7:0] t_r25_c12_2;
  wire [7:0] t_r25_c12_3;
  wire [7:0] t_r25_c12_4;
  wire [7:0] t_r25_c12_5;
  wire [7:0] t_r25_c12_6;
  wire [7:0] t_r25_c12_7;
  wire [7:0] t_r25_c12_8;
  wire [7:0] t_r25_c12_9;
  wire [7:0] t_r25_c12_10;
  wire [7:0] t_r25_c12_11;
  wire [7:0] t_r25_c12_12;
  wire [7:0] t_r25_c13_0;
  wire [7:0] t_r25_c13_1;
  wire [7:0] t_r25_c13_2;
  wire [7:0] t_r25_c13_3;
  wire [7:0] t_r25_c13_4;
  wire [7:0] t_r25_c13_5;
  wire [7:0] t_r25_c13_6;
  wire [7:0] t_r25_c13_7;
  wire [7:0] t_r25_c13_8;
  wire [7:0] t_r25_c13_9;
  wire [7:0] t_r25_c13_10;
  wire [7:0] t_r25_c13_11;
  wire [7:0] t_r25_c13_12;
  wire [7:0] t_r25_c14_0;
  wire [7:0] t_r25_c14_1;
  wire [7:0] t_r25_c14_2;
  wire [7:0] t_r25_c14_3;
  wire [7:0] t_r25_c14_4;
  wire [7:0] t_r25_c14_5;
  wire [7:0] t_r25_c14_6;
  wire [7:0] t_r25_c14_7;
  wire [7:0] t_r25_c14_8;
  wire [7:0] t_r25_c14_9;
  wire [7:0] t_r25_c14_10;
  wire [7:0] t_r25_c14_11;
  wire [7:0] t_r25_c14_12;
  wire [7:0] t_r25_c15_0;
  wire [7:0] t_r25_c15_1;
  wire [7:0] t_r25_c15_2;
  wire [7:0] t_r25_c15_3;
  wire [7:0] t_r25_c15_4;
  wire [7:0] t_r25_c15_5;
  wire [7:0] t_r25_c15_6;
  wire [7:0] t_r25_c15_7;
  wire [7:0] t_r25_c15_8;
  wire [7:0] t_r25_c15_9;
  wire [7:0] t_r25_c15_10;
  wire [7:0] t_r25_c15_11;
  wire [7:0] t_r25_c15_12;
  wire [7:0] t_r25_c16_0;
  wire [7:0] t_r25_c16_1;
  wire [7:0] t_r25_c16_2;
  wire [7:0] t_r25_c16_3;
  wire [7:0] t_r25_c16_4;
  wire [7:0] t_r25_c16_5;
  wire [7:0] t_r25_c16_6;
  wire [7:0] t_r25_c16_7;
  wire [7:0] t_r25_c16_8;
  wire [7:0] t_r25_c16_9;
  wire [7:0] t_r25_c16_10;
  wire [7:0] t_r25_c16_11;
  wire [7:0] t_r25_c16_12;
  wire [7:0] t_r25_c17_0;
  wire [7:0] t_r25_c17_1;
  wire [7:0] t_r25_c17_2;
  wire [7:0] t_r25_c17_3;
  wire [7:0] t_r25_c17_4;
  wire [7:0] t_r25_c17_5;
  wire [7:0] t_r25_c17_6;
  wire [7:0] t_r25_c17_7;
  wire [7:0] t_r25_c17_8;
  wire [7:0] t_r25_c17_9;
  wire [7:0] t_r25_c17_10;
  wire [7:0] t_r25_c17_11;
  wire [7:0] t_r25_c17_12;
  wire [7:0] t_r25_c18_0;
  wire [7:0] t_r25_c18_1;
  wire [7:0] t_r25_c18_2;
  wire [7:0] t_r25_c18_3;
  wire [7:0] t_r25_c18_4;
  wire [7:0] t_r25_c18_5;
  wire [7:0] t_r25_c18_6;
  wire [7:0] t_r25_c18_7;
  wire [7:0] t_r25_c18_8;
  wire [7:0] t_r25_c18_9;
  wire [7:0] t_r25_c18_10;
  wire [7:0] t_r25_c18_11;
  wire [7:0] t_r25_c18_12;
  wire [7:0] t_r25_c19_0;
  wire [7:0] t_r25_c19_1;
  wire [7:0] t_r25_c19_2;
  wire [7:0] t_r25_c19_3;
  wire [7:0] t_r25_c19_4;
  wire [7:0] t_r25_c19_5;
  wire [7:0] t_r25_c19_6;
  wire [7:0] t_r25_c19_7;
  wire [7:0] t_r25_c19_8;
  wire [7:0] t_r25_c19_9;
  wire [7:0] t_r25_c19_10;
  wire [7:0] t_r25_c19_11;
  wire [7:0] t_r25_c19_12;
  wire [7:0] t_r25_c20_0;
  wire [7:0] t_r25_c20_1;
  wire [7:0] t_r25_c20_2;
  wire [7:0] t_r25_c20_3;
  wire [7:0] t_r25_c20_4;
  wire [7:0] t_r25_c20_5;
  wire [7:0] t_r25_c20_6;
  wire [7:0] t_r25_c20_7;
  wire [7:0] t_r25_c20_8;
  wire [7:0] t_r25_c20_9;
  wire [7:0] t_r25_c20_10;
  wire [7:0] t_r25_c20_11;
  wire [7:0] t_r25_c20_12;
  wire [7:0] t_r25_c21_0;
  wire [7:0] t_r25_c21_1;
  wire [7:0] t_r25_c21_2;
  wire [7:0] t_r25_c21_3;
  wire [7:0] t_r25_c21_4;
  wire [7:0] t_r25_c21_5;
  wire [7:0] t_r25_c21_6;
  wire [7:0] t_r25_c21_7;
  wire [7:0] t_r25_c21_8;
  wire [7:0] t_r25_c21_9;
  wire [7:0] t_r25_c21_10;
  wire [7:0] t_r25_c21_11;
  wire [7:0] t_r25_c21_12;
  wire [7:0] t_r25_c22_0;
  wire [7:0] t_r25_c22_1;
  wire [7:0] t_r25_c22_2;
  wire [7:0] t_r25_c22_3;
  wire [7:0] t_r25_c22_4;
  wire [7:0] t_r25_c22_5;
  wire [7:0] t_r25_c22_6;
  wire [7:0] t_r25_c22_7;
  wire [7:0] t_r25_c22_8;
  wire [7:0] t_r25_c22_9;
  wire [7:0] t_r25_c22_10;
  wire [7:0] t_r25_c22_11;
  wire [7:0] t_r25_c22_12;
  wire [7:0] t_r25_c23_0;
  wire [7:0] t_r25_c23_1;
  wire [7:0] t_r25_c23_2;
  wire [7:0] t_r25_c23_3;
  wire [7:0] t_r25_c23_4;
  wire [7:0] t_r25_c23_5;
  wire [7:0] t_r25_c23_6;
  wire [7:0] t_r25_c23_7;
  wire [7:0] t_r25_c23_8;
  wire [7:0] t_r25_c23_9;
  wire [7:0] t_r25_c23_10;
  wire [7:0] t_r25_c23_11;
  wire [7:0] t_r25_c23_12;
  wire [7:0] t_r25_c24_0;
  wire [7:0] t_r25_c24_1;
  wire [7:0] t_r25_c24_2;
  wire [7:0] t_r25_c24_3;
  wire [7:0] t_r25_c24_4;
  wire [7:0] t_r25_c24_5;
  wire [7:0] t_r25_c24_6;
  wire [7:0] t_r25_c24_7;
  wire [7:0] t_r25_c24_8;
  wire [7:0] t_r25_c24_9;
  wire [7:0] t_r25_c24_10;
  wire [7:0] t_r25_c24_11;
  wire [7:0] t_r25_c24_12;
  wire [7:0] t_r25_c25_0;
  wire [7:0] t_r25_c25_1;
  wire [7:0] t_r25_c25_2;
  wire [7:0] t_r25_c25_3;
  wire [7:0] t_r25_c25_4;
  wire [7:0] t_r25_c25_5;
  wire [7:0] t_r25_c25_6;
  wire [7:0] t_r25_c25_7;
  wire [7:0] t_r25_c25_8;
  wire [7:0] t_r25_c25_9;
  wire [7:0] t_r25_c25_10;
  wire [7:0] t_r25_c25_11;
  wire [7:0] t_r25_c25_12;
  wire [7:0] t_r25_c26_0;
  wire [7:0] t_r25_c26_1;
  wire [7:0] t_r25_c26_2;
  wire [7:0] t_r25_c26_3;
  wire [7:0] t_r25_c26_4;
  wire [7:0] t_r25_c26_5;
  wire [7:0] t_r25_c26_6;
  wire [7:0] t_r25_c26_7;
  wire [7:0] t_r25_c26_8;
  wire [7:0] t_r25_c26_9;
  wire [7:0] t_r25_c26_10;
  wire [7:0] t_r25_c26_11;
  wire [7:0] t_r25_c26_12;
  wire [7:0] t_r25_c27_0;
  wire [7:0] t_r25_c27_1;
  wire [7:0] t_r25_c27_2;
  wire [7:0] t_r25_c27_3;
  wire [7:0] t_r25_c27_4;
  wire [7:0] t_r25_c27_5;
  wire [7:0] t_r25_c27_6;
  wire [7:0] t_r25_c27_7;
  wire [7:0] t_r25_c27_8;
  wire [7:0] t_r25_c27_9;
  wire [7:0] t_r25_c27_10;
  wire [7:0] t_r25_c27_11;
  wire [7:0] t_r25_c27_12;
  wire [7:0] t_r25_c28_0;
  wire [7:0] t_r25_c28_1;
  wire [7:0] t_r25_c28_2;
  wire [7:0] t_r25_c28_3;
  wire [7:0] t_r25_c28_4;
  wire [7:0] t_r25_c28_5;
  wire [7:0] t_r25_c28_6;
  wire [7:0] t_r25_c28_7;
  wire [7:0] t_r25_c28_8;
  wire [7:0] t_r25_c28_9;
  wire [7:0] t_r25_c28_10;
  wire [7:0] t_r25_c28_11;
  wire [7:0] t_r25_c28_12;
  wire [7:0] t_r25_c29_0;
  wire [7:0] t_r25_c29_1;
  wire [7:0] t_r25_c29_2;
  wire [7:0] t_r25_c29_3;
  wire [7:0] t_r25_c29_4;
  wire [7:0] t_r25_c29_5;
  wire [7:0] t_r25_c29_6;
  wire [7:0] t_r25_c29_7;
  wire [7:0] t_r25_c29_8;
  wire [7:0] t_r25_c29_9;
  wire [7:0] t_r25_c29_10;
  wire [7:0] t_r25_c29_11;
  wire [7:0] t_r25_c29_12;
  wire [7:0] t_r25_c30_0;
  wire [7:0] t_r25_c30_1;
  wire [7:0] t_r25_c30_2;
  wire [7:0] t_r25_c30_3;
  wire [7:0] t_r25_c30_4;
  wire [7:0] t_r25_c30_5;
  wire [7:0] t_r25_c30_6;
  wire [7:0] t_r25_c30_7;
  wire [7:0] t_r25_c30_8;
  wire [7:0] t_r25_c30_9;
  wire [7:0] t_r25_c30_10;
  wire [7:0] t_r25_c30_11;
  wire [7:0] t_r25_c30_12;
  wire [7:0] t_r25_c31_0;
  wire [7:0] t_r25_c31_1;
  wire [7:0] t_r25_c31_2;
  wire [7:0] t_r25_c31_3;
  wire [7:0] t_r25_c31_4;
  wire [7:0] t_r25_c31_5;
  wire [7:0] t_r25_c31_6;
  wire [7:0] t_r25_c31_7;
  wire [7:0] t_r25_c31_8;
  wire [7:0] t_r25_c31_9;
  wire [7:0] t_r25_c31_10;
  wire [7:0] t_r25_c31_11;
  wire [7:0] t_r25_c31_12;
  wire [7:0] t_r25_c32_0;
  wire [7:0] t_r25_c32_1;
  wire [7:0] t_r25_c32_2;
  wire [7:0] t_r25_c32_3;
  wire [7:0] t_r25_c32_4;
  wire [7:0] t_r25_c32_5;
  wire [7:0] t_r25_c32_6;
  wire [7:0] t_r25_c32_7;
  wire [7:0] t_r25_c32_8;
  wire [7:0] t_r25_c32_9;
  wire [7:0] t_r25_c32_10;
  wire [7:0] t_r25_c32_11;
  wire [7:0] t_r25_c32_12;
  wire [7:0] t_r25_c33_0;
  wire [7:0] t_r25_c33_1;
  wire [7:0] t_r25_c33_2;
  wire [7:0] t_r25_c33_3;
  wire [7:0] t_r25_c33_4;
  wire [7:0] t_r25_c33_5;
  wire [7:0] t_r25_c33_6;
  wire [7:0] t_r25_c33_7;
  wire [7:0] t_r25_c33_8;
  wire [7:0] t_r25_c33_9;
  wire [7:0] t_r25_c33_10;
  wire [7:0] t_r25_c33_11;
  wire [7:0] t_r25_c33_12;
  wire [7:0] t_r25_c34_0;
  wire [7:0] t_r25_c34_1;
  wire [7:0] t_r25_c34_2;
  wire [7:0] t_r25_c34_3;
  wire [7:0] t_r25_c34_4;
  wire [7:0] t_r25_c34_5;
  wire [7:0] t_r25_c34_6;
  wire [7:0] t_r25_c34_7;
  wire [7:0] t_r25_c34_8;
  wire [7:0] t_r25_c34_9;
  wire [7:0] t_r25_c34_10;
  wire [7:0] t_r25_c34_11;
  wire [7:0] t_r25_c34_12;
  wire [7:0] t_r25_c35_0;
  wire [7:0] t_r25_c35_1;
  wire [7:0] t_r25_c35_2;
  wire [7:0] t_r25_c35_3;
  wire [7:0] t_r25_c35_4;
  wire [7:0] t_r25_c35_5;
  wire [7:0] t_r25_c35_6;
  wire [7:0] t_r25_c35_7;
  wire [7:0] t_r25_c35_8;
  wire [7:0] t_r25_c35_9;
  wire [7:0] t_r25_c35_10;
  wire [7:0] t_r25_c35_11;
  wire [7:0] t_r25_c35_12;
  wire [7:0] t_r25_c36_0;
  wire [7:0] t_r25_c36_1;
  wire [7:0] t_r25_c36_2;
  wire [7:0] t_r25_c36_3;
  wire [7:0] t_r25_c36_4;
  wire [7:0] t_r25_c36_5;
  wire [7:0] t_r25_c36_6;
  wire [7:0] t_r25_c36_7;
  wire [7:0] t_r25_c36_8;
  wire [7:0] t_r25_c36_9;
  wire [7:0] t_r25_c36_10;
  wire [7:0] t_r25_c36_11;
  wire [7:0] t_r25_c36_12;
  wire [7:0] t_r25_c37_0;
  wire [7:0] t_r25_c37_1;
  wire [7:0] t_r25_c37_2;
  wire [7:0] t_r25_c37_3;
  wire [7:0] t_r25_c37_4;
  wire [7:0] t_r25_c37_5;
  wire [7:0] t_r25_c37_6;
  wire [7:0] t_r25_c37_7;
  wire [7:0] t_r25_c37_8;
  wire [7:0] t_r25_c37_9;
  wire [7:0] t_r25_c37_10;
  wire [7:0] t_r25_c37_11;
  wire [7:0] t_r25_c37_12;
  wire [7:0] t_r25_c38_0;
  wire [7:0] t_r25_c38_1;
  wire [7:0] t_r25_c38_2;
  wire [7:0] t_r25_c38_3;
  wire [7:0] t_r25_c38_4;
  wire [7:0] t_r25_c38_5;
  wire [7:0] t_r25_c38_6;
  wire [7:0] t_r25_c38_7;
  wire [7:0] t_r25_c38_8;
  wire [7:0] t_r25_c38_9;
  wire [7:0] t_r25_c38_10;
  wire [7:0] t_r25_c38_11;
  wire [7:0] t_r25_c38_12;
  wire [7:0] t_r25_c39_0;
  wire [7:0] t_r25_c39_1;
  wire [7:0] t_r25_c39_2;
  wire [7:0] t_r25_c39_3;
  wire [7:0] t_r25_c39_4;
  wire [7:0] t_r25_c39_5;
  wire [7:0] t_r25_c39_6;
  wire [7:0] t_r25_c39_7;
  wire [7:0] t_r25_c39_8;
  wire [7:0] t_r25_c39_9;
  wire [7:0] t_r25_c39_10;
  wire [7:0] t_r25_c39_11;
  wire [7:0] t_r25_c39_12;
  wire [7:0] t_r25_c40_0;
  wire [7:0] t_r25_c40_1;
  wire [7:0] t_r25_c40_2;
  wire [7:0] t_r25_c40_3;
  wire [7:0] t_r25_c40_4;
  wire [7:0] t_r25_c40_5;
  wire [7:0] t_r25_c40_6;
  wire [7:0] t_r25_c40_7;
  wire [7:0] t_r25_c40_8;
  wire [7:0] t_r25_c40_9;
  wire [7:0] t_r25_c40_10;
  wire [7:0] t_r25_c40_11;
  wire [7:0] t_r25_c40_12;
  wire [7:0] t_r25_c41_0;
  wire [7:0] t_r25_c41_1;
  wire [7:0] t_r25_c41_2;
  wire [7:0] t_r25_c41_3;
  wire [7:0] t_r25_c41_4;
  wire [7:0] t_r25_c41_5;
  wire [7:0] t_r25_c41_6;
  wire [7:0] t_r25_c41_7;
  wire [7:0] t_r25_c41_8;
  wire [7:0] t_r25_c41_9;
  wire [7:0] t_r25_c41_10;
  wire [7:0] t_r25_c41_11;
  wire [7:0] t_r25_c41_12;
  wire [7:0] t_r25_c42_0;
  wire [7:0] t_r25_c42_1;
  wire [7:0] t_r25_c42_2;
  wire [7:0] t_r25_c42_3;
  wire [7:0] t_r25_c42_4;
  wire [7:0] t_r25_c42_5;
  wire [7:0] t_r25_c42_6;
  wire [7:0] t_r25_c42_7;
  wire [7:0] t_r25_c42_8;
  wire [7:0] t_r25_c42_9;
  wire [7:0] t_r25_c42_10;
  wire [7:0] t_r25_c42_11;
  wire [7:0] t_r25_c42_12;
  wire [7:0] t_r25_c43_0;
  wire [7:0] t_r25_c43_1;
  wire [7:0] t_r25_c43_2;
  wire [7:0] t_r25_c43_3;
  wire [7:0] t_r25_c43_4;
  wire [7:0] t_r25_c43_5;
  wire [7:0] t_r25_c43_6;
  wire [7:0] t_r25_c43_7;
  wire [7:0] t_r25_c43_8;
  wire [7:0] t_r25_c43_9;
  wire [7:0] t_r25_c43_10;
  wire [7:0] t_r25_c43_11;
  wire [7:0] t_r25_c43_12;
  wire [7:0] t_r25_c44_0;
  wire [7:0] t_r25_c44_1;
  wire [7:0] t_r25_c44_2;
  wire [7:0] t_r25_c44_3;
  wire [7:0] t_r25_c44_4;
  wire [7:0] t_r25_c44_5;
  wire [7:0] t_r25_c44_6;
  wire [7:0] t_r25_c44_7;
  wire [7:0] t_r25_c44_8;
  wire [7:0] t_r25_c44_9;
  wire [7:0] t_r25_c44_10;
  wire [7:0] t_r25_c44_11;
  wire [7:0] t_r25_c44_12;
  wire [7:0] t_r25_c45_0;
  wire [7:0] t_r25_c45_1;
  wire [7:0] t_r25_c45_2;
  wire [7:0] t_r25_c45_3;
  wire [7:0] t_r25_c45_4;
  wire [7:0] t_r25_c45_5;
  wire [7:0] t_r25_c45_6;
  wire [7:0] t_r25_c45_7;
  wire [7:0] t_r25_c45_8;
  wire [7:0] t_r25_c45_9;
  wire [7:0] t_r25_c45_10;
  wire [7:0] t_r25_c45_11;
  wire [7:0] t_r25_c45_12;
  wire [7:0] t_r25_c46_0;
  wire [7:0] t_r25_c46_1;
  wire [7:0] t_r25_c46_2;
  wire [7:0] t_r25_c46_3;
  wire [7:0] t_r25_c46_4;
  wire [7:0] t_r25_c46_5;
  wire [7:0] t_r25_c46_6;
  wire [7:0] t_r25_c46_7;
  wire [7:0] t_r25_c46_8;
  wire [7:0] t_r25_c46_9;
  wire [7:0] t_r25_c46_10;
  wire [7:0] t_r25_c46_11;
  wire [7:0] t_r25_c46_12;
  wire [7:0] t_r25_c47_0;
  wire [7:0] t_r25_c47_1;
  wire [7:0] t_r25_c47_2;
  wire [7:0] t_r25_c47_3;
  wire [7:0] t_r25_c47_4;
  wire [7:0] t_r25_c47_5;
  wire [7:0] t_r25_c47_6;
  wire [7:0] t_r25_c47_7;
  wire [7:0] t_r25_c47_8;
  wire [7:0] t_r25_c47_9;
  wire [7:0] t_r25_c47_10;
  wire [7:0] t_r25_c47_11;
  wire [7:0] t_r25_c47_12;
  wire [7:0] t_r25_c48_0;
  wire [7:0] t_r25_c48_1;
  wire [7:0] t_r25_c48_2;
  wire [7:0] t_r25_c48_3;
  wire [7:0] t_r25_c48_4;
  wire [7:0] t_r25_c48_5;
  wire [7:0] t_r25_c48_6;
  wire [7:0] t_r25_c48_7;
  wire [7:0] t_r25_c48_8;
  wire [7:0] t_r25_c48_9;
  wire [7:0] t_r25_c48_10;
  wire [7:0] t_r25_c48_11;
  wire [7:0] t_r25_c48_12;
  wire [7:0] t_r25_c49_0;
  wire [7:0] t_r25_c49_1;
  wire [7:0] t_r25_c49_2;
  wire [7:0] t_r25_c49_3;
  wire [7:0] t_r25_c49_4;
  wire [7:0] t_r25_c49_5;
  wire [7:0] t_r25_c49_6;
  wire [7:0] t_r25_c49_7;
  wire [7:0] t_r25_c49_8;
  wire [7:0] t_r25_c49_9;
  wire [7:0] t_r25_c49_10;
  wire [7:0] t_r25_c49_11;
  wire [7:0] t_r25_c49_12;
  wire [7:0] t_r25_c50_0;
  wire [7:0] t_r25_c50_1;
  wire [7:0] t_r25_c50_2;
  wire [7:0] t_r25_c50_3;
  wire [7:0] t_r25_c50_4;
  wire [7:0] t_r25_c50_5;
  wire [7:0] t_r25_c50_6;
  wire [7:0] t_r25_c50_7;
  wire [7:0] t_r25_c50_8;
  wire [7:0] t_r25_c50_9;
  wire [7:0] t_r25_c50_10;
  wire [7:0] t_r25_c50_11;
  wire [7:0] t_r25_c50_12;
  wire [7:0] t_r25_c51_0;
  wire [7:0] t_r25_c51_1;
  wire [7:0] t_r25_c51_2;
  wire [7:0] t_r25_c51_3;
  wire [7:0] t_r25_c51_4;
  wire [7:0] t_r25_c51_5;
  wire [7:0] t_r25_c51_6;
  wire [7:0] t_r25_c51_7;
  wire [7:0] t_r25_c51_8;
  wire [7:0] t_r25_c51_9;
  wire [7:0] t_r25_c51_10;
  wire [7:0] t_r25_c51_11;
  wire [7:0] t_r25_c51_12;
  wire [7:0] t_r25_c52_0;
  wire [7:0] t_r25_c52_1;
  wire [7:0] t_r25_c52_2;
  wire [7:0] t_r25_c52_3;
  wire [7:0] t_r25_c52_4;
  wire [7:0] t_r25_c52_5;
  wire [7:0] t_r25_c52_6;
  wire [7:0] t_r25_c52_7;
  wire [7:0] t_r25_c52_8;
  wire [7:0] t_r25_c52_9;
  wire [7:0] t_r25_c52_10;
  wire [7:0] t_r25_c52_11;
  wire [7:0] t_r25_c52_12;
  wire [7:0] t_r25_c53_0;
  wire [7:0] t_r25_c53_1;
  wire [7:0] t_r25_c53_2;
  wire [7:0] t_r25_c53_3;
  wire [7:0] t_r25_c53_4;
  wire [7:0] t_r25_c53_5;
  wire [7:0] t_r25_c53_6;
  wire [7:0] t_r25_c53_7;
  wire [7:0] t_r25_c53_8;
  wire [7:0] t_r25_c53_9;
  wire [7:0] t_r25_c53_10;
  wire [7:0] t_r25_c53_11;
  wire [7:0] t_r25_c53_12;
  wire [7:0] t_r25_c54_0;
  wire [7:0] t_r25_c54_1;
  wire [7:0] t_r25_c54_2;
  wire [7:0] t_r25_c54_3;
  wire [7:0] t_r25_c54_4;
  wire [7:0] t_r25_c54_5;
  wire [7:0] t_r25_c54_6;
  wire [7:0] t_r25_c54_7;
  wire [7:0] t_r25_c54_8;
  wire [7:0] t_r25_c54_9;
  wire [7:0] t_r25_c54_10;
  wire [7:0] t_r25_c54_11;
  wire [7:0] t_r25_c54_12;
  wire [7:0] t_r25_c55_0;
  wire [7:0] t_r25_c55_1;
  wire [7:0] t_r25_c55_2;
  wire [7:0] t_r25_c55_3;
  wire [7:0] t_r25_c55_4;
  wire [7:0] t_r25_c55_5;
  wire [7:0] t_r25_c55_6;
  wire [7:0] t_r25_c55_7;
  wire [7:0] t_r25_c55_8;
  wire [7:0] t_r25_c55_9;
  wire [7:0] t_r25_c55_10;
  wire [7:0] t_r25_c55_11;
  wire [7:0] t_r25_c55_12;
  wire [7:0] t_r25_c56_0;
  wire [7:0] t_r25_c56_1;
  wire [7:0] t_r25_c56_2;
  wire [7:0] t_r25_c56_3;
  wire [7:0] t_r25_c56_4;
  wire [7:0] t_r25_c56_5;
  wire [7:0] t_r25_c56_6;
  wire [7:0] t_r25_c56_7;
  wire [7:0] t_r25_c56_8;
  wire [7:0] t_r25_c56_9;
  wire [7:0] t_r25_c56_10;
  wire [7:0] t_r25_c56_11;
  wire [7:0] t_r25_c56_12;
  wire [7:0] t_r25_c57_0;
  wire [7:0] t_r25_c57_1;
  wire [7:0] t_r25_c57_2;
  wire [7:0] t_r25_c57_3;
  wire [7:0] t_r25_c57_4;
  wire [7:0] t_r25_c57_5;
  wire [7:0] t_r25_c57_6;
  wire [7:0] t_r25_c57_7;
  wire [7:0] t_r25_c57_8;
  wire [7:0] t_r25_c57_9;
  wire [7:0] t_r25_c57_10;
  wire [7:0] t_r25_c57_11;
  wire [7:0] t_r25_c57_12;
  wire [7:0] t_r25_c58_0;
  wire [7:0] t_r25_c58_1;
  wire [7:0] t_r25_c58_2;
  wire [7:0] t_r25_c58_3;
  wire [7:0] t_r25_c58_4;
  wire [7:0] t_r25_c58_5;
  wire [7:0] t_r25_c58_6;
  wire [7:0] t_r25_c58_7;
  wire [7:0] t_r25_c58_8;
  wire [7:0] t_r25_c58_9;
  wire [7:0] t_r25_c58_10;
  wire [7:0] t_r25_c58_11;
  wire [7:0] t_r25_c58_12;
  wire [7:0] t_r25_c59_0;
  wire [7:0] t_r25_c59_1;
  wire [7:0] t_r25_c59_2;
  wire [7:0] t_r25_c59_3;
  wire [7:0] t_r25_c59_4;
  wire [7:0] t_r25_c59_5;
  wire [7:0] t_r25_c59_6;
  wire [7:0] t_r25_c59_7;
  wire [7:0] t_r25_c59_8;
  wire [7:0] t_r25_c59_9;
  wire [7:0] t_r25_c59_10;
  wire [7:0] t_r25_c59_11;
  wire [7:0] t_r25_c59_12;
  wire [7:0] t_r25_c60_0;
  wire [7:0] t_r25_c60_1;
  wire [7:0] t_r25_c60_2;
  wire [7:0] t_r25_c60_3;
  wire [7:0] t_r25_c60_4;
  wire [7:0] t_r25_c60_5;
  wire [7:0] t_r25_c60_6;
  wire [7:0] t_r25_c60_7;
  wire [7:0] t_r25_c60_8;
  wire [7:0] t_r25_c60_9;
  wire [7:0] t_r25_c60_10;
  wire [7:0] t_r25_c60_11;
  wire [7:0] t_r25_c60_12;
  wire [7:0] t_r25_c61_0;
  wire [7:0] t_r25_c61_1;
  wire [7:0] t_r25_c61_2;
  wire [7:0] t_r25_c61_3;
  wire [7:0] t_r25_c61_4;
  wire [7:0] t_r25_c61_5;
  wire [7:0] t_r25_c61_6;
  wire [7:0] t_r25_c61_7;
  wire [7:0] t_r25_c61_8;
  wire [7:0] t_r25_c61_9;
  wire [7:0] t_r25_c61_10;
  wire [7:0] t_r25_c61_11;
  wire [7:0] t_r25_c61_12;
  wire [7:0] t_r25_c62_0;
  wire [7:0] t_r25_c62_1;
  wire [7:0] t_r25_c62_2;
  wire [7:0] t_r25_c62_3;
  wire [7:0] t_r25_c62_4;
  wire [7:0] t_r25_c62_5;
  wire [7:0] t_r25_c62_6;
  wire [7:0] t_r25_c62_7;
  wire [7:0] t_r25_c62_8;
  wire [7:0] t_r25_c62_9;
  wire [7:0] t_r25_c62_10;
  wire [7:0] t_r25_c62_11;
  wire [7:0] t_r25_c62_12;
  wire [7:0] t_r25_c63_0;
  wire [7:0] t_r25_c63_1;
  wire [7:0] t_r25_c63_2;
  wire [7:0] t_r25_c63_3;
  wire [7:0] t_r25_c63_4;
  wire [7:0] t_r25_c63_5;
  wire [7:0] t_r25_c63_6;
  wire [7:0] t_r25_c63_7;
  wire [7:0] t_r25_c63_8;
  wire [7:0] t_r25_c63_9;
  wire [7:0] t_r25_c63_10;
  wire [7:0] t_r25_c63_11;
  wire [7:0] t_r25_c63_12;
  wire [7:0] t_r25_c64_0;
  wire [7:0] t_r25_c64_1;
  wire [7:0] t_r25_c64_2;
  wire [7:0] t_r25_c64_3;
  wire [7:0] t_r25_c64_4;
  wire [7:0] t_r25_c64_5;
  wire [7:0] t_r25_c64_6;
  wire [7:0] t_r25_c64_7;
  wire [7:0] t_r25_c64_8;
  wire [7:0] t_r25_c64_9;
  wire [7:0] t_r25_c64_10;
  wire [7:0] t_r25_c64_11;
  wire [7:0] t_r25_c64_12;
  wire [7:0] t_r25_c65_0;
  wire [7:0] t_r25_c65_1;
  wire [7:0] t_r25_c65_2;
  wire [7:0] t_r25_c65_3;
  wire [7:0] t_r25_c65_4;
  wire [7:0] t_r25_c65_5;
  wire [7:0] t_r25_c65_6;
  wire [7:0] t_r25_c65_7;
  wire [7:0] t_r25_c65_8;
  wire [7:0] t_r25_c65_9;
  wire [7:0] t_r25_c65_10;
  wire [7:0] t_r25_c65_11;
  wire [7:0] t_r25_c65_12;
  wire [7:0] t_r26_c0_0;
  wire [7:0] t_r26_c0_1;
  wire [7:0] t_r26_c0_2;
  wire [7:0] t_r26_c0_3;
  wire [7:0] t_r26_c0_4;
  wire [7:0] t_r26_c0_5;
  wire [7:0] t_r26_c0_6;
  wire [7:0] t_r26_c0_7;
  wire [7:0] t_r26_c0_8;
  wire [7:0] t_r26_c0_9;
  wire [7:0] t_r26_c0_10;
  wire [7:0] t_r26_c0_11;
  wire [7:0] t_r26_c0_12;
  wire [7:0] t_r26_c1_0;
  wire [7:0] t_r26_c1_1;
  wire [7:0] t_r26_c1_2;
  wire [7:0] t_r26_c1_3;
  wire [7:0] t_r26_c1_4;
  wire [7:0] t_r26_c1_5;
  wire [7:0] t_r26_c1_6;
  wire [7:0] t_r26_c1_7;
  wire [7:0] t_r26_c1_8;
  wire [7:0] t_r26_c1_9;
  wire [7:0] t_r26_c1_10;
  wire [7:0] t_r26_c1_11;
  wire [7:0] t_r26_c1_12;
  wire [7:0] t_r26_c2_0;
  wire [7:0] t_r26_c2_1;
  wire [7:0] t_r26_c2_2;
  wire [7:0] t_r26_c2_3;
  wire [7:0] t_r26_c2_4;
  wire [7:0] t_r26_c2_5;
  wire [7:0] t_r26_c2_6;
  wire [7:0] t_r26_c2_7;
  wire [7:0] t_r26_c2_8;
  wire [7:0] t_r26_c2_9;
  wire [7:0] t_r26_c2_10;
  wire [7:0] t_r26_c2_11;
  wire [7:0] t_r26_c2_12;
  wire [7:0] t_r26_c3_0;
  wire [7:0] t_r26_c3_1;
  wire [7:0] t_r26_c3_2;
  wire [7:0] t_r26_c3_3;
  wire [7:0] t_r26_c3_4;
  wire [7:0] t_r26_c3_5;
  wire [7:0] t_r26_c3_6;
  wire [7:0] t_r26_c3_7;
  wire [7:0] t_r26_c3_8;
  wire [7:0] t_r26_c3_9;
  wire [7:0] t_r26_c3_10;
  wire [7:0] t_r26_c3_11;
  wire [7:0] t_r26_c3_12;
  wire [7:0] t_r26_c4_0;
  wire [7:0] t_r26_c4_1;
  wire [7:0] t_r26_c4_2;
  wire [7:0] t_r26_c4_3;
  wire [7:0] t_r26_c4_4;
  wire [7:0] t_r26_c4_5;
  wire [7:0] t_r26_c4_6;
  wire [7:0] t_r26_c4_7;
  wire [7:0] t_r26_c4_8;
  wire [7:0] t_r26_c4_9;
  wire [7:0] t_r26_c4_10;
  wire [7:0] t_r26_c4_11;
  wire [7:0] t_r26_c4_12;
  wire [7:0] t_r26_c5_0;
  wire [7:0] t_r26_c5_1;
  wire [7:0] t_r26_c5_2;
  wire [7:0] t_r26_c5_3;
  wire [7:0] t_r26_c5_4;
  wire [7:0] t_r26_c5_5;
  wire [7:0] t_r26_c5_6;
  wire [7:0] t_r26_c5_7;
  wire [7:0] t_r26_c5_8;
  wire [7:0] t_r26_c5_9;
  wire [7:0] t_r26_c5_10;
  wire [7:0] t_r26_c5_11;
  wire [7:0] t_r26_c5_12;
  wire [7:0] t_r26_c6_0;
  wire [7:0] t_r26_c6_1;
  wire [7:0] t_r26_c6_2;
  wire [7:0] t_r26_c6_3;
  wire [7:0] t_r26_c6_4;
  wire [7:0] t_r26_c6_5;
  wire [7:0] t_r26_c6_6;
  wire [7:0] t_r26_c6_7;
  wire [7:0] t_r26_c6_8;
  wire [7:0] t_r26_c6_9;
  wire [7:0] t_r26_c6_10;
  wire [7:0] t_r26_c6_11;
  wire [7:0] t_r26_c6_12;
  wire [7:0] t_r26_c7_0;
  wire [7:0] t_r26_c7_1;
  wire [7:0] t_r26_c7_2;
  wire [7:0] t_r26_c7_3;
  wire [7:0] t_r26_c7_4;
  wire [7:0] t_r26_c7_5;
  wire [7:0] t_r26_c7_6;
  wire [7:0] t_r26_c7_7;
  wire [7:0] t_r26_c7_8;
  wire [7:0] t_r26_c7_9;
  wire [7:0] t_r26_c7_10;
  wire [7:0] t_r26_c7_11;
  wire [7:0] t_r26_c7_12;
  wire [7:0] t_r26_c8_0;
  wire [7:0] t_r26_c8_1;
  wire [7:0] t_r26_c8_2;
  wire [7:0] t_r26_c8_3;
  wire [7:0] t_r26_c8_4;
  wire [7:0] t_r26_c8_5;
  wire [7:0] t_r26_c8_6;
  wire [7:0] t_r26_c8_7;
  wire [7:0] t_r26_c8_8;
  wire [7:0] t_r26_c8_9;
  wire [7:0] t_r26_c8_10;
  wire [7:0] t_r26_c8_11;
  wire [7:0] t_r26_c8_12;
  wire [7:0] t_r26_c9_0;
  wire [7:0] t_r26_c9_1;
  wire [7:0] t_r26_c9_2;
  wire [7:0] t_r26_c9_3;
  wire [7:0] t_r26_c9_4;
  wire [7:0] t_r26_c9_5;
  wire [7:0] t_r26_c9_6;
  wire [7:0] t_r26_c9_7;
  wire [7:0] t_r26_c9_8;
  wire [7:0] t_r26_c9_9;
  wire [7:0] t_r26_c9_10;
  wire [7:0] t_r26_c9_11;
  wire [7:0] t_r26_c9_12;
  wire [7:0] t_r26_c10_0;
  wire [7:0] t_r26_c10_1;
  wire [7:0] t_r26_c10_2;
  wire [7:0] t_r26_c10_3;
  wire [7:0] t_r26_c10_4;
  wire [7:0] t_r26_c10_5;
  wire [7:0] t_r26_c10_6;
  wire [7:0] t_r26_c10_7;
  wire [7:0] t_r26_c10_8;
  wire [7:0] t_r26_c10_9;
  wire [7:0] t_r26_c10_10;
  wire [7:0] t_r26_c10_11;
  wire [7:0] t_r26_c10_12;
  wire [7:0] t_r26_c11_0;
  wire [7:0] t_r26_c11_1;
  wire [7:0] t_r26_c11_2;
  wire [7:0] t_r26_c11_3;
  wire [7:0] t_r26_c11_4;
  wire [7:0] t_r26_c11_5;
  wire [7:0] t_r26_c11_6;
  wire [7:0] t_r26_c11_7;
  wire [7:0] t_r26_c11_8;
  wire [7:0] t_r26_c11_9;
  wire [7:0] t_r26_c11_10;
  wire [7:0] t_r26_c11_11;
  wire [7:0] t_r26_c11_12;
  wire [7:0] t_r26_c12_0;
  wire [7:0] t_r26_c12_1;
  wire [7:0] t_r26_c12_2;
  wire [7:0] t_r26_c12_3;
  wire [7:0] t_r26_c12_4;
  wire [7:0] t_r26_c12_5;
  wire [7:0] t_r26_c12_6;
  wire [7:0] t_r26_c12_7;
  wire [7:0] t_r26_c12_8;
  wire [7:0] t_r26_c12_9;
  wire [7:0] t_r26_c12_10;
  wire [7:0] t_r26_c12_11;
  wire [7:0] t_r26_c12_12;
  wire [7:0] t_r26_c13_0;
  wire [7:0] t_r26_c13_1;
  wire [7:0] t_r26_c13_2;
  wire [7:0] t_r26_c13_3;
  wire [7:0] t_r26_c13_4;
  wire [7:0] t_r26_c13_5;
  wire [7:0] t_r26_c13_6;
  wire [7:0] t_r26_c13_7;
  wire [7:0] t_r26_c13_8;
  wire [7:0] t_r26_c13_9;
  wire [7:0] t_r26_c13_10;
  wire [7:0] t_r26_c13_11;
  wire [7:0] t_r26_c13_12;
  wire [7:0] t_r26_c14_0;
  wire [7:0] t_r26_c14_1;
  wire [7:0] t_r26_c14_2;
  wire [7:0] t_r26_c14_3;
  wire [7:0] t_r26_c14_4;
  wire [7:0] t_r26_c14_5;
  wire [7:0] t_r26_c14_6;
  wire [7:0] t_r26_c14_7;
  wire [7:0] t_r26_c14_8;
  wire [7:0] t_r26_c14_9;
  wire [7:0] t_r26_c14_10;
  wire [7:0] t_r26_c14_11;
  wire [7:0] t_r26_c14_12;
  wire [7:0] t_r26_c15_0;
  wire [7:0] t_r26_c15_1;
  wire [7:0] t_r26_c15_2;
  wire [7:0] t_r26_c15_3;
  wire [7:0] t_r26_c15_4;
  wire [7:0] t_r26_c15_5;
  wire [7:0] t_r26_c15_6;
  wire [7:0] t_r26_c15_7;
  wire [7:0] t_r26_c15_8;
  wire [7:0] t_r26_c15_9;
  wire [7:0] t_r26_c15_10;
  wire [7:0] t_r26_c15_11;
  wire [7:0] t_r26_c15_12;
  wire [7:0] t_r26_c16_0;
  wire [7:0] t_r26_c16_1;
  wire [7:0] t_r26_c16_2;
  wire [7:0] t_r26_c16_3;
  wire [7:0] t_r26_c16_4;
  wire [7:0] t_r26_c16_5;
  wire [7:0] t_r26_c16_6;
  wire [7:0] t_r26_c16_7;
  wire [7:0] t_r26_c16_8;
  wire [7:0] t_r26_c16_9;
  wire [7:0] t_r26_c16_10;
  wire [7:0] t_r26_c16_11;
  wire [7:0] t_r26_c16_12;
  wire [7:0] t_r26_c17_0;
  wire [7:0] t_r26_c17_1;
  wire [7:0] t_r26_c17_2;
  wire [7:0] t_r26_c17_3;
  wire [7:0] t_r26_c17_4;
  wire [7:0] t_r26_c17_5;
  wire [7:0] t_r26_c17_6;
  wire [7:0] t_r26_c17_7;
  wire [7:0] t_r26_c17_8;
  wire [7:0] t_r26_c17_9;
  wire [7:0] t_r26_c17_10;
  wire [7:0] t_r26_c17_11;
  wire [7:0] t_r26_c17_12;
  wire [7:0] t_r26_c18_0;
  wire [7:0] t_r26_c18_1;
  wire [7:0] t_r26_c18_2;
  wire [7:0] t_r26_c18_3;
  wire [7:0] t_r26_c18_4;
  wire [7:0] t_r26_c18_5;
  wire [7:0] t_r26_c18_6;
  wire [7:0] t_r26_c18_7;
  wire [7:0] t_r26_c18_8;
  wire [7:0] t_r26_c18_9;
  wire [7:0] t_r26_c18_10;
  wire [7:0] t_r26_c18_11;
  wire [7:0] t_r26_c18_12;
  wire [7:0] t_r26_c19_0;
  wire [7:0] t_r26_c19_1;
  wire [7:0] t_r26_c19_2;
  wire [7:0] t_r26_c19_3;
  wire [7:0] t_r26_c19_4;
  wire [7:0] t_r26_c19_5;
  wire [7:0] t_r26_c19_6;
  wire [7:0] t_r26_c19_7;
  wire [7:0] t_r26_c19_8;
  wire [7:0] t_r26_c19_9;
  wire [7:0] t_r26_c19_10;
  wire [7:0] t_r26_c19_11;
  wire [7:0] t_r26_c19_12;
  wire [7:0] t_r26_c20_0;
  wire [7:0] t_r26_c20_1;
  wire [7:0] t_r26_c20_2;
  wire [7:0] t_r26_c20_3;
  wire [7:0] t_r26_c20_4;
  wire [7:0] t_r26_c20_5;
  wire [7:0] t_r26_c20_6;
  wire [7:0] t_r26_c20_7;
  wire [7:0] t_r26_c20_8;
  wire [7:0] t_r26_c20_9;
  wire [7:0] t_r26_c20_10;
  wire [7:0] t_r26_c20_11;
  wire [7:0] t_r26_c20_12;
  wire [7:0] t_r26_c21_0;
  wire [7:0] t_r26_c21_1;
  wire [7:0] t_r26_c21_2;
  wire [7:0] t_r26_c21_3;
  wire [7:0] t_r26_c21_4;
  wire [7:0] t_r26_c21_5;
  wire [7:0] t_r26_c21_6;
  wire [7:0] t_r26_c21_7;
  wire [7:0] t_r26_c21_8;
  wire [7:0] t_r26_c21_9;
  wire [7:0] t_r26_c21_10;
  wire [7:0] t_r26_c21_11;
  wire [7:0] t_r26_c21_12;
  wire [7:0] t_r26_c22_0;
  wire [7:0] t_r26_c22_1;
  wire [7:0] t_r26_c22_2;
  wire [7:0] t_r26_c22_3;
  wire [7:0] t_r26_c22_4;
  wire [7:0] t_r26_c22_5;
  wire [7:0] t_r26_c22_6;
  wire [7:0] t_r26_c22_7;
  wire [7:0] t_r26_c22_8;
  wire [7:0] t_r26_c22_9;
  wire [7:0] t_r26_c22_10;
  wire [7:0] t_r26_c22_11;
  wire [7:0] t_r26_c22_12;
  wire [7:0] t_r26_c23_0;
  wire [7:0] t_r26_c23_1;
  wire [7:0] t_r26_c23_2;
  wire [7:0] t_r26_c23_3;
  wire [7:0] t_r26_c23_4;
  wire [7:0] t_r26_c23_5;
  wire [7:0] t_r26_c23_6;
  wire [7:0] t_r26_c23_7;
  wire [7:0] t_r26_c23_8;
  wire [7:0] t_r26_c23_9;
  wire [7:0] t_r26_c23_10;
  wire [7:0] t_r26_c23_11;
  wire [7:0] t_r26_c23_12;
  wire [7:0] t_r26_c24_0;
  wire [7:0] t_r26_c24_1;
  wire [7:0] t_r26_c24_2;
  wire [7:0] t_r26_c24_3;
  wire [7:0] t_r26_c24_4;
  wire [7:0] t_r26_c24_5;
  wire [7:0] t_r26_c24_6;
  wire [7:0] t_r26_c24_7;
  wire [7:0] t_r26_c24_8;
  wire [7:0] t_r26_c24_9;
  wire [7:0] t_r26_c24_10;
  wire [7:0] t_r26_c24_11;
  wire [7:0] t_r26_c24_12;
  wire [7:0] t_r26_c25_0;
  wire [7:0] t_r26_c25_1;
  wire [7:0] t_r26_c25_2;
  wire [7:0] t_r26_c25_3;
  wire [7:0] t_r26_c25_4;
  wire [7:0] t_r26_c25_5;
  wire [7:0] t_r26_c25_6;
  wire [7:0] t_r26_c25_7;
  wire [7:0] t_r26_c25_8;
  wire [7:0] t_r26_c25_9;
  wire [7:0] t_r26_c25_10;
  wire [7:0] t_r26_c25_11;
  wire [7:0] t_r26_c25_12;
  wire [7:0] t_r26_c26_0;
  wire [7:0] t_r26_c26_1;
  wire [7:0] t_r26_c26_2;
  wire [7:0] t_r26_c26_3;
  wire [7:0] t_r26_c26_4;
  wire [7:0] t_r26_c26_5;
  wire [7:0] t_r26_c26_6;
  wire [7:0] t_r26_c26_7;
  wire [7:0] t_r26_c26_8;
  wire [7:0] t_r26_c26_9;
  wire [7:0] t_r26_c26_10;
  wire [7:0] t_r26_c26_11;
  wire [7:0] t_r26_c26_12;
  wire [7:0] t_r26_c27_0;
  wire [7:0] t_r26_c27_1;
  wire [7:0] t_r26_c27_2;
  wire [7:0] t_r26_c27_3;
  wire [7:0] t_r26_c27_4;
  wire [7:0] t_r26_c27_5;
  wire [7:0] t_r26_c27_6;
  wire [7:0] t_r26_c27_7;
  wire [7:0] t_r26_c27_8;
  wire [7:0] t_r26_c27_9;
  wire [7:0] t_r26_c27_10;
  wire [7:0] t_r26_c27_11;
  wire [7:0] t_r26_c27_12;
  wire [7:0] t_r26_c28_0;
  wire [7:0] t_r26_c28_1;
  wire [7:0] t_r26_c28_2;
  wire [7:0] t_r26_c28_3;
  wire [7:0] t_r26_c28_4;
  wire [7:0] t_r26_c28_5;
  wire [7:0] t_r26_c28_6;
  wire [7:0] t_r26_c28_7;
  wire [7:0] t_r26_c28_8;
  wire [7:0] t_r26_c28_9;
  wire [7:0] t_r26_c28_10;
  wire [7:0] t_r26_c28_11;
  wire [7:0] t_r26_c28_12;
  wire [7:0] t_r26_c29_0;
  wire [7:0] t_r26_c29_1;
  wire [7:0] t_r26_c29_2;
  wire [7:0] t_r26_c29_3;
  wire [7:0] t_r26_c29_4;
  wire [7:0] t_r26_c29_5;
  wire [7:0] t_r26_c29_6;
  wire [7:0] t_r26_c29_7;
  wire [7:0] t_r26_c29_8;
  wire [7:0] t_r26_c29_9;
  wire [7:0] t_r26_c29_10;
  wire [7:0] t_r26_c29_11;
  wire [7:0] t_r26_c29_12;
  wire [7:0] t_r26_c30_0;
  wire [7:0] t_r26_c30_1;
  wire [7:0] t_r26_c30_2;
  wire [7:0] t_r26_c30_3;
  wire [7:0] t_r26_c30_4;
  wire [7:0] t_r26_c30_5;
  wire [7:0] t_r26_c30_6;
  wire [7:0] t_r26_c30_7;
  wire [7:0] t_r26_c30_8;
  wire [7:0] t_r26_c30_9;
  wire [7:0] t_r26_c30_10;
  wire [7:0] t_r26_c30_11;
  wire [7:0] t_r26_c30_12;
  wire [7:0] t_r26_c31_0;
  wire [7:0] t_r26_c31_1;
  wire [7:0] t_r26_c31_2;
  wire [7:0] t_r26_c31_3;
  wire [7:0] t_r26_c31_4;
  wire [7:0] t_r26_c31_5;
  wire [7:0] t_r26_c31_6;
  wire [7:0] t_r26_c31_7;
  wire [7:0] t_r26_c31_8;
  wire [7:0] t_r26_c31_9;
  wire [7:0] t_r26_c31_10;
  wire [7:0] t_r26_c31_11;
  wire [7:0] t_r26_c31_12;
  wire [7:0] t_r26_c32_0;
  wire [7:0] t_r26_c32_1;
  wire [7:0] t_r26_c32_2;
  wire [7:0] t_r26_c32_3;
  wire [7:0] t_r26_c32_4;
  wire [7:0] t_r26_c32_5;
  wire [7:0] t_r26_c32_6;
  wire [7:0] t_r26_c32_7;
  wire [7:0] t_r26_c32_8;
  wire [7:0] t_r26_c32_9;
  wire [7:0] t_r26_c32_10;
  wire [7:0] t_r26_c32_11;
  wire [7:0] t_r26_c32_12;
  wire [7:0] t_r26_c33_0;
  wire [7:0] t_r26_c33_1;
  wire [7:0] t_r26_c33_2;
  wire [7:0] t_r26_c33_3;
  wire [7:0] t_r26_c33_4;
  wire [7:0] t_r26_c33_5;
  wire [7:0] t_r26_c33_6;
  wire [7:0] t_r26_c33_7;
  wire [7:0] t_r26_c33_8;
  wire [7:0] t_r26_c33_9;
  wire [7:0] t_r26_c33_10;
  wire [7:0] t_r26_c33_11;
  wire [7:0] t_r26_c33_12;
  wire [7:0] t_r26_c34_0;
  wire [7:0] t_r26_c34_1;
  wire [7:0] t_r26_c34_2;
  wire [7:0] t_r26_c34_3;
  wire [7:0] t_r26_c34_4;
  wire [7:0] t_r26_c34_5;
  wire [7:0] t_r26_c34_6;
  wire [7:0] t_r26_c34_7;
  wire [7:0] t_r26_c34_8;
  wire [7:0] t_r26_c34_9;
  wire [7:0] t_r26_c34_10;
  wire [7:0] t_r26_c34_11;
  wire [7:0] t_r26_c34_12;
  wire [7:0] t_r26_c35_0;
  wire [7:0] t_r26_c35_1;
  wire [7:0] t_r26_c35_2;
  wire [7:0] t_r26_c35_3;
  wire [7:0] t_r26_c35_4;
  wire [7:0] t_r26_c35_5;
  wire [7:0] t_r26_c35_6;
  wire [7:0] t_r26_c35_7;
  wire [7:0] t_r26_c35_8;
  wire [7:0] t_r26_c35_9;
  wire [7:0] t_r26_c35_10;
  wire [7:0] t_r26_c35_11;
  wire [7:0] t_r26_c35_12;
  wire [7:0] t_r26_c36_0;
  wire [7:0] t_r26_c36_1;
  wire [7:0] t_r26_c36_2;
  wire [7:0] t_r26_c36_3;
  wire [7:0] t_r26_c36_4;
  wire [7:0] t_r26_c36_5;
  wire [7:0] t_r26_c36_6;
  wire [7:0] t_r26_c36_7;
  wire [7:0] t_r26_c36_8;
  wire [7:0] t_r26_c36_9;
  wire [7:0] t_r26_c36_10;
  wire [7:0] t_r26_c36_11;
  wire [7:0] t_r26_c36_12;
  wire [7:0] t_r26_c37_0;
  wire [7:0] t_r26_c37_1;
  wire [7:0] t_r26_c37_2;
  wire [7:0] t_r26_c37_3;
  wire [7:0] t_r26_c37_4;
  wire [7:0] t_r26_c37_5;
  wire [7:0] t_r26_c37_6;
  wire [7:0] t_r26_c37_7;
  wire [7:0] t_r26_c37_8;
  wire [7:0] t_r26_c37_9;
  wire [7:0] t_r26_c37_10;
  wire [7:0] t_r26_c37_11;
  wire [7:0] t_r26_c37_12;
  wire [7:0] t_r26_c38_0;
  wire [7:0] t_r26_c38_1;
  wire [7:0] t_r26_c38_2;
  wire [7:0] t_r26_c38_3;
  wire [7:0] t_r26_c38_4;
  wire [7:0] t_r26_c38_5;
  wire [7:0] t_r26_c38_6;
  wire [7:0] t_r26_c38_7;
  wire [7:0] t_r26_c38_8;
  wire [7:0] t_r26_c38_9;
  wire [7:0] t_r26_c38_10;
  wire [7:0] t_r26_c38_11;
  wire [7:0] t_r26_c38_12;
  wire [7:0] t_r26_c39_0;
  wire [7:0] t_r26_c39_1;
  wire [7:0] t_r26_c39_2;
  wire [7:0] t_r26_c39_3;
  wire [7:0] t_r26_c39_4;
  wire [7:0] t_r26_c39_5;
  wire [7:0] t_r26_c39_6;
  wire [7:0] t_r26_c39_7;
  wire [7:0] t_r26_c39_8;
  wire [7:0] t_r26_c39_9;
  wire [7:0] t_r26_c39_10;
  wire [7:0] t_r26_c39_11;
  wire [7:0] t_r26_c39_12;
  wire [7:0] t_r26_c40_0;
  wire [7:0] t_r26_c40_1;
  wire [7:0] t_r26_c40_2;
  wire [7:0] t_r26_c40_3;
  wire [7:0] t_r26_c40_4;
  wire [7:0] t_r26_c40_5;
  wire [7:0] t_r26_c40_6;
  wire [7:0] t_r26_c40_7;
  wire [7:0] t_r26_c40_8;
  wire [7:0] t_r26_c40_9;
  wire [7:0] t_r26_c40_10;
  wire [7:0] t_r26_c40_11;
  wire [7:0] t_r26_c40_12;
  wire [7:0] t_r26_c41_0;
  wire [7:0] t_r26_c41_1;
  wire [7:0] t_r26_c41_2;
  wire [7:0] t_r26_c41_3;
  wire [7:0] t_r26_c41_4;
  wire [7:0] t_r26_c41_5;
  wire [7:0] t_r26_c41_6;
  wire [7:0] t_r26_c41_7;
  wire [7:0] t_r26_c41_8;
  wire [7:0] t_r26_c41_9;
  wire [7:0] t_r26_c41_10;
  wire [7:0] t_r26_c41_11;
  wire [7:0] t_r26_c41_12;
  wire [7:0] t_r26_c42_0;
  wire [7:0] t_r26_c42_1;
  wire [7:0] t_r26_c42_2;
  wire [7:0] t_r26_c42_3;
  wire [7:0] t_r26_c42_4;
  wire [7:0] t_r26_c42_5;
  wire [7:0] t_r26_c42_6;
  wire [7:0] t_r26_c42_7;
  wire [7:0] t_r26_c42_8;
  wire [7:0] t_r26_c42_9;
  wire [7:0] t_r26_c42_10;
  wire [7:0] t_r26_c42_11;
  wire [7:0] t_r26_c42_12;
  wire [7:0] t_r26_c43_0;
  wire [7:0] t_r26_c43_1;
  wire [7:0] t_r26_c43_2;
  wire [7:0] t_r26_c43_3;
  wire [7:0] t_r26_c43_4;
  wire [7:0] t_r26_c43_5;
  wire [7:0] t_r26_c43_6;
  wire [7:0] t_r26_c43_7;
  wire [7:0] t_r26_c43_8;
  wire [7:0] t_r26_c43_9;
  wire [7:0] t_r26_c43_10;
  wire [7:0] t_r26_c43_11;
  wire [7:0] t_r26_c43_12;
  wire [7:0] t_r26_c44_0;
  wire [7:0] t_r26_c44_1;
  wire [7:0] t_r26_c44_2;
  wire [7:0] t_r26_c44_3;
  wire [7:0] t_r26_c44_4;
  wire [7:0] t_r26_c44_5;
  wire [7:0] t_r26_c44_6;
  wire [7:0] t_r26_c44_7;
  wire [7:0] t_r26_c44_8;
  wire [7:0] t_r26_c44_9;
  wire [7:0] t_r26_c44_10;
  wire [7:0] t_r26_c44_11;
  wire [7:0] t_r26_c44_12;
  wire [7:0] t_r26_c45_0;
  wire [7:0] t_r26_c45_1;
  wire [7:0] t_r26_c45_2;
  wire [7:0] t_r26_c45_3;
  wire [7:0] t_r26_c45_4;
  wire [7:0] t_r26_c45_5;
  wire [7:0] t_r26_c45_6;
  wire [7:0] t_r26_c45_7;
  wire [7:0] t_r26_c45_8;
  wire [7:0] t_r26_c45_9;
  wire [7:0] t_r26_c45_10;
  wire [7:0] t_r26_c45_11;
  wire [7:0] t_r26_c45_12;
  wire [7:0] t_r26_c46_0;
  wire [7:0] t_r26_c46_1;
  wire [7:0] t_r26_c46_2;
  wire [7:0] t_r26_c46_3;
  wire [7:0] t_r26_c46_4;
  wire [7:0] t_r26_c46_5;
  wire [7:0] t_r26_c46_6;
  wire [7:0] t_r26_c46_7;
  wire [7:0] t_r26_c46_8;
  wire [7:0] t_r26_c46_9;
  wire [7:0] t_r26_c46_10;
  wire [7:0] t_r26_c46_11;
  wire [7:0] t_r26_c46_12;
  wire [7:0] t_r26_c47_0;
  wire [7:0] t_r26_c47_1;
  wire [7:0] t_r26_c47_2;
  wire [7:0] t_r26_c47_3;
  wire [7:0] t_r26_c47_4;
  wire [7:0] t_r26_c47_5;
  wire [7:0] t_r26_c47_6;
  wire [7:0] t_r26_c47_7;
  wire [7:0] t_r26_c47_8;
  wire [7:0] t_r26_c47_9;
  wire [7:0] t_r26_c47_10;
  wire [7:0] t_r26_c47_11;
  wire [7:0] t_r26_c47_12;
  wire [7:0] t_r26_c48_0;
  wire [7:0] t_r26_c48_1;
  wire [7:0] t_r26_c48_2;
  wire [7:0] t_r26_c48_3;
  wire [7:0] t_r26_c48_4;
  wire [7:0] t_r26_c48_5;
  wire [7:0] t_r26_c48_6;
  wire [7:0] t_r26_c48_7;
  wire [7:0] t_r26_c48_8;
  wire [7:0] t_r26_c48_9;
  wire [7:0] t_r26_c48_10;
  wire [7:0] t_r26_c48_11;
  wire [7:0] t_r26_c48_12;
  wire [7:0] t_r26_c49_0;
  wire [7:0] t_r26_c49_1;
  wire [7:0] t_r26_c49_2;
  wire [7:0] t_r26_c49_3;
  wire [7:0] t_r26_c49_4;
  wire [7:0] t_r26_c49_5;
  wire [7:0] t_r26_c49_6;
  wire [7:0] t_r26_c49_7;
  wire [7:0] t_r26_c49_8;
  wire [7:0] t_r26_c49_9;
  wire [7:0] t_r26_c49_10;
  wire [7:0] t_r26_c49_11;
  wire [7:0] t_r26_c49_12;
  wire [7:0] t_r26_c50_0;
  wire [7:0] t_r26_c50_1;
  wire [7:0] t_r26_c50_2;
  wire [7:0] t_r26_c50_3;
  wire [7:0] t_r26_c50_4;
  wire [7:0] t_r26_c50_5;
  wire [7:0] t_r26_c50_6;
  wire [7:0] t_r26_c50_7;
  wire [7:0] t_r26_c50_8;
  wire [7:0] t_r26_c50_9;
  wire [7:0] t_r26_c50_10;
  wire [7:0] t_r26_c50_11;
  wire [7:0] t_r26_c50_12;
  wire [7:0] t_r26_c51_0;
  wire [7:0] t_r26_c51_1;
  wire [7:0] t_r26_c51_2;
  wire [7:0] t_r26_c51_3;
  wire [7:0] t_r26_c51_4;
  wire [7:0] t_r26_c51_5;
  wire [7:0] t_r26_c51_6;
  wire [7:0] t_r26_c51_7;
  wire [7:0] t_r26_c51_8;
  wire [7:0] t_r26_c51_9;
  wire [7:0] t_r26_c51_10;
  wire [7:0] t_r26_c51_11;
  wire [7:0] t_r26_c51_12;
  wire [7:0] t_r26_c52_0;
  wire [7:0] t_r26_c52_1;
  wire [7:0] t_r26_c52_2;
  wire [7:0] t_r26_c52_3;
  wire [7:0] t_r26_c52_4;
  wire [7:0] t_r26_c52_5;
  wire [7:0] t_r26_c52_6;
  wire [7:0] t_r26_c52_7;
  wire [7:0] t_r26_c52_8;
  wire [7:0] t_r26_c52_9;
  wire [7:0] t_r26_c52_10;
  wire [7:0] t_r26_c52_11;
  wire [7:0] t_r26_c52_12;
  wire [7:0] t_r26_c53_0;
  wire [7:0] t_r26_c53_1;
  wire [7:0] t_r26_c53_2;
  wire [7:0] t_r26_c53_3;
  wire [7:0] t_r26_c53_4;
  wire [7:0] t_r26_c53_5;
  wire [7:0] t_r26_c53_6;
  wire [7:0] t_r26_c53_7;
  wire [7:0] t_r26_c53_8;
  wire [7:0] t_r26_c53_9;
  wire [7:0] t_r26_c53_10;
  wire [7:0] t_r26_c53_11;
  wire [7:0] t_r26_c53_12;
  wire [7:0] t_r26_c54_0;
  wire [7:0] t_r26_c54_1;
  wire [7:0] t_r26_c54_2;
  wire [7:0] t_r26_c54_3;
  wire [7:0] t_r26_c54_4;
  wire [7:0] t_r26_c54_5;
  wire [7:0] t_r26_c54_6;
  wire [7:0] t_r26_c54_7;
  wire [7:0] t_r26_c54_8;
  wire [7:0] t_r26_c54_9;
  wire [7:0] t_r26_c54_10;
  wire [7:0] t_r26_c54_11;
  wire [7:0] t_r26_c54_12;
  wire [7:0] t_r26_c55_0;
  wire [7:0] t_r26_c55_1;
  wire [7:0] t_r26_c55_2;
  wire [7:0] t_r26_c55_3;
  wire [7:0] t_r26_c55_4;
  wire [7:0] t_r26_c55_5;
  wire [7:0] t_r26_c55_6;
  wire [7:0] t_r26_c55_7;
  wire [7:0] t_r26_c55_8;
  wire [7:0] t_r26_c55_9;
  wire [7:0] t_r26_c55_10;
  wire [7:0] t_r26_c55_11;
  wire [7:0] t_r26_c55_12;
  wire [7:0] t_r26_c56_0;
  wire [7:0] t_r26_c56_1;
  wire [7:0] t_r26_c56_2;
  wire [7:0] t_r26_c56_3;
  wire [7:0] t_r26_c56_4;
  wire [7:0] t_r26_c56_5;
  wire [7:0] t_r26_c56_6;
  wire [7:0] t_r26_c56_7;
  wire [7:0] t_r26_c56_8;
  wire [7:0] t_r26_c56_9;
  wire [7:0] t_r26_c56_10;
  wire [7:0] t_r26_c56_11;
  wire [7:0] t_r26_c56_12;
  wire [7:0] t_r26_c57_0;
  wire [7:0] t_r26_c57_1;
  wire [7:0] t_r26_c57_2;
  wire [7:0] t_r26_c57_3;
  wire [7:0] t_r26_c57_4;
  wire [7:0] t_r26_c57_5;
  wire [7:0] t_r26_c57_6;
  wire [7:0] t_r26_c57_7;
  wire [7:0] t_r26_c57_8;
  wire [7:0] t_r26_c57_9;
  wire [7:0] t_r26_c57_10;
  wire [7:0] t_r26_c57_11;
  wire [7:0] t_r26_c57_12;
  wire [7:0] t_r26_c58_0;
  wire [7:0] t_r26_c58_1;
  wire [7:0] t_r26_c58_2;
  wire [7:0] t_r26_c58_3;
  wire [7:0] t_r26_c58_4;
  wire [7:0] t_r26_c58_5;
  wire [7:0] t_r26_c58_6;
  wire [7:0] t_r26_c58_7;
  wire [7:0] t_r26_c58_8;
  wire [7:0] t_r26_c58_9;
  wire [7:0] t_r26_c58_10;
  wire [7:0] t_r26_c58_11;
  wire [7:0] t_r26_c58_12;
  wire [7:0] t_r26_c59_0;
  wire [7:0] t_r26_c59_1;
  wire [7:0] t_r26_c59_2;
  wire [7:0] t_r26_c59_3;
  wire [7:0] t_r26_c59_4;
  wire [7:0] t_r26_c59_5;
  wire [7:0] t_r26_c59_6;
  wire [7:0] t_r26_c59_7;
  wire [7:0] t_r26_c59_8;
  wire [7:0] t_r26_c59_9;
  wire [7:0] t_r26_c59_10;
  wire [7:0] t_r26_c59_11;
  wire [7:0] t_r26_c59_12;
  wire [7:0] t_r26_c60_0;
  wire [7:0] t_r26_c60_1;
  wire [7:0] t_r26_c60_2;
  wire [7:0] t_r26_c60_3;
  wire [7:0] t_r26_c60_4;
  wire [7:0] t_r26_c60_5;
  wire [7:0] t_r26_c60_6;
  wire [7:0] t_r26_c60_7;
  wire [7:0] t_r26_c60_8;
  wire [7:0] t_r26_c60_9;
  wire [7:0] t_r26_c60_10;
  wire [7:0] t_r26_c60_11;
  wire [7:0] t_r26_c60_12;
  wire [7:0] t_r26_c61_0;
  wire [7:0] t_r26_c61_1;
  wire [7:0] t_r26_c61_2;
  wire [7:0] t_r26_c61_3;
  wire [7:0] t_r26_c61_4;
  wire [7:0] t_r26_c61_5;
  wire [7:0] t_r26_c61_6;
  wire [7:0] t_r26_c61_7;
  wire [7:0] t_r26_c61_8;
  wire [7:0] t_r26_c61_9;
  wire [7:0] t_r26_c61_10;
  wire [7:0] t_r26_c61_11;
  wire [7:0] t_r26_c61_12;
  wire [7:0] t_r26_c62_0;
  wire [7:0] t_r26_c62_1;
  wire [7:0] t_r26_c62_2;
  wire [7:0] t_r26_c62_3;
  wire [7:0] t_r26_c62_4;
  wire [7:0] t_r26_c62_5;
  wire [7:0] t_r26_c62_6;
  wire [7:0] t_r26_c62_7;
  wire [7:0] t_r26_c62_8;
  wire [7:0] t_r26_c62_9;
  wire [7:0] t_r26_c62_10;
  wire [7:0] t_r26_c62_11;
  wire [7:0] t_r26_c62_12;
  wire [7:0] t_r26_c63_0;
  wire [7:0] t_r26_c63_1;
  wire [7:0] t_r26_c63_2;
  wire [7:0] t_r26_c63_3;
  wire [7:0] t_r26_c63_4;
  wire [7:0] t_r26_c63_5;
  wire [7:0] t_r26_c63_6;
  wire [7:0] t_r26_c63_7;
  wire [7:0] t_r26_c63_8;
  wire [7:0] t_r26_c63_9;
  wire [7:0] t_r26_c63_10;
  wire [7:0] t_r26_c63_11;
  wire [7:0] t_r26_c63_12;
  wire [7:0] t_r26_c64_0;
  wire [7:0] t_r26_c64_1;
  wire [7:0] t_r26_c64_2;
  wire [7:0] t_r26_c64_3;
  wire [7:0] t_r26_c64_4;
  wire [7:0] t_r26_c64_5;
  wire [7:0] t_r26_c64_6;
  wire [7:0] t_r26_c64_7;
  wire [7:0] t_r26_c64_8;
  wire [7:0] t_r26_c64_9;
  wire [7:0] t_r26_c64_10;
  wire [7:0] t_r26_c64_11;
  wire [7:0] t_r26_c64_12;
  wire [7:0] t_r26_c65_0;
  wire [7:0] t_r26_c65_1;
  wire [7:0] t_r26_c65_2;
  wire [7:0] t_r26_c65_3;
  wire [7:0] t_r26_c65_4;
  wire [7:0] t_r26_c65_5;
  wire [7:0] t_r26_c65_6;
  wire [7:0] t_r26_c65_7;
  wire [7:0] t_r26_c65_8;
  wire [7:0] t_r26_c65_9;
  wire [7:0] t_r26_c65_10;
  wire [7:0] t_r26_c65_11;
  wire [7:0] t_r26_c65_12;
  wire [7:0] t_r27_c0_0;
  wire [7:0] t_r27_c0_1;
  wire [7:0] t_r27_c0_2;
  wire [7:0] t_r27_c0_3;
  wire [7:0] t_r27_c0_4;
  wire [7:0] t_r27_c0_5;
  wire [7:0] t_r27_c0_6;
  wire [7:0] t_r27_c0_7;
  wire [7:0] t_r27_c0_8;
  wire [7:0] t_r27_c0_9;
  wire [7:0] t_r27_c0_10;
  wire [7:0] t_r27_c0_11;
  wire [7:0] t_r27_c0_12;
  wire [7:0] t_r27_c1_0;
  wire [7:0] t_r27_c1_1;
  wire [7:0] t_r27_c1_2;
  wire [7:0] t_r27_c1_3;
  wire [7:0] t_r27_c1_4;
  wire [7:0] t_r27_c1_5;
  wire [7:0] t_r27_c1_6;
  wire [7:0] t_r27_c1_7;
  wire [7:0] t_r27_c1_8;
  wire [7:0] t_r27_c1_9;
  wire [7:0] t_r27_c1_10;
  wire [7:0] t_r27_c1_11;
  wire [7:0] t_r27_c1_12;
  wire [7:0] t_r27_c2_0;
  wire [7:0] t_r27_c2_1;
  wire [7:0] t_r27_c2_2;
  wire [7:0] t_r27_c2_3;
  wire [7:0] t_r27_c2_4;
  wire [7:0] t_r27_c2_5;
  wire [7:0] t_r27_c2_6;
  wire [7:0] t_r27_c2_7;
  wire [7:0] t_r27_c2_8;
  wire [7:0] t_r27_c2_9;
  wire [7:0] t_r27_c2_10;
  wire [7:0] t_r27_c2_11;
  wire [7:0] t_r27_c2_12;
  wire [7:0] t_r27_c3_0;
  wire [7:0] t_r27_c3_1;
  wire [7:0] t_r27_c3_2;
  wire [7:0] t_r27_c3_3;
  wire [7:0] t_r27_c3_4;
  wire [7:0] t_r27_c3_5;
  wire [7:0] t_r27_c3_6;
  wire [7:0] t_r27_c3_7;
  wire [7:0] t_r27_c3_8;
  wire [7:0] t_r27_c3_9;
  wire [7:0] t_r27_c3_10;
  wire [7:0] t_r27_c3_11;
  wire [7:0] t_r27_c3_12;
  wire [7:0] t_r27_c4_0;
  wire [7:0] t_r27_c4_1;
  wire [7:0] t_r27_c4_2;
  wire [7:0] t_r27_c4_3;
  wire [7:0] t_r27_c4_4;
  wire [7:0] t_r27_c4_5;
  wire [7:0] t_r27_c4_6;
  wire [7:0] t_r27_c4_7;
  wire [7:0] t_r27_c4_8;
  wire [7:0] t_r27_c4_9;
  wire [7:0] t_r27_c4_10;
  wire [7:0] t_r27_c4_11;
  wire [7:0] t_r27_c4_12;
  wire [7:0] t_r27_c5_0;
  wire [7:0] t_r27_c5_1;
  wire [7:0] t_r27_c5_2;
  wire [7:0] t_r27_c5_3;
  wire [7:0] t_r27_c5_4;
  wire [7:0] t_r27_c5_5;
  wire [7:0] t_r27_c5_6;
  wire [7:0] t_r27_c5_7;
  wire [7:0] t_r27_c5_8;
  wire [7:0] t_r27_c5_9;
  wire [7:0] t_r27_c5_10;
  wire [7:0] t_r27_c5_11;
  wire [7:0] t_r27_c5_12;
  wire [7:0] t_r27_c6_0;
  wire [7:0] t_r27_c6_1;
  wire [7:0] t_r27_c6_2;
  wire [7:0] t_r27_c6_3;
  wire [7:0] t_r27_c6_4;
  wire [7:0] t_r27_c6_5;
  wire [7:0] t_r27_c6_6;
  wire [7:0] t_r27_c6_7;
  wire [7:0] t_r27_c6_8;
  wire [7:0] t_r27_c6_9;
  wire [7:0] t_r27_c6_10;
  wire [7:0] t_r27_c6_11;
  wire [7:0] t_r27_c6_12;
  wire [7:0] t_r27_c7_0;
  wire [7:0] t_r27_c7_1;
  wire [7:0] t_r27_c7_2;
  wire [7:0] t_r27_c7_3;
  wire [7:0] t_r27_c7_4;
  wire [7:0] t_r27_c7_5;
  wire [7:0] t_r27_c7_6;
  wire [7:0] t_r27_c7_7;
  wire [7:0] t_r27_c7_8;
  wire [7:0] t_r27_c7_9;
  wire [7:0] t_r27_c7_10;
  wire [7:0] t_r27_c7_11;
  wire [7:0] t_r27_c7_12;
  wire [7:0] t_r27_c8_0;
  wire [7:0] t_r27_c8_1;
  wire [7:0] t_r27_c8_2;
  wire [7:0] t_r27_c8_3;
  wire [7:0] t_r27_c8_4;
  wire [7:0] t_r27_c8_5;
  wire [7:0] t_r27_c8_6;
  wire [7:0] t_r27_c8_7;
  wire [7:0] t_r27_c8_8;
  wire [7:0] t_r27_c8_9;
  wire [7:0] t_r27_c8_10;
  wire [7:0] t_r27_c8_11;
  wire [7:0] t_r27_c8_12;
  wire [7:0] t_r27_c9_0;
  wire [7:0] t_r27_c9_1;
  wire [7:0] t_r27_c9_2;
  wire [7:0] t_r27_c9_3;
  wire [7:0] t_r27_c9_4;
  wire [7:0] t_r27_c9_5;
  wire [7:0] t_r27_c9_6;
  wire [7:0] t_r27_c9_7;
  wire [7:0] t_r27_c9_8;
  wire [7:0] t_r27_c9_9;
  wire [7:0] t_r27_c9_10;
  wire [7:0] t_r27_c9_11;
  wire [7:0] t_r27_c9_12;
  wire [7:0] t_r27_c10_0;
  wire [7:0] t_r27_c10_1;
  wire [7:0] t_r27_c10_2;
  wire [7:0] t_r27_c10_3;
  wire [7:0] t_r27_c10_4;
  wire [7:0] t_r27_c10_5;
  wire [7:0] t_r27_c10_6;
  wire [7:0] t_r27_c10_7;
  wire [7:0] t_r27_c10_8;
  wire [7:0] t_r27_c10_9;
  wire [7:0] t_r27_c10_10;
  wire [7:0] t_r27_c10_11;
  wire [7:0] t_r27_c10_12;
  wire [7:0] t_r27_c11_0;
  wire [7:0] t_r27_c11_1;
  wire [7:0] t_r27_c11_2;
  wire [7:0] t_r27_c11_3;
  wire [7:0] t_r27_c11_4;
  wire [7:0] t_r27_c11_5;
  wire [7:0] t_r27_c11_6;
  wire [7:0] t_r27_c11_7;
  wire [7:0] t_r27_c11_8;
  wire [7:0] t_r27_c11_9;
  wire [7:0] t_r27_c11_10;
  wire [7:0] t_r27_c11_11;
  wire [7:0] t_r27_c11_12;
  wire [7:0] t_r27_c12_0;
  wire [7:0] t_r27_c12_1;
  wire [7:0] t_r27_c12_2;
  wire [7:0] t_r27_c12_3;
  wire [7:0] t_r27_c12_4;
  wire [7:0] t_r27_c12_5;
  wire [7:0] t_r27_c12_6;
  wire [7:0] t_r27_c12_7;
  wire [7:0] t_r27_c12_8;
  wire [7:0] t_r27_c12_9;
  wire [7:0] t_r27_c12_10;
  wire [7:0] t_r27_c12_11;
  wire [7:0] t_r27_c12_12;
  wire [7:0] t_r27_c13_0;
  wire [7:0] t_r27_c13_1;
  wire [7:0] t_r27_c13_2;
  wire [7:0] t_r27_c13_3;
  wire [7:0] t_r27_c13_4;
  wire [7:0] t_r27_c13_5;
  wire [7:0] t_r27_c13_6;
  wire [7:0] t_r27_c13_7;
  wire [7:0] t_r27_c13_8;
  wire [7:0] t_r27_c13_9;
  wire [7:0] t_r27_c13_10;
  wire [7:0] t_r27_c13_11;
  wire [7:0] t_r27_c13_12;
  wire [7:0] t_r27_c14_0;
  wire [7:0] t_r27_c14_1;
  wire [7:0] t_r27_c14_2;
  wire [7:0] t_r27_c14_3;
  wire [7:0] t_r27_c14_4;
  wire [7:0] t_r27_c14_5;
  wire [7:0] t_r27_c14_6;
  wire [7:0] t_r27_c14_7;
  wire [7:0] t_r27_c14_8;
  wire [7:0] t_r27_c14_9;
  wire [7:0] t_r27_c14_10;
  wire [7:0] t_r27_c14_11;
  wire [7:0] t_r27_c14_12;
  wire [7:0] t_r27_c15_0;
  wire [7:0] t_r27_c15_1;
  wire [7:0] t_r27_c15_2;
  wire [7:0] t_r27_c15_3;
  wire [7:0] t_r27_c15_4;
  wire [7:0] t_r27_c15_5;
  wire [7:0] t_r27_c15_6;
  wire [7:0] t_r27_c15_7;
  wire [7:0] t_r27_c15_8;
  wire [7:0] t_r27_c15_9;
  wire [7:0] t_r27_c15_10;
  wire [7:0] t_r27_c15_11;
  wire [7:0] t_r27_c15_12;
  wire [7:0] t_r27_c16_0;
  wire [7:0] t_r27_c16_1;
  wire [7:0] t_r27_c16_2;
  wire [7:0] t_r27_c16_3;
  wire [7:0] t_r27_c16_4;
  wire [7:0] t_r27_c16_5;
  wire [7:0] t_r27_c16_6;
  wire [7:0] t_r27_c16_7;
  wire [7:0] t_r27_c16_8;
  wire [7:0] t_r27_c16_9;
  wire [7:0] t_r27_c16_10;
  wire [7:0] t_r27_c16_11;
  wire [7:0] t_r27_c16_12;
  wire [7:0] t_r27_c17_0;
  wire [7:0] t_r27_c17_1;
  wire [7:0] t_r27_c17_2;
  wire [7:0] t_r27_c17_3;
  wire [7:0] t_r27_c17_4;
  wire [7:0] t_r27_c17_5;
  wire [7:0] t_r27_c17_6;
  wire [7:0] t_r27_c17_7;
  wire [7:0] t_r27_c17_8;
  wire [7:0] t_r27_c17_9;
  wire [7:0] t_r27_c17_10;
  wire [7:0] t_r27_c17_11;
  wire [7:0] t_r27_c17_12;
  wire [7:0] t_r27_c18_0;
  wire [7:0] t_r27_c18_1;
  wire [7:0] t_r27_c18_2;
  wire [7:0] t_r27_c18_3;
  wire [7:0] t_r27_c18_4;
  wire [7:0] t_r27_c18_5;
  wire [7:0] t_r27_c18_6;
  wire [7:0] t_r27_c18_7;
  wire [7:0] t_r27_c18_8;
  wire [7:0] t_r27_c18_9;
  wire [7:0] t_r27_c18_10;
  wire [7:0] t_r27_c18_11;
  wire [7:0] t_r27_c18_12;
  wire [7:0] t_r27_c19_0;
  wire [7:0] t_r27_c19_1;
  wire [7:0] t_r27_c19_2;
  wire [7:0] t_r27_c19_3;
  wire [7:0] t_r27_c19_4;
  wire [7:0] t_r27_c19_5;
  wire [7:0] t_r27_c19_6;
  wire [7:0] t_r27_c19_7;
  wire [7:0] t_r27_c19_8;
  wire [7:0] t_r27_c19_9;
  wire [7:0] t_r27_c19_10;
  wire [7:0] t_r27_c19_11;
  wire [7:0] t_r27_c19_12;
  wire [7:0] t_r27_c20_0;
  wire [7:0] t_r27_c20_1;
  wire [7:0] t_r27_c20_2;
  wire [7:0] t_r27_c20_3;
  wire [7:0] t_r27_c20_4;
  wire [7:0] t_r27_c20_5;
  wire [7:0] t_r27_c20_6;
  wire [7:0] t_r27_c20_7;
  wire [7:0] t_r27_c20_8;
  wire [7:0] t_r27_c20_9;
  wire [7:0] t_r27_c20_10;
  wire [7:0] t_r27_c20_11;
  wire [7:0] t_r27_c20_12;
  wire [7:0] t_r27_c21_0;
  wire [7:0] t_r27_c21_1;
  wire [7:0] t_r27_c21_2;
  wire [7:0] t_r27_c21_3;
  wire [7:0] t_r27_c21_4;
  wire [7:0] t_r27_c21_5;
  wire [7:0] t_r27_c21_6;
  wire [7:0] t_r27_c21_7;
  wire [7:0] t_r27_c21_8;
  wire [7:0] t_r27_c21_9;
  wire [7:0] t_r27_c21_10;
  wire [7:0] t_r27_c21_11;
  wire [7:0] t_r27_c21_12;
  wire [7:0] t_r27_c22_0;
  wire [7:0] t_r27_c22_1;
  wire [7:0] t_r27_c22_2;
  wire [7:0] t_r27_c22_3;
  wire [7:0] t_r27_c22_4;
  wire [7:0] t_r27_c22_5;
  wire [7:0] t_r27_c22_6;
  wire [7:0] t_r27_c22_7;
  wire [7:0] t_r27_c22_8;
  wire [7:0] t_r27_c22_9;
  wire [7:0] t_r27_c22_10;
  wire [7:0] t_r27_c22_11;
  wire [7:0] t_r27_c22_12;
  wire [7:0] t_r27_c23_0;
  wire [7:0] t_r27_c23_1;
  wire [7:0] t_r27_c23_2;
  wire [7:0] t_r27_c23_3;
  wire [7:0] t_r27_c23_4;
  wire [7:0] t_r27_c23_5;
  wire [7:0] t_r27_c23_6;
  wire [7:0] t_r27_c23_7;
  wire [7:0] t_r27_c23_8;
  wire [7:0] t_r27_c23_9;
  wire [7:0] t_r27_c23_10;
  wire [7:0] t_r27_c23_11;
  wire [7:0] t_r27_c23_12;
  wire [7:0] t_r27_c24_0;
  wire [7:0] t_r27_c24_1;
  wire [7:0] t_r27_c24_2;
  wire [7:0] t_r27_c24_3;
  wire [7:0] t_r27_c24_4;
  wire [7:0] t_r27_c24_5;
  wire [7:0] t_r27_c24_6;
  wire [7:0] t_r27_c24_7;
  wire [7:0] t_r27_c24_8;
  wire [7:0] t_r27_c24_9;
  wire [7:0] t_r27_c24_10;
  wire [7:0] t_r27_c24_11;
  wire [7:0] t_r27_c24_12;
  wire [7:0] t_r27_c25_0;
  wire [7:0] t_r27_c25_1;
  wire [7:0] t_r27_c25_2;
  wire [7:0] t_r27_c25_3;
  wire [7:0] t_r27_c25_4;
  wire [7:0] t_r27_c25_5;
  wire [7:0] t_r27_c25_6;
  wire [7:0] t_r27_c25_7;
  wire [7:0] t_r27_c25_8;
  wire [7:0] t_r27_c25_9;
  wire [7:0] t_r27_c25_10;
  wire [7:0] t_r27_c25_11;
  wire [7:0] t_r27_c25_12;
  wire [7:0] t_r27_c26_0;
  wire [7:0] t_r27_c26_1;
  wire [7:0] t_r27_c26_2;
  wire [7:0] t_r27_c26_3;
  wire [7:0] t_r27_c26_4;
  wire [7:0] t_r27_c26_5;
  wire [7:0] t_r27_c26_6;
  wire [7:0] t_r27_c26_7;
  wire [7:0] t_r27_c26_8;
  wire [7:0] t_r27_c26_9;
  wire [7:0] t_r27_c26_10;
  wire [7:0] t_r27_c26_11;
  wire [7:0] t_r27_c26_12;
  wire [7:0] t_r27_c27_0;
  wire [7:0] t_r27_c27_1;
  wire [7:0] t_r27_c27_2;
  wire [7:0] t_r27_c27_3;
  wire [7:0] t_r27_c27_4;
  wire [7:0] t_r27_c27_5;
  wire [7:0] t_r27_c27_6;
  wire [7:0] t_r27_c27_7;
  wire [7:0] t_r27_c27_8;
  wire [7:0] t_r27_c27_9;
  wire [7:0] t_r27_c27_10;
  wire [7:0] t_r27_c27_11;
  wire [7:0] t_r27_c27_12;
  wire [7:0] t_r27_c28_0;
  wire [7:0] t_r27_c28_1;
  wire [7:0] t_r27_c28_2;
  wire [7:0] t_r27_c28_3;
  wire [7:0] t_r27_c28_4;
  wire [7:0] t_r27_c28_5;
  wire [7:0] t_r27_c28_6;
  wire [7:0] t_r27_c28_7;
  wire [7:0] t_r27_c28_8;
  wire [7:0] t_r27_c28_9;
  wire [7:0] t_r27_c28_10;
  wire [7:0] t_r27_c28_11;
  wire [7:0] t_r27_c28_12;
  wire [7:0] t_r27_c29_0;
  wire [7:0] t_r27_c29_1;
  wire [7:0] t_r27_c29_2;
  wire [7:0] t_r27_c29_3;
  wire [7:0] t_r27_c29_4;
  wire [7:0] t_r27_c29_5;
  wire [7:0] t_r27_c29_6;
  wire [7:0] t_r27_c29_7;
  wire [7:0] t_r27_c29_8;
  wire [7:0] t_r27_c29_9;
  wire [7:0] t_r27_c29_10;
  wire [7:0] t_r27_c29_11;
  wire [7:0] t_r27_c29_12;
  wire [7:0] t_r27_c30_0;
  wire [7:0] t_r27_c30_1;
  wire [7:0] t_r27_c30_2;
  wire [7:0] t_r27_c30_3;
  wire [7:0] t_r27_c30_4;
  wire [7:0] t_r27_c30_5;
  wire [7:0] t_r27_c30_6;
  wire [7:0] t_r27_c30_7;
  wire [7:0] t_r27_c30_8;
  wire [7:0] t_r27_c30_9;
  wire [7:0] t_r27_c30_10;
  wire [7:0] t_r27_c30_11;
  wire [7:0] t_r27_c30_12;
  wire [7:0] t_r27_c31_0;
  wire [7:0] t_r27_c31_1;
  wire [7:0] t_r27_c31_2;
  wire [7:0] t_r27_c31_3;
  wire [7:0] t_r27_c31_4;
  wire [7:0] t_r27_c31_5;
  wire [7:0] t_r27_c31_6;
  wire [7:0] t_r27_c31_7;
  wire [7:0] t_r27_c31_8;
  wire [7:0] t_r27_c31_9;
  wire [7:0] t_r27_c31_10;
  wire [7:0] t_r27_c31_11;
  wire [7:0] t_r27_c31_12;
  wire [7:0] t_r27_c32_0;
  wire [7:0] t_r27_c32_1;
  wire [7:0] t_r27_c32_2;
  wire [7:0] t_r27_c32_3;
  wire [7:0] t_r27_c32_4;
  wire [7:0] t_r27_c32_5;
  wire [7:0] t_r27_c32_6;
  wire [7:0] t_r27_c32_7;
  wire [7:0] t_r27_c32_8;
  wire [7:0] t_r27_c32_9;
  wire [7:0] t_r27_c32_10;
  wire [7:0] t_r27_c32_11;
  wire [7:0] t_r27_c32_12;
  wire [7:0] t_r27_c33_0;
  wire [7:0] t_r27_c33_1;
  wire [7:0] t_r27_c33_2;
  wire [7:0] t_r27_c33_3;
  wire [7:0] t_r27_c33_4;
  wire [7:0] t_r27_c33_5;
  wire [7:0] t_r27_c33_6;
  wire [7:0] t_r27_c33_7;
  wire [7:0] t_r27_c33_8;
  wire [7:0] t_r27_c33_9;
  wire [7:0] t_r27_c33_10;
  wire [7:0] t_r27_c33_11;
  wire [7:0] t_r27_c33_12;
  wire [7:0] t_r27_c34_0;
  wire [7:0] t_r27_c34_1;
  wire [7:0] t_r27_c34_2;
  wire [7:0] t_r27_c34_3;
  wire [7:0] t_r27_c34_4;
  wire [7:0] t_r27_c34_5;
  wire [7:0] t_r27_c34_6;
  wire [7:0] t_r27_c34_7;
  wire [7:0] t_r27_c34_8;
  wire [7:0] t_r27_c34_9;
  wire [7:0] t_r27_c34_10;
  wire [7:0] t_r27_c34_11;
  wire [7:0] t_r27_c34_12;
  wire [7:0] t_r27_c35_0;
  wire [7:0] t_r27_c35_1;
  wire [7:0] t_r27_c35_2;
  wire [7:0] t_r27_c35_3;
  wire [7:0] t_r27_c35_4;
  wire [7:0] t_r27_c35_5;
  wire [7:0] t_r27_c35_6;
  wire [7:0] t_r27_c35_7;
  wire [7:0] t_r27_c35_8;
  wire [7:0] t_r27_c35_9;
  wire [7:0] t_r27_c35_10;
  wire [7:0] t_r27_c35_11;
  wire [7:0] t_r27_c35_12;
  wire [7:0] t_r27_c36_0;
  wire [7:0] t_r27_c36_1;
  wire [7:0] t_r27_c36_2;
  wire [7:0] t_r27_c36_3;
  wire [7:0] t_r27_c36_4;
  wire [7:0] t_r27_c36_5;
  wire [7:0] t_r27_c36_6;
  wire [7:0] t_r27_c36_7;
  wire [7:0] t_r27_c36_8;
  wire [7:0] t_r27_c36_9;
  wire [7:0] t_r27_c36_10;
  wire [7:0] t_r27_c36_11;
  wire [7:0] t_r27_c36_12;
  wire [7:0] t_r27_c37_0;
  wire [7:0] t_r27_c37_1;
  wire [7:0] t_r27_c37_2;
  wire [7:0] t_r27_c37_3;
  wire [7:0] t_r27_c37_4;
  wire [7:0] t_r27_c37_5;
  wire [7:0] t_r27_c37_6;
  wire [7:0] t_r27_c37_7;
  wire [7:0] t_r27_c37_8;
  wire [7:0] t_r27_c37_9;
  wire [7:0] t_r27_c37_10;
  wire [7:0] t_r27_c37_11;
  wire [7:0] t_r27_c37_12;
  wire [7:0] t_r27_c38_0;
  wire [7:0] t_r27_c38_1;
  wire [7:0] t_r27_c38_2;
  wire [7:0] t_r27_c38_3;
  wire [7:0] t_r27_c38_4;
  wire [7:0] t_r27_c38_5;
  wire [7:0] t_r27_c38_6;
  wire [7:0] t_r27_c38_7;
  wire [7:0] t_r27_c38_8;
  wire [7:0] t_r27_c38_9;
  wire [7:0] t_r27_c38_10;
  wire [7:0] t_r27_c38_11;
  wire [7:0] t_r27_c38_12;
  wire [7:0] t_r27_c39_0;
  wire [7:0] t_r27_c39_1;
  wire [7:0] t_r27_c39_2;
  wire [7:0] t_r27_c39_3;
  wire [7:0] t_r27_c39_4;
  wire [7:0] t_r27_c39_5;
  wire [7:0] t_r27_c39_6;
  wire [7:0] t_r27_c39_7;
  wire [7:0] t_r27_c39_8;
  wire [7:0] t_r27_c39_9;
  wire [7:0] t_r27_c39_10;
  wire [7:0] t_r27_c39_11;
  wire [7:0] t_r27_c39_12;
  wire [7:0] t_r27_c40_0;
  wire [7:0] t_r27_c40_1;
  wire [7:0] t_r27_c40_2;
  wire [7:0] t_r27_c40_3;
  wire [7:0] t_r27_c40_4;
  wire [7:0] t_r27_c40_5;
  wire [7:0] t_r27_c40_6;
  wire [7:0] t_r27_c40_7;
  wire [7:0] t_r27_c40_8;
  wire [7:0] t_r27_c40_9;
  wire [7:0] t_r27_c40_10;
  wire [7:0] t_r27_c40_11;
  wire [7:0] t_r27_c40_12;
  wire [7:0] t_r27_c41_0;
  wire [7:0] t_r27_c41_1;
  wire [7:0] t_r27_c41_2;
  wire [7:0] t_r27_c41_3;
  wire [7:0] t_r27_c41_4;
  wire [7:0] t_r27_c41_5;
  wire [7:0] t_r27_c41_6;
  wire [7:0] t_r27_c41_7;
  wire [7:0] t_r27_c41_8;
  wire [7:0] t_r27_c41_9;
  wire [7:0] t_r27_c41_10;
  wire [7:0] t_r27_c41_11;
  wire [7:0] t_r27_c41_12;
  wire [7:0] t_r27_c42_0;
  wire [7:0] t_r27_c42_1;
  wire [7:0] t_r27_c42_2;
  wire [7:0] t_r27_c42_3;
  wire [7:0] t_r27_c42_4;
  wire [7:0] t_r27_c42_5;
  wire [7:0] t_r27_c42_6;
  wire [7:0] t_r27_c42_7;
  wire [7:0] t_r27_c42_8;
  wire [7:0] t_r27_c42_9;
  wire [7:0] t_r27_c42_10;
  wire [7:0] t_r27_c42_11;
  wire [7:0] t_r27_c42_12;
  wire [7:0] t_r27_c43_0;
  wire [7:0] t_r27_c43_1;
  wire [7:0] t_r27_c43_2;
  wire [7:0] t_r27_c43_3;
  wire [7:0] t_r27_c43_4;
  wire [7:0] t_r27_c43_5;
  wire [7:0] t_r27_c43_6;
  wire [7:0] t_r27_c43_7;
  wire [7:0] t_r27_c43_8;
  wire [7:0] t_r27_c43_9;
  wire [7:0] t_r27_c43_10;
  wire [7:0] t_r27_c43_11;
  wire [7:0] t_r27_c43_12;
  wire [7:0] t_r27_c44_0;
  wire [7:0] t_r27_c44_1;
  wire [7:0] t_r27_c44_2;
  wire [7:0] t_r27_c44_3;
  wire [7:0] t_r27_c44_4;
  wire [7:0] t_r27_c44_5;
  wire [7:0] t_r27_c44_6;
  wire [7:0] t_r27_c44_7;
  wire [7:0] t_r27_c44_8;
  wire [7:0] t_r27_c44_9;
  wire [7:0] t_r27_c44_10;
  wire [7:0] t_r27_c44_11;
  wire [7:0] t_r27_c44_12;
  wire [7:0] t_r27_c45_0;
  wire [7:0] t_r27_c45_1;
  wire [7:0] t_r27_c45_2;
  wire [7:0] t_r27_c45_3;
  wire [7:0] t_r27_c45_4;
  wire [7:0] t_r27_c45_5;
  wire [7:0] t_r27_c45_6;
  wire [7:0] t_r27_c45_7;
  wire [7:0] t_r27_c45_8;
  wire [7:0] t_r27_c45_9;
  wire [7:0] t_r27_c45_10;
  wire [7:0] t_r27_c45_11;
  wire [7:0] t_r27_c45_12;
  wire [7:0] t_r27_c46_0;
  wire [7:0] t_r27_c46_1;
  wire [7:0] t_r27_c46_2;
  wire [7:0] t_r27_c46_3;
  wire [7:0] t_r27_c46_4;
  wire [7:0] t_r27_c46_5;
  wire [7:0] t_r27_c46_6;
  wire [7:0] t_r27_c46_7;
  wire [7:0] t_r27_c46_8;
  wire [7:0] t_r27_c46_9;
  wire [7:0] t_r27_c46_10;
  wire [7:0] t_r27_c46_11;
  wire [7:0] t_r27_c46_12;
  wire [7:0] t_r27_c47_0;
  wire [7:0] t_r27_c47_1;
  wire [7:0] t_r27_c47_2;
  wire [7:0] t_r27_c47_3;
  wire [7:0] t_r27_c47_4;
  wire [7:0] t_r27_c47_5;
  wire [7:0] t_r27_c47_6;
  wire [7:0] t_r27_c47_7;
  wire [7:0] t_r27_c47_8;
  wire [7:0] t_r27_c47_9;
  wire [7:0] t_r27_c47_10;
  wire [7:0] t_r27_c47_11;
  wire [7:0] t_r27_c47_12;
  wire [7:0] t_r27_c48_0;
  wire [7:0] t_r27_c48_1;
  wire [7:0] t_r27_c48_2;
  wire [7:0] t_r27_c48_3;
  wire [7:0] t_r27_c48_4;
  wire [7:0] t_r27_c48_5;
  wire [7:0] t_r27_c48_6;
  wire [7:0] t_r27_c48_7;
  wire [7:0] t_r27_c48_8;
  wire [7:0] t_r27_c48_9;
  wire [7:0] t_r27_c48_10;
  wire [7:0] t_r27_c48_11;
  wire [7:0] t_r27_c48_12;
  wire [7:0] t_r27_c49_0;
  wire [7:0] t_r27_c49_1;
  wire [7:0] t_r27_c49_2;
  wire [7:0] t_r27_c49_3;
  wire [7:0] t_r27_c49_4;
  wire [7:0] t_r27_c49_5;
  wire [7:0] t_r27_c49_6;
  wire [7:0] t_r27_c49_7;
  wire [7:0] t_r27_c49_8;
  wire [7:0] t_r27_c49_9;
  wire [7:0] t_r27_c49_10;
  wire [7:0] t_r27_c49_11;
  wire [7:0] t_r27_c49_12;
  wire [7:0] t_r27_c50_0;
  wire [7:0] t_r27_c50_1;
  wire [7:0] t_r27_c50_2;
  wire [7:0] t_r27_c50_3;
  wire [7:0] t_r27_c50_4;
  wire [7:0] t_r27_c50_5;
  wire [7:0] t_r27_c50_6;
  wire [7:0] t_r27_c50_7;
  wire [7:0] t_r27_c50_8;
  wire [7:0] t_r27_c50_9;
  wire [7:0] t_r27_c50_10;
  wire [7:0] t_r27_c50_11;
  wire [7:0] t_r27_c50_12;
  wire [7:0] t_r27_c51_0;
  wire [7:0] t_r27_c51_1;
  wire [7:0] t_r27_c51_2;
  wire [7:0] t_r27_c51_3;
  wire [7:0] t_r27_c51_4;
  wire [7:0] t_r27_c51_5;
  wire [7:0] t_r27_c51_6;
  wire [7:0] t_r27_c51_7;
  wire [7:0] t_r27_c51_8;
  wire [7:0] t_r27_c51_9;
  wire [7:0] t_r27_c51_10;
  wire [7:0] t_r27_c51_11;
  wire [7:0] t_r27_c51_12;
  wire [7:0] t_r27_c52_0;
  wire [7:0] t_r27_c52_1;
  wire [7:0] t_r27_c52_2;
  wire [7:0] t_r27_c52_3;
  wire [7:0] t_r27_c52_4;
  wire [7:0] t_r27_c52_5;
  wire [7:0] t_r27_c52_6;
  wire [7:0] t_r27_c52_7;
  wire [7:0] t_r27_c52_8;
  wire [7:0] t_r27_c52_9;
  wire [7:0] t_r27_c52_10;
  wire [7:0] t_r27_c52_11;
  wire [7:0] t_r27_c52_12;
  wire [7:0] t_r27_c53_0;
  wire [7:0] t_r27_c53_1;
  wire [7:0] t_r27_c53_2;
  wire [7:0] t_r27_c53_3;
  wire [7:0] t_r27_c53_4;
  wire [7:0] t_r27_c53_5;
  wire [7:0] t_r27_c53_6;
  wire [7:0] t_r27_c53_7;
  wire [7:0] t_r27_c53_8;
  wire [7:0] t_r27_c53_9;
  wire [7:0] t_r27_c53_10;
  wire [7:0] t_r27_c53_11;
  wire [7:0] t_r27_c53_12;
  wire [7:0] t_r27_c54_0;
  wire [7:0] t_r27_c54_1;
  wire [7:0] t_r27_c54_2;
  wire [7:0] t_r27_c54_3;
  wire [7:0] t_r27_c54_4;
  wire [7:0] t_r27_c54_5;
  wire [7:0] t_r27_c54_6;
  wire [7:0] t_r27_c54_7;
  wire [7:0] t_r27_c54_8;
  wire [7:0] t_r27_c54_9;
  wire [7:0] t_r27_c54_10;
  wire [7:0] t_r27_c54_11;
  wire [7:0] t_r27_c54_12;
  wire [7:0] t_r27_c55_0;
  wire [7:0] t_r27_c55_1;
  wire [7:0] t_r27_c55_2;
  wire [7:0] t_r27_c55_3;
  wire [7:0] t_r27_c55_4;
  wire [7:0] t_r27_c55_5;
  wire [7:0] t_r27_c55_6;
  wire [7:0] t_r27_c55_7;
  wire [7:0] t_r27_c55_8;
  wire [7:0] t_r27_c55_9;
  wire [7:0] t_r27_c55_10;
  wire [7:0] t_r27_c55_11;
  wire [7:0] t_r27_c55_12;
  wire [7:0] t_r27_c56_0;
  wire [7:0] t_r27_c56_1;
  wire [7:0] t_r27_c56_2;
  wire [7:0] t_r27_c56_3;
  wire [7:0] t_r27_c56_4;
  wire [7:0] t_r27_c56_5;
  wire [7:0] t_r27_c56_6;
  wire [7:0] t_r27_c56_7;
  wire [7:0] t_r27_c56_8;
  wire [7:0] t_r27_c56_9;
  wire [7:0] t_r27_c56_10;
  wire [7:0] t_r27_c56_11;
  wire [7:0] t_r27_c56_12;
  wire [7:0] t_r27_c57_0;
  wire [7:0] t_r27_c57_1;
  wire [7:0] t_r27_c57_2;
  wire [7:0] t_r27_c57_3;
  wire [7:0] t_r27_c57_4;
  wire [7:0] t_r27_c57_5;
  wire [7:0] t_r27_c57_6;
  wire [7:0] t_r27_c57_7;
  wire [7:0] t_r27_c57_8;
  wire [7:0] t_r27_c57_9;
  wire [7:0] t_r27_c57_10;
  wire [7:0] t_r27_c57_11;
  wire [7:0] t_r27_c57_12;
  wire [7:0] t_r27_c58_0;
  wire [7:0] t_r27_c58_1;
  wire [7:0] t_r27_c58_2;
  wire [7:0] t_r27_c58_3;
  wire [7:0] t_r27_c58_4;
  wire [7:0] t_r27_c58_5;
  wire [7:0] t_r27_c58_6;
  wire [7:0] t_r27_c58_7;
  wire [7:0] t_r27_c58_8;
  wire [7:0] t_r27_c58_9;
  wire [7:0] t_r27_c58_10;
  wire [7:0] t_r27_c58_11;
  wire [7:0] t_r27_c58_12;
  wire [7:0] t_r27_c59_0;
  wire [7:0] t_r27_c59_1;
  wire [7:0] t_r27_c59_2;
  wire [7:0] t_r27_c59_3;
  wire [7:0] t_r27_c59_4;
  wire [7:0] t_r27_c59_5;
  wire [7:0] t_r27_c59_6;
  wire [7:0] t_r27_c59_7;
  wire [7:0] t_r27_c59_8;
  wire [7:0] t_r27_c59_9;
  wire [7:0] t_r27_c59_10;
  wire [7:0] t_r27_c59_11;
  wire [7:0] t_r27_c59_12;
  wire [7:0] t_r27_c60_0;
  wire [7:0] t_r27_c60_1;
  wire [7:0] t_r27_c60_2;
  wire [7:0] t_r27_c60_3;
  wire [7:0] t_r27_c60_4;
  wire [7:0] t_r27_c60_5;
  wire [7:0] t_r27_c60_6;
  wire [7:0] t_r27_c60_7;
  wire [7:0] t_r27_c60_8;
  wire [7:0] t_r27_c60_9;
  wire [7:0] t_r27_c60_10;
  wire [7:0] t_r27_c60_11;
  wire [7:0] t_r27_c60_12;
  wire [7:0] t_r27_c61_0;
  wire [7:0] t_r27_c61_1;
  wire [7:0] t_r27_c61_2;
  wire [7:0] t_r27_c61_3;
  wire [7:0] t_r27_c61_4;
  wire [7:0] t_r27_c61_5;
  wire [7:0] t_r27_c61_6;
  wire [7:0] t_r27_c61_7;
  wire [7:0] t_r27_c61_8;
  wire [7:0] t_r27_c61_9;
  wire [7:0] t_r27_c61_10;
  wire [7:0] t_r27_c61_11;
  wire [7:0] t_r27_c61_12;
  wire [7:0] t_r27_c62_0;
  wire [7:0] t_r27_c62_1;
  wire [7:0] t_r27_c62_2;
  wire [7:0] t_r27_c62_3;
  wire [7:0] t_r27_c62_4;
  wire [7:0] t_r27_c62_5;
  wire [7:0] t_r27_c62_6;
  wire [7:0] t_r27_c62_7;
  wire [7:0] t_r27_c62_8;
  wire [7:0] t_r27_c62_9;
  wire [7:0] t_r27_c62_10;
  wire [7:0] t_r27_c62_11;
  wire [7:0] t_r27_c62_12;
  wire [7:0] t_r27_c63_0;
  wire [7:0] t_r27_c63_1;
  wire [7:0] t_r27_c63_2;
  wire [7:0] t_r27_c63_3;
  wire [7:0] t_r27_c63_4;
  wire [7:0] t_r27_c63_5;
  wire [7:0] t_r27_c63_6;
  wire [7:0] t_r27_c63_7;
  wire [7:0] t_r27_c63_8;
  wire [7:0] t_r27_c63_9;
  wire [7:0] t_r27_c63_10;
  wire [7:0] t_r27_c63_11;
  wire [7:0] t_r27_c63_12;
  wire [7:0] t_r27_c64_0;
  wire [7:0] t_r27_c64_1;
  wire [7:0] t_r27_c64_2;
  wire [7:0] t_r27_c64_3;
  wire [7:0] t_r27_c64_4;
  wire [7:0] t_r27_c64_5;
  wire [7:0] t_r27_c64_6;
  wire [7:0] t_r27_c64_7;
  wire [7:0] t_r27_c64_8;
  wire [7:0] t_r27_c64_9;
  wire [7:0] t_r27_c64_10;
  wire [7:0] t_r27_c64_11;
  wire [7:0] t_r27_c64_12;
  wire [7:0] t_r27_c65_0;
  wire [7:0] t_r27_c65_1;
  wire [7:0] t_r27_c65_2;
  wire [7:0] t_r27_c65_3;
  wire [7:0] t_r27_c65_4;
  wire [7:0] t_r27_c65_5;
  wire [7:0] t_r27_c65_6;
  wire [7:0] t_r27_c65_7;
  wire [7:0] t_r27_c65_8;
  wire [7:0] t_r27_c65_9;
  wire [7:0] t_r27_c65_10;
  wire [7:0] t_r27_c65_11;
  wire [7:0] t_r27_c65_12;
  wire [7:0] t_r28_c0_0;
  wire [7:0] t_r28_c0_1;
  wire [7:0] t_r28_c0_2;
  wire [7:0] t_r28_c0_3;
  wire [7:0] t_r28_c0_4;
  wire [7:0] t_r28_c0_5;
  wire [7:0] t_r28_c0_6;
  wire [7:0] t_r28_c0_7;
  wire [7:0] t_r28_c0_8;
  wire [7:0] t_r28_c0_9;
  wire [7:0] t_r28_c0_10;
  wire [7:0] t_r28_c0_11;
  wire [7:0] t_r28_c0_12;
  wire [7:0] t_r28_c1_0;
  wire [7:0] t_r28_c1_1;
  wire [7:0] t_r28_c1_2;
  wire [7:0] t_r28_c1_3;
  wire [7:0] t_r28_c1_4;
  wire [7:0] t_r28_c1_5;
  wire [7:0] t_r28_c1_6;
  wire [7:0] t_r28_c1_7;
  wire [7:0] t_r28_c1_8;
  wire [7:0] t_r28_c1_9;
  wire [7:0] t_r28_c1_10;
  wire [7:0] t_r28_c1_11;
  wire [7:0] t_r28_c1_12;
  wire [7:0] t_r28_c2_0;
  wire [7:0] t_r28_c2_1;
  wire [7:0] t_r28_c2_2;
  wire [7:0] t_r28_c2_3;
  wire [7:0] t_r28_c2_4;
  wire [7:0] t_r28_c2_5;
  wire [7:0] t_r28_c2_6;
  wire [7:0] t_r28_c2_7;
  wire [7:0] t_r28_c2_8;
  wire [7:0] t_r28_c2_9;
  wire [7:0] t_r28_c2_10;
  wire [7:0] t_r28_c2_11;
  wire [7:0] t_r28_c2_12;
  wire [7:0] t_r28_c3_0;
  wire [7:0] t_r28_c3_1;
  wire [7:0] t_r28_c3_2;
  wire [7:0] t_r28_c3_3;
  wire [7:0] t_r28_c3_4;
  wire [7:0] t_r28_c3_5;
  wire [7:0] t_r28_c3_6;
  wire [7:0] t_r28_c3_7;
  wire [7:0] t_r28_c3_8;
  wire [7:0] t_r28_c3_9;
  wire [7:0] t_r28_c3_10;
  wire [7:0] t_r28_c3_11;
  wire [7:0] t_r28_c3_12;
  wire [7:0] t_r28_c4_0;
  wire [7:0] t_r28_c4_1;
  wire [7:0] t_r28_c4_2;
  wire [7:0] t_r28_c4_3;
  wire [7:0] t_r28_c4_4;
  wire [7:0] t_r28_c4_5;
  wire [7:0] t_r28_c4_6;
  wire [7:0] t_r28_c4_7;
  wire [7:0] t_r28_c4_8;
  wire [7:0] t_r28_c4_9;
  wire [7:0] t_r28_c4_10;
  wire [7:0] t_r28_c4_11;
  wire [7:0] t_r28_c4_12;
  wire [7:0] t_r28_c5_0;
  wire [7:0] t_r28_c5_1;
  wire [7:0] t_r28_c5_2;
  wire [7:0] t_r28_c5_3;
  wire [7:0] t_r28_c5_4;
  wire [7:0] t_r28_c5_5;
  wire [7:0] t_r28_c5_6;
  wire [7:0] t_r28_c5_7;
  wire [7:0] t_r28_c5_8;
  wire [7:0] t_r28_c5_9;
  wire [7:0] t_r28_c5_10;
  wire [7:0] t_r28_c5_11;
  wire [7:0] t_r28_c5_12;
  wire [7:0] t_r28_c6_0;
  wire [7:0] t_r28_c6_1;
  wire [7:0] t_r28_c6_2;
  wire [7:0] t_r28_c6_3;
  wire [7:0] t_r28_c6_4;
  wire [7:0] t_r28_c6_5;
  wire [7:0] t_r28_c6_6;
  wire [7:0] t_r28_c6_7;
  wire [7:0] t_r28_c6_8;
  wire [7:0] t_r28_c6_9;
  wire [7:0] t_r28_c6_10;
  wire [7:0] t_r28_c6_11;
  wire [7:0] t_r28_c6_12;
  wire [7:0] t_r28_c7_0;
  wire [7:0] t_r28_c7_1;
  wire [7:0] t_r28_c7_2;
  wire [7:0] t_r28_c7_3;
  wire [7:0] t_r28_c7_4;
  wire [7:0] t_r28_c7_5;
  wire [7:0] t_r28_c7_6;
  wire [7:0] t_r28_c7_7;
  wire [7:0] t_r28_c7_8;
  wire [7:0] t_r28_c7_9;
  wire [7:0] t_r28_c7_10;
  wire [7:0] t_r28_c7_11;
  wire [7:0] t_r28_c7_12;
  wire [7:0] t_r28_c8_0;
  wire [7:0] t_r28_c8_1;
  wire [7:0] t_r28_c8_2;
  wire [7:0] t_r28_c8_3;
  wire [7:0] t_r28_c8_4;
  wire [7:0] t_r28_c8_5;
  wire [7:0] t_r28_c8_6;
  wire [7:0] t_r28_c8_7;
  wire [7:0] t_r28_c8_8;
  wire [7:0] t_r28_c8_9;
  wire [7:0] t_r28_c8_10;
  wire [7:0] t_r28_c8_11;
  wire [7:0] t_r28_c8_12;
  wire [7:0] t_r28_c9_0;
  wire [7:0] t_r28_c9_1;
  wire [7:0] t_r28_c9_2;
  wire [7:0] t_r28_c9_3;
  wire [7:0] t_r28_c9_4;
  wire [7:0] t_r28_c9_5;
  wire [7:0] t_r28_c9_6;
  wire [7:0] t_r28_c9_7;
  wire [7:0] t_r28_c9_8;
  wire [7:0] t_r28_c9_9;
  wire [7:0] t_r28_c9_10;
  wire [7:0] t_r28_c9_11;
  wire [7:0] t_r28_c9_12;
  wire [7:0] t_r28_c10_0;
  wire [7:0] t_r28_c10_1;
  wire [7:0] t_r28_c10_2;
  wire [7:0] t_r28_c10_3;
  wire [7:0] t_r28_c10_4;
  wire [7:0] t_r28_c10_5;
  wire [7:0] t_r28_c10_6;
  wire [7:0] t_r28_c10_7;
  wire [7:0] t_r28_c10_8;
  wire [7:0] t_r28_c10_9;
  wire [7:0] t_r28_c10_10;
  wire [7:0] t_r28_c10_11;
  wire [7:0] t_r28_c10_12;
  wire [7:0] t_r28_c11_0;
  wire [7:0] t_r28_c11_1;
  wire [7:0] t_r28_c11_2;
  wire [7:0] t_r28_c11_3;
  wire [7:0] t_r28_c11_4;
  wire [7:0] t_r28_c11_5;
  wire [7:0] t_r28_c11_6;
  wire [7:0] t_r28_c11_7;
  wire [7:0] t_r28_c11_8;
  wire [7:0] t_r28_c11_9;
  wire [7:0] t_r28_c11_10;
  wire [7:0] t_r28_c11_11;
  wire [7:0] t_r28_c11_12;
  wire [7:0] t_r28_c12_0;
  wire [7:0] t_r28_c12_1;
  wire [7:0] t_r28_c12_2;
  wire [7:0] t_r28_c12_3;
  wire [7:0] t_r28_c12_4;
  wire [7:0] t_r28_c12_5;
  wire [7:0] t_r28_c12_6;
  wire [7:0] t_r28_c12_7;
  wire [7:0] t_r28_c12_8;
  wire [7:0] t_r28_c12_9;
  wire [7:0] t_r28_c12_10;
  wire [7:0] t_r28_c12_11;
  wire [7:0] t_r28_c12_12;
  wire [7:0] t_r28_c13_0;
  wire [7:0] t_r28_c13_1;
  wire [7:0] t_r28_c13_2;
  wire [7:0] t_r28_c13_3;
  wire [7:0] t_r28_c13_4;
  wire [7:0] t_r28_c13_5;
  wire [7:0] t_r28_c13_6;
  wire [7:0] t_r28_c13_7;
  wire [7:0] t_r28_c13_8;
  wire [7:0] t_r28_c13_9;
  wire [7:0] t_r28_c13_10;
  wire [7:0] t_r28_c13_11;
  wire [7:0] t_r28_c13_12;
  wire [7:0] t_r28_c14_0;
  wire [7:0] t_r28_c14_1;
  wire [7:0] t_r28_c14_2;
  wire [7:0] t_r28_c14_3;
  wire [7:0] t_r28_c14_4;
  wire [7:0] t_r28_c14_5;
  wire [7:0] t_r28_c14_6;
  wire [7:0] t_r28_c14_7;
  wire [7:0] t_r28_c14_8;
  wire [7:0] t_r28_c14_9;
  wire [7:0] t_r28_c14_10;
  wire [7:0] t_r28_c14_11;
  wire [7:0] t_r28_c14_12;
  wire [7:0] t_r28_c15_0;
  wire [7:0] t_r28_c15_1;
  wire [7:0] t_r28_c15_2;
  wire [7:0] t_r28_c15_3;
  wire [7:0] t_r28_c15_4;
  wire [7:0] t_r28_c15_5;
  wire [7:0] t_r28_c15_6;
  wire [7:0] t_r28_c15_7;
  wire [7:0] t_r28_c15_8;
  wire [7:0] t_r28_c15_9;
  wire [7:0] t_r28_c15_10;
  wire [7:0] t_r28_c15_11;
  wire [7:0] t_r28_c15_12;
  wire [7:0] t_r28_c16_0;
  wire [7:0] t_r28_c16_1;
  wire [7:0] t_r28_c16_2;
  wire [7:0] t_r28_c16_3;
  wire [7:0] t_r28_c16_4;
  wire [7:0] t_r28_c16_5;
  wire [7:0] t_r28_c16_6;
  wire [7:0] t_r28_c16_7;
  wire [7:0] t_r28_c16_8;
  wire [7:0] t_r28_c16_9;
  wire [7:0] t_r28_c16_10;
  wire [7:0] t_r28_c16_11;
  wire [7:0] t_r28_c16_12;
  wire [7:0] t_r28_c17_0;
  wire [7:0] t_r28_c17_1;
  wire [7:0] t_r28_c17_2;
  wire [7:0] t_r28_c17_3;
  wire [7:0] t_r28_c17_4;
  wire [7:0] t_r28_c17_5;
  wire [7:0] t_r28_c17_6;
  wire [7:0] t_r28_c17_7;
  wire [7:0] t_r28_c17_8;
  wire [7:0] t_r28_c17_9;
  wire [7:0] t_r28_c17_10;
  wire [7:0] t_r28_c17_11;
  wire [7:0] t_r28_c17_12;
  wire [7:0] t_r28_c18_0;
  wire [7:0] t_r28_c18_1;
  wire [7:0] t_r28_c18_2;
  wire [7:0] t_r28_c18_3;
  wire [7:0] t_r28_c18_4;
  wire [7:0] t_r28_c18_5;
  wire [7:0] t_r28_c18_6;
  wire [7:0] t_r28_c18_7;
  wire [7:0] t_r28_c18_8;
  wire [7:0] t_r28_c18_9;
  wire [7:0] t_r28_c18_10;
  wire [7:0] t_r28_c18_11;
  wire [7:0] t_r28_c18_12;
  wire [7:0] t_r28_c19_0;
  wire [7:0] t_r28_c19_1;
  wire [7:0] t_r28_c19_2;
  wire [7:0] t_r28_c19_3;
  wire [7:0] t_r28_c19_4;
  wire [7:0] t_r28_c19_5;
  wire [7:0] t_r28_c19_6;
  wire [7:0] t_r28_c19_7;
  wire [7:0] t_r28_c19_8;
  wire [7:0] t_r28_c19_9;
  wire [7:0] t_r28_c19_10;
  wire [7:0] t_r28_c19_11;
  wire [7:0] t_r28_c19_12;
  wire [7:0] t_r28_c20_0;
  wire [7:0] t_r28_c20_1;
  wire [7:0] t_r28_c20_2;
  wire [7:0] t_r28_c20_3;
  wire [7:0] t_r28_c20_4;
  wire [7:0] t_r28_c20_5;
  wire [7:0] t_r28_c20_6;
  wire [7:0] t_r28_c20_7;
  wire [7:0] t_r28_c20_8;
  wire [7:0] t_r28_c20_9;
  wire [7:0] t_r28_c20_10;
  wire [7:0] t_r28_c20_11;
  wire [7:0] t_r28_c20_12;
  wire [7:0] t_r28_c21_0;
  wire [7:0] t_r28_c21_1;
  wire [7:0] t_r28_c21_2;
  wire [7:0] t_r28_c21_3;
  wire [7:0] t_r28_c21_4;
  wire [7:0] t_r28_c21_5;
  wire [7:0] t_r28_c21_6;
  wire [7:0] t_r28_c21_7;
  wire [7:0] t_r28_c21_8;
  wire [7:0] t_r28_c21_9;
  wire [7:0] t_r28_c21_10;
  wire [7:0] t_r28_c21_11;
  wire [7:0] t_r28_c21_12;
  wire [7:0] t_r28_c22_0;
  wire [7:0] t_r28_c22_1;
  wire [7:0] t_r28_c22_2;
  wire [7:0] t_r28_c22_3;
  wire [7:0] t_r28_c22_4;
  wire [7:0] t_r28_c22_5;
  wire [7:0] t_r28_c22_6;
  wire [7:0] t_r28_c22_7;
  wire [7:0] t_r28_c22_8;
  wire [7:0] t_r28_c22_9;
  wire [7:0] t_r28_c22_10;
  wire [7:0] t_r28_c22_11;
  wire [7:0] t_r28_c22_12;
  wire [7:0] t_r28_c23_0;
  wire [7:0] t_r28_c23_1;
  wire [7:0] t_r28_c23_2;
  wire [7:0] t_r28_c23_3;
  wire [7:0] t_r28_c23_4;
  wire [7:0] t_r28_c23_5;
  wire [7:0] t_r28_c23_6;
  wire [7:0] t_r28_c23_7;
  wire [7:0] t_r28_c23_8;
  wire [7:0] t_r28_c23_9;
  wire [7:0] t_r28_c23_10;
  wire [7:0] t_r28_c23_11;
  wire [7:0] t_r28_c23_12;
  wire [7:0] t_r28_c24_0;
  wire [7:0] t_r28_c24_1;
  wire [7:0] t_r28_c24_2;
  wire [7:0] t_r28_c24_3;
  wire [7:0] t_r28_c24_4;
  wire [7:0] t_r28_c24_5;
  wire [7:0] t_r28_c24_6;
  wire [7:0] t_r28_c24_7;
  wire [7:0] t_r28_c24_8;
  wire [7:0] t_r28_c24_9;
  wire [7:0] t_r28_c24_10;
  wire [7:0] t_r28_c24_11;
  wire [7:0] t_r28_c24_12;
  wire [7:0] t_r28_c25_0;
  wire [7:0] t_r28_c25_1;
  wire [7:0] t_r28_c25_2;
  wire [7:0] t_r28_c25_3;
  wire [7:0] t_r28_c25_4;
  wire [7:0] t_r28_c25_5;
  wire [7:0] t_r28_c25_6;
  wire [7:0] t_r28_c25_7;
  wire [7:0] t_r28_c25_8;
  wire [7:0] t_r28_c25_9;
  wire [7:0] t_r28_c25_10;
  wire [7:0] t_r28_c25_11;
  wire [7:0] t_r28_c25_12;
  wire [7:0] t_r28_c26_0;
  wire [7:0] t_r28_c26_1;
  wire [7:0] t_r28_c26_2;
  wire [7:0] t_r28_c26_3;
  wire [7:0] t_r28_c26_4;
  wire [7:0] t_r28_c26_5;
  wire [7:0] t_r28_c26_6;
  wire [7:0] t_r28_c26_7;
  wire [7:0] t_r28_c26_8;
  wire [7:0] t_r28_c26_9;
  wire [7:0] t_r28_c26_10;
  wire [7:0] t_r28_c26_11;
  wire [7:0] t_r28_c26_12;
  wire [7:0] t_r28_c27_0;
  wire [7:0] t_r28_c27_1;
  wire [7:0] t_r28_c27_2;
  wire [7:0] t_r28_c27_3;
  wire [7:0] t_r28_c27_4;
  wire [7:0] t_r28_c27_5;
  wire [7:0] t_r28_c27_6;
  wire [7:0] t_r28_c27_7;
  wire [7:0] t_r28_c27_8;
  wire [7:0] t_r28_c27_9;
  wire [7:0] t_r28_c27_10;
  wire [7:0] t_r28_c27_11;
  wire [7:0] t_r28_c27_12;
  wire [7:0] t_r28_c28_0;
  wire [7:0] t_r28_c28_1;
  wire [7:0] t_r28_c28_2;
  wire [7:0] t_r28_c28_3;
  wire [7:0] t_r28_c28_4;
  wire [7:0] t_r28_c28_5;
  wire [7:0] t_r28_c28_6;
  wire [7:0] t_r28_c28_7;
  wire [7:0] t_r28_c28_8;
  wire [7:0] t_r28_c28_9;
  wire [7:0] t_r28_c28_10;
  wire [7:0] t_r28_c28_11;
  wire [7:0] t_r28_c28_12;
  wire [7:0] t_r28_c29_0;
  wire [7:0] t_r28_c29_1;
  wire [7:0] t_r28_c29_2;
  wire [7:0] t_r28_c29_3;
  wire [7:0] t_r28_c29_4;
  wire [7:0] t_r28_c29_5;
  wire [7:0] t_r28_c29_6;
  wire [7:0] t_r28_c29_7;
  wire [7:0] t_r28_c29_8;
  wire [7:0] t_r28_c29_9;
  wire [7:0] t_r28_c29_10;
  wire [7:0] t_r28_c29_11;
  wire [7:0] t_r28_c29_12;
  wire [7:0] t_r28_c30_0;
  wire [7:0] t_r28_c30_1;
  wire [7:0] t_r28_c30_2;
  wire [7:0] t_r28_c30_3;
  wire [7:0] t_r28_c30_4;
  wire [7:0] t_r28_c30_5;
  wire [7:0] t_r28_c30_6;
  wire [7:0] t_r28_c30_7;
  wire [7:0] t_r28_c30_8;
  wire [7:0] t_r28_c30_9;
  wire [7:0] t_r28_c30_10;
  wire [7:0] t_r28_c30_11;
  wire [7:0] t_r28_c30_12;
  wire [7:0] t_r28_c31_0;
  wire [7:0] t_r28_c31_1;
  wire [7:0] t_r28_c31_2;
  wire [7:0] t_r28_c31_3;
  wire [7:0] t_r28_c31_4;
  wire [7:0] t_r28_c31_5;
  wire [7:0] t_r28_c31_6;
  wire [7:0] t_r28_c31_7;
  wire [7:0] t_r28_c31_8;
  wire [7:0] t_r28_c31_9;
  wire [7:0] t_r28_c31_10;
  wire [7:0] t_r28_c31_11;
  wire [7:0] t_r28_c31_12;
  wire [7:0] t_r28_c32_0;
  wire [7:0] t_r28_c32_1;
  wire [7:0] t_r28_c32_2;
  wire [7:0] t_r28_c32_3;
  wire [7:0] t_r28_c32_4;
  wire [7:0] t_r28_c32_5;
  wire [7:0] t_r28_c32_6;
  wire [7:0] t_r28_c32_7;
  wire [7:0] t_r28_c32_8;
  wire [7:0] t_r28_c32_9;
  wire [7:0] t_r28_c32_10;
  wire [7:0] t_r28_c32_11;
  wire [7:0] t_r28_c32_12;
  wire [7:0] t_r28_c33_0;
  wire [7:0] t_r28_c33_1;
  wire [7:0] t_r28_c33_2;
  wire [7:0] t_r28_c33_3;
  wire [7:0] t_r28_c33_4;
  wire [7:0] t_r28_c33_5;
  wire [7:0] t_r28_c33_6;
  wire [7:0] t_r28_c33_7;
  wire [7:0] t_r28_c33_8;
  wire [7:0] t_r28_c33_9;
  wire [7:0] t_r28_c33_10;
  wire [7:0] t_r28_c33_11;
  wire [7:0] t_r28_c33_12;
  wire [7:0] t_r28_c34_0;
  wire [7:0] t_r28_c34_1;
  wire [7:0] t_r28_c34_2;
  wire [7:0] t_r28_c34_3;
  wire [7:0] t_r28_c34_4;
  wire [7:0] t_r28_c34_5;
  wire [7:0] t_r28_c34_6;
  wire [7:0] t_r28_c34_7;
  wire [7:0] t_r28_c34_8;
  wire [7:0] t_r28_c34_9;
  wire [7:0] t_r28_c34_10;
  wire [7:0] t_r28_c34_11;
  wire [7:0] t_r28_c34_12;
  wire [7:0] t_r28_c35_0;
  wire [7:0] t_r28_c35_1;
  wire [7:0] t_r28_c35_2;
  wire [7:0] t_r28_c35_3;
  wire [7:0] t_r28_c35_4;
  wire [7:0] t_r28_c35_5;
  wire [7:0] t_r28_c35_6;
  wire [7:0] t_r28_c35_7;
  wire [7:0] t_r28_c35_8;
  wire [7:0] t_r28_c35_9;
  wire [7:0] t_r28_c35_10;
  wire [7:0] t_r28_c35_11;
  wire [7:0] t_r28_c35_12;
  wire [7:0] t_r28_c36_0;
  wire [7:0] t_r28_c36_1;
  wire [7:0] t_r28_c36_2;
  wire [7:0] t_r28_c36_3;
  wire [7:0] t_r28_c36_4;
  wire [7:0] t_r28_c36_5;
  wire [7:0] t_r28_c36_6;
  wire [7:0] t_r28_c36_7;
  wire [7:0] t_r28_c36_8;
  wire [7:0] t_r28_c36_9;
  wire [7:0] t_r28_c36_10;
  wire [7:0] t_r28_c36_11;
  wire [7:0] t_r28_c36_12;
  wire [7:0] t_r28_c37_0;
  wire [7:0] t_r28_c37_1;
  wire [7:0] t_r28_c37_2;
  wire [7:0] t_r28_c37_3;
  wire [7:0] t_r28_c37_4;
  wire [7:0] t_r28_c37_5;
  wire [7:0] t_r28_c37_6;
  wire [7:0] t_r28_c37_7;
  wire [7:0] t_r28_c37_8;
  wire [7:0] t_r28_c37_9;
  wire [7:0] t_r28_c37_10;
  wire [7:0] t_r28_c37_11;
  wire [7:0] t_r28_c37_12;
  wire [7:0] t_r28_c38_0;
  wire [7:0] t_r28_c38_1;
  wire [7:0] t_r28_c38_2;
  wire [7:0] t_r28_c38_3;
  wire [7:0] t_r28_c38_4;
  wire [7:0] t_r28_c38_5;
  wire [7:0] t_r28_c38_6;
  wire [7:0] t_r28_c38_7;
  wire [7:0] t_r28_c38_8;
  wire [7:0] t_r28_c38_9;
  wire [7:0] t_r28_c38_10;
  wire [7:0] t_r28_c38_11;
  wire [7:0] t_r28_c38_12;
  wire [7:0] t_r28_c39_0;
  wire [7:0] t_r28_c39_1;
  wire [7:0] t_r28_c39_2;
  wire [7:0] t_r28_c39_3;
  wire [7:0] t_r28_c39_4;
  wire [7:0] t_r28_c39_5;
  wire [7:0] t_r28_c39_6;
  wire [7:0] t_r28_c39_7;
  wire [7:0] t_r28_c39_8;
  wire [7:0] t_r28_c39_9;
  wire [7:0] t_r28_c39_10;
  wire [7:0] t_r28_c39_11;
  wire [7:0] t_r28_c39_12;
  wire [7:0] t_r28_c40_0;
  wire [7:0] t_r28_c40_1;
  wire [7:0] t_r28_c40_2;
  wire [7:0] t_r28_c40_3;
  wire [7:0] t_r28_c40_4;
  wire [7:0] t_r28_c40_5;
  wire [7:0] t_r28_c40_6;
  wire [7:0] t_r28_c40_7;
  wire [7:0] t_r28_c40_8;
  wire [7:0] t_r28_c40_9;
  wire [7:0] t_r28_c40_10;
  wire [7:0] t_r28_c40_11;
  wire [7:0] t_r28_c40_12;
  wire [7:0] t_r28_c41_0;
  wire [7:0] t_r28_c41_1;
  wire [7:0] t_r28_c41_2;
  wire [7:0] t_r28_c41_3;
  wire [7:0] t_r28_c41_4;
  wire [7:0] t_r28_c41_5;
  wire [7:0] t_r28_c41_6;
  wire [7:0] t_r28_c41_7;
  wire [7:0] t_r28_c41_8;
  wire [7:0] t_r28_c41_9;
  wire [7:0] t_r28_c41_10;
  wire [7:0] t_r28_c41_11;
  wire [7:0] t_r28_c41_12;
  wire [7:0] t_r28_c42_0;
  wire [7:0] t_r28_c42_1;
  wire [7:0] t_r28_c42_2;
  wire [7:0] t_r28_c42_3;
  wire [7:0] t_r28_c42_4;
  wire [7:0] t_r28_c42_5;
  wire [7:0] t_r28_c42_6;
  wire [7:0] t_r28_c42_7;
  wire [7:0] t_r28_c42_8;
  wire [7:0] t_r28_c42_9;
  wire [7:0] t_r28_c42_10;
  wire [7:0] t_r28_c42_11;
  wire [7:0] t_r28_c42_12;
  wire [7:0] t_r28_c43_0;
  wire [7:0] t_r28_c43_1;
  wire [7:0] t_r28_c43_2;
  wire [7:0] t_r28_c43_3;
  wire [7:0] t_r28_c43_4;
  wire [7:0] t_r28_c43_5;
  wire [7:0] t_r28_c43_6;
  wire [7:0] t_r28_c43_7;
  wire [7:0] t_r28_c43_8;
  wire [7:0] t_r28_c43_9;
  wire [7:0] t_r28_c43_10;
  wire [7:0] t_r28_c43_11;
  wire [7:0] t_r28_c43_12;
  wire [7:0] t_r28_c44_0;
  wire [7:0] t_r28_c44_1;
  wire [7:0] t_r28_c44_2;
  wire [7:0] t_r28_c44_3;
  wire [7:0] t_r28_c44_4;
  wire [7:0] t_r28_c44_5;
  wire [7:0] t_r28_c44_6;
  wire [7:0] t_r28_c44_7;
  wire [7:0] t_r28_c44_8;
  wire [7:0] t_r28_c44_9;
  wire [7:0] t_r28_c44_10;
  wire [7:0] t_r28_c44_11;
  wire [7:0] t_r28_c44_12;
  wire [7:0] t_r28_c45_0;
  wire [7:0] t_r28_c45_1;
  wire [7:0] t_r28_c45_2;
  wire [7:0] t_r28_c45_3;
  wire [7:0] t_r28_c45_4;
  wire [7:0] t_r28_c45_5;
  wire [7:0] t_r28_c45_6;
  wire [7:0] t_r28_c45_7;
  wire [7:0] t_r28_c45_8;
  wire [7:0] t_r28_c45_9;
  wire [7:0] t_r28_c45_10;
  wire [7:0] t_r28_c45_11;
  wire [7:0] t_r28_c45_12;
  wire [7:0] t_r28_c46_0;
  wire [7:0] t_r28_c46_1;
  wire [7:0] t_r28_c46_2;
  wire [7:0] t_r28_c46_3;
  wire [7:0] t_r28_c46_4;
  wire [7:0] t_r28_c46_5;
  wire [7:0] t_r28_c46_6;
  wire [7:0] t_r28_c46_7;
  wire [7:0] t_r28_c46_8;
  wire [7:0] t_r28_c46_9;
  wire [7:0] t_r28_c46_10;
  wire [7:0] t_r28_c46_11;
  wire [7:0] t_r28_c46_12;
  wire [7:0] t_r28_c47_0;
  wire [7:0] t_r28_c47_1;
  wire [7:0] t_r28_c47_2;
  wire [7:0] t_r28_c47_3;
  wire [7:0] t_r28_c47_4;
  wire [7:0] t_r28_c47_5;
  wire [7:0] t_r28_c47_6;
  wire [7:0] t_r28_c47_7;
  wire [7:0] t_r28_c47_8;
  wire [7:0] t_r28_c47_9;
  wire [7:0] t_r28_c47_10;
  wire [7:0] t_r28_c47_11;
  wire [7:0] t_r28_c47_12;
  wire [7:0] t_r28_c48_0;
  wire [7:0] t_r28_c48_1;
  wire [7:0] t_r28_c48_2;
  wire [7:0] t_r28_c48_3;
  wire [7:0] t_r28_c48_4;
  wire [7:0] t_r28_c48_5;
  wire [7:0] t_r28_c48_6;
  wire [7:0] t_r28_c48_7;
  wire [7:0] t_r28_c48_8;
  wire [7:0] t_r28_c48_9;
  wire [7:0] t_r28_c48_10;
  wire [7:0] t_r28_c48_11;
  wire [7:0] t_r28_c48_12;
  wire [7:0] t_r28_c49_0;
  wire [7:0] t_r28_c49_1;
  wire [7:0] t_r28_c49_2;
  wire [7:0] t_r28_c49_3;
  wire [7:0] t_r28_c49_4;
  wire [7:0] t_r28_c49_5;
  wire [7:0] t_r28_c49_6;
  wire [7:0] t_r28_c49_7;
  wire [7:0] t_r28_c49_8;
  wire [7:0] t_r28_c49_9;
  wire [7:0] t_r28_c49_10;
  wire [7:0] t_r28_c49_11;
  wire [7:0] t_r28_c49_12;
  wire [7:0] t_r28_c50_0;
  wire [7:0] t_r28_c50_1;
  wire [7:0] t_r28_c50_2;
  wire [7:0] t_r28_c50_3;
  wire [7:0] t_r28_c50_4;
  wire [7:0] t_r28_c50_5;
  wire [7:0] t_r28_c50_6;
  wire [7:0] t_r28_c50_7;
  wire [7:0] t_r28_c50_8;
  wire [7:0] t_r28_c50_9;
  wire [7:0] t_r28_c50_10;
  wire [7:0] t_r28_c50_11;
  wire [7:0] t_r28_c50_12;
  wire [7:0] t_r28_c51_0;
  wire [7:0] t_r28_c51_1;
  wire [7:0] t_r28_c51_2;
  wire [7:0] t_r28_c51_3;
  wire [7:0] t_r28_c51_4;
  wire [7:0] t_r28_c51_5;
  wire [7:0] t_r28_c51_6;
  wire [7:0] t_r28_c51_7;
  wire [7:0] t_r28_c51_8;
  wire [7:0] t_r28_c51_9;
  wire [7:0] t_r28_c51_10;
  wire [7:0] t_r28_c51_11;
  wire [7:0] t_r28_c51_12;
  wire [7:0] t_r28_c52_0;
  wire [7:0] t_r28_c52_1;
  wire [7:0] t_r28_c52_2;
  wire [7:0] t_r28_c52_3;
  wire [7:0] t_r28_c52_4;
  wire [7:0] t_r28_c52_5;
  wire [7:0] t_r28_c52_6;
  wire [7:0] t_r28_c52_7;
  wire [7:0] t_r28_c52_8;
  wire [7:0] t_r28_c52_9;
  wire [7:0] t_r28_c52_10;
  wire [7:0] t_r28_c52_11;
  wire [7:0] t_r28_c52_12;
  wire [7:0] t_r28_c53_0;
  wire [7:0] t_r28_c53_1;
  wire [7:0] t_r28_c53_2;
  wire [7:0] t_r28_c53_3;
  wire [7:0] t_r28_c53_4;
  wire [7:0] t_r28_c53_5;
  wire [7:0] t_r28_c53_6;
  wire [7:0] t_r28_c53_7;
  wire [7:0] t_r28_c53_8;
  wire [7:0] t_r28_c53_9;
  wire [7:0] t_r28_c53_10;
  wire [7:0] t_r28_c53_11;
  wire [7:0] t_r28_c53_12;
  wire [7:0] t_r28_c54_0;
  wire [7:0] t_r28_c54_1;
  wire [7:0] t_r28_c54_2;
  wire [7:0] t_r28_c54_3;
  wire [7:0] t_r28_c54_4;
  wire [7:0] t_r28_c54_5;
  wire [7:0] t_r28_c54_6;
  wire [7:0] t_r28_c54_7;
  wire [7:0] t_r28_c54_8;
  wire [7:0] t_r28_c54_9;
  wire [7:0] t_r28_c54_10;
  wire [7:0] t_r28_c54_11;
  wire [7:0] t_r28_c54_12;
  wire [7:0] t_r28_c55_0;
  wire [7:0] t_r28_c55_1;
  wire [7:0] t_r28_c55_2;
  wire [7:0] t_r28_c55_3;
  wire [7:0] t_r28_c55_4;
  wire [7:0] t_r28_c55_5;
  wire [7:0] t_r28_c55_6;
  wire [7:0] t_r28_c55_7;
  wire [7:0] t_r28_c55_8;
  wire [7:0] t_r28_c55_9;
  wire [7:0] t_r28_c55_10;
  wire [7:0] t_r28_c55_11;
  wire [7:0] t_r28_c55_12;
  wire [7:0] t_r28_c56_0;
  wire [7:0] t_r28_c56_1;
  wire [7:0] t_r28_c56_2;
  wire [7:0] t_r28_c56_3;
  wire [7:0] t_r28_c56_4;
  wire [7:0] t_r28_c56_5;
  wire [7:0] t_r28_c56_6;
  wire [7:0] t_r28_c56_7;
  wire [7:0] t_r28_c56_8;
  wire [7:0] t_r28_c56_9;
  wire [7:0] t_r28_c56_10;
  wire [7:0] t_r28_c56_11;
  wire [7:0] t_r28_c56_12;
  wire [7:0] t_r28_c57_0;
  wire [7:0] t_r28_c57_1;
  wire [7:0] t_r28_c57_2;
  wire [7:0] t_r28_c57_3;
  wire [7:0] t_r28_c57_4;
  wire [7:0] t_r28_c57_5;
  wire [7:0] t_r28_c57_6;
  wire [7:0] t_r28_c57_7;
  wire [7:0] t_r28_c57_8;
  wire [7:0] t_r28_c57_9;
  wire [7:0] t_r28_c57_10;
  wire [7:0] t_r28_c57_11;
  wire [7:0] t_r28_c57_12;
  wire [7:0] t_r28_c58_0;
  wire [7:0] t_r28_c58_1;
  wire [7:0] t_r28_c58_2;
  wire [7:0] t_r28_c58_3;
  wire [7:0] t_r28_c58_4;
  wire [7:0] t_r28_c58_5;
  wire [7:0] t_r28_c58_6;
  wire [7:0] t_r28_c58_7;
  wire [7:0] t_r28_c58_8;
  wire [7:0] t_r28_c58_9;
  wire [7:0] t_r28_c58_10;
  wire [7:0] t_r28_c58_11;
  wire [7:0] t_r28_c58_12;
  wire [7:0] t_r28_c59_0;
  wire [7:0] t_r28_c59_1;
  wire [7:0] t_r28_c59_2;
  wire [7:0] t_r28_c59_3;
  wire [7:0] t_r28_c59_4;
  wire [7:0] t_r28_c59_5;
  wire [7:0] t_r28_c59_6;
  wire [7:0] t_r28_c59_7;
  wire [7:0] t_r28_c59_8;
  wire [7:0] t_r28_c59_9;
  wire [7:0] t_r28_c59_10;
  wire [7:0] t_r28_c59_11;
  wire [7:0] t_r28_c59_12;
  wire [7:0] t_r28_c60_0;
  wire [7:0] t_r28_c60_1;
  wire [7:0] t_r28_c60_2;
  wire [7:0] t_r28_c60_3;
  wire [7:0] t_r28_c60_4;
  wire [7:0] t_r28_c60_5;
  wire [7:0] t_r28_c60_6;
  wire [7:0] t_r28_c60_7;
  wire [7:0] t_r28_c60_8;
  wire [7:0] t_r28_c60_9;
  wire [7:0] t_r28_c60_10;
  wire [7:0] t_r28_c60_11;
  wire [7:0] t_r28_c60_12;
  wire [7:0] t_r28_c61_0;
  wire [7:0] t_r28_c61_1;
  wire [7:0] t_r28_c61_2;
  wire [7:0] t_r28_c61_3;
  wire [7:0] t_r28_c61_4;
  wire [7:0] t_r28_c61_5;
  wire [7:0] t_r28_c61_6;
  wire [7:0] t_r28_c61_7;
  wire [7:0] t_r28_c61_8;
  wire [7:0] t_r28_c61_9;
  wire [7:0] t_r28_c61_10;
  wire [7:0] t_r28_c61_11;
  wire [7:0] t_r28_c61_12;
  wire [7:0] t_r28_c62_0;
  wire [7:0] t_r28_c62_1;
  wire [7:0] t_r28_c62_2;
  wire [7:0] t_r28_c62_3;
  wire [7:0] t_r28_c62_4;
  wire [7:0] t_r28_c62_5;
  wire [7:0] t_r28_c62_6;
  wire [7:0] t_r28_c62_7;
  wire [7:0] t_r28_c62_8;
  wire [7:0] t_r28_c62_9;
  wire [7:0] t_r28_c62_10;
  wire [7:0] t_r28_c62_11;
  wire [7:0] t_r28_c62_12;
  wire [7:0] t_r28_c63_0;
  wire [7:0] t_r28_c63_1;
  wire [7:0] t_r28_c63_2;
  wire [7:0] t_r28_c63_3;
  wire [7:0] t_r28_c63_4;
  wire [7:0] t_r28_c63_5;
  wire [7:0] t_r28_c63_6;
  wire [7:0] t_r28_c63_7;
  wire [7:0] t_r28_c63_8;
  wire [7:0] t_r28_c63_9;
  wire [7:0] t_r28_c63_10;
  wire [7:0] t_r28_c63_11;
  wire [7:0] t_r28_c63_12;
  wire [7:0] t_r28_c64_0;
  wire [7:0] t_r28_c64_1;
  wire [7:0] t_r28_c64_2;
  wire [7:0] t_r28_c64_3;
  wire [7:0] t_r28_c64_4;
  wire [7:0] t_r28_c64_5;
  wire [7:0] t_r28_c64_6;
  wire [7:0] t_r28_c64_7;
  wire [7:0] t_r28_c64_8;
  wire [7:0] t_r28_c64_9;
  wire [7:0] t_r28_c64_10;
  wire [7:0] t_r28_c64_11;
  wire [7:0] t_r28_c64_12;
  wire [7:0] t_r28_c65_0;
  wire [7:0] t_r28_c65_1;
  wire [7:0] t_r28_c65_2;
  wire [7:0] t_r28_c65_3;
  wire [7:0] t_r28_c65_4;
  wire [7:0] t_r28_c65_5;
  wire [7:0] t_r28_c65_6;
  wire [7:0] t_r28_c65_7;
  wire [7:0] t_r28_c65_8;
  wire [7:0] t_r28_c65_9;
  wire [7:0] t_r28_c65_10;
  wire [7:0] t_r28_c65_11;
  wire [7:0] t_r28_c65_12;
  wire [7:0] t_r29_c0_0;
  wire [7:0] t_r29_c0_1;
  wire [7:0] t_r29_c0_2;
  wire [7:0] t_r29_c0_3;
  wire [7:0] t_r29_c0_4;
  wire [7:0] t_r29_c0_5;
  wire [7:0] t_r29_c0_6;
  wire [7:0] t_r29_c0_7;
  wire [7:0] t_r29_c0_8;
  wire [7:0] t_r29_c0_9;
  wire [7:0] t_r29_c0_10;
  wire [7:0] t_r29_c0_11;
  wire [7:0] t_r29_c0_12;
  wire [7:0] t_r29_c1_0;
  wire [7:0] t_r29_c1_1;
  wire [7:0] t_r29_c1_2;
  wire [7:0] t_r29_c1_3;
  wire [7:0] t_r29_c1_4;
  wire [7:0] t_r29_c1_5;
  wire [7:0] t_r29_c1_6;
  wire [7:0] t_r29_c1_7;
  wire [7:0] t_r29_c1_8;
  wire [7:0] t_r29_c1_9;
  wire [7:0] t_r29_c1_10;
  wire [7:0] t_r29_c1_11;
  wire [7:0] t_r29_c1_12;
  wire [7:0] t_r29_c2_0;
  wire [7:0] t_r29_c2_1;
  wire [7:0] t_r29_c2_2;
  wire [7:0] t_r29_c2_3;
  wire [7:0] t_r29_c2_4;
  wire [7:0] t_r29_c2_5;
  wire [7:0] t_r29_c2_6;
  wire [7:0] t_r29_c2_7;
  wire [7:0] t_r29_c2_8;
  wire [7:0] t_r29_c2_9;
  wire [7:0] t_r29_c2_10;
  wire [7:0] t_r29_c2_11;
  wire [7:0] t_r29_c2_12;
  wire [7:0] t_r29_c3_0;
  wire [7:0] t_r29_c3_1;
  wire [7:0] t_r29_c3_2;
  wire [7:0] t_r29_c3_3;
  wire [7:0] t_r29_c3_4;
  wire [7:0] t_r29_c3_5;
  wire [7:0] t_r29_c3_6;
  wire [7:0] t_r29_c3_7;
  wire [7:0] t_r29_c3_8;
  wire [7:0] t_r29_c3_9;
  wire [7:0] t_r29_c3_10;
  wire [7:0] t_r29_c3_11;
  wire [7:0] t_r29_c3_12;
  wire [7:0] t_r29_c4_0;
  wire [7:0] t_r29_c4_1;
  wire [7:0] t_r29_c4_2;
  wire [7:0] t_r29_c4_3;
  wire [7:0] t_r29_c4_4;
  wire [7:0] t_r29_c4_5;
  wire [7:0] t_r29_c4_6;
  wire [7:0] t_r29_c4_7;
  wire [7:0] t_r29_c4_8;
  wire [7:0] t_r29_c4_9;
  wire [7:0] t_r29_c4_10;
  wire [7:0] t_r29_c4_11;
  wire [7:0] t_r29_c4_12;
  wire [7:0] t_r29_c5_0;
  wire [7:0] t_r29_c5_1;
  wire [7:0] t_r29_c5_2;
  wire [7:0] t_r29_c5_3;
  wire [7:0] t_r29_c5_4;
  wire [7:0] t_r29_c5_5;
  wire [7:0] t_r29_c5_6;
  wire [7:0] t_r29_c5_7;
  wire [7:0] t_r29_c5_8;
  wire [7:0] t_r29_c5_9;
  wire [7:0] t_r29_c5_10;
  wire [7:0] t_r29_c5_11;
  wire [7:0] t_r29_c5_12;
  wire [7:0] t_r29_c6_0;
  wire [7:0] t_r29_c6_1;
  wire [7:0] t_r29_c6_2;
  wire [7:0] t_r29_c6_3;
  wire [7:0] t_r29_c6_4;
  wire [7:0] t_r29_c6_5;
  wire [7:0] t_r29_c6_6;
  wire [7:0] t_r29_c6_7;
  wire [7:0] t_r29_c6_8;
  wire [7:0] t_r29_c6_9;
  wire [7:0] t_r29_c6_10;
  wire [7:0] t_r29_c6_11;
  wire [7:0] t_r29_c6_12;
  wire [7:0] t_r29_c7_0;
  wire [7:0] t_r29_c7_1;
  wire [7:0] t_r29_c7_2;
  wire [7:0] t_r29_c7_3;
  wire [7:0] t_r29_c7_4;
  wire [7:0] t_r29_c7_5;
  wire [7:0] t_r29_c7_6;
  wire [7:0] t_r29_c7_7;
  wire [7:0] t_r29_c7_8;
  wire [7:0] t_r29_c7_9;
  wire [7:0] t_r29_c7_10;
  wire [7:0] t_r29_c7_11;
  wire [7:0] t_r29_c7_12;
  wire [7:0] t_r29_c8_0;
  wire [7:0] t_r29_c8_1;
  wire [7:0] t_r29_c8_2;
  wire [7:0] t_r29_c8_3;
  wire [7:0] t_r29_c8_4;
  wire [7:0] t_r29_c8_5;
  wire [7:0] t_r29_c8_6;
  wire [7:0] t_r29_c8_7;
  wire [7:0] t_r29_c8_8;
  wire [7:0] t_r29_c8_9;
  wire [7:0] t_r29_c8_10;
  wire [7:0] t_r29_c8_11;
  wire [7:0] t_r29_c8_12;
  wire [7:0] t_r29_c9_0;
  wire [7:0] t_r29_c9_1;
  wire [7:0] t_r29_c9_2;
  wire [7:0] t_r29_c9_3;
  wire [7:0] t_r29_c9_4;
  wire [7:0] t_r29_c9_5;
  wire [7:0] t_r29_c9_6;
  wire [7:0] t_r29_c9_7;
  wire [7:0] t_r29_c9_8;
  wire [7:0] t_r29_c9_9;
  wire [7:0] t_r29_c9_10;
  wire [7:0] t_r29_c9_11;
  wire [7:0] t_r29_c9_12;
  wire [7:0] t_r29_c10_0;
  wire [7:0] t_r29_c10_1;
  wire [7:0] t_r29_c10_2;
  wire [7:0] t_r29_c10_3;
  wire [7:0] t_r29_c10_4;
  wire [7:0] t_r29_c10_5;
  wire [7:0] t_r29_c10_6;
  wire [7:0] t_r29_c10_7;
  wire [7:0] t_r29_c10_8;
  wire [7:0] t_r29_c10_9;
  wire [7:0] t_r29_c10_10;
  wire [7:0] t_r29_c10_11;
  wire [7:0] t_r29_c10_12;
  wire [7:0] t_r29_c11_0;
  wire [7:0] t_r29_c11_1;
  wire [7:0] t_r29_c11_2;
  wire [7:0] t_r29_c11_3;
  wire [7:0] t_r29_c11_4;
  wire [7:0] t_r29_c11_5;
  wire [7:0] t_r29_c11_6;
  wire [7:0] t_r29_c11_7;
  wire [7:0] t_r29_c11_8;
  wire [7:0] t_r29_c11_9;
  wire [7:0] t_r29_c11_10;
  wire [7:0] t_r29_c11_11;
  wire [7:0] t_r29_c11_12;
  wire [7:0] t_r29_c12_0;
  wire [7:0] t_r29_c12_1;
  wire [7:0] t_r29_c12_2;
  wire [7:0] t_r29_c12_3;
  wire [7:0] t_r29_c12_4;
  wire [7:0] t_r29_c12_5;
  wire [7:0] t_r29_c12_6;
  wire [7:0] t_r29_c12_7;
  wire [7:0] t_r29_c12_8;
  wire [7:0] t_r29_c12_9;
  wire [7:0] t_r29_c12_10;
  wire [7:0] t_r29_c12_11;
  wire [7:0] t_r29_c12_12;
  wire [7:0] t_r29_c13_0;
  wire [7:0] t_r29_c13_1;
  wire [7:0] t_r29_c13_2;
  wire [7:0] t_r29_c13_3;
  wire [7:0] t_r29_c13_4;
  wire [7:0] t_r29_c13_5;
  wire [7:0] t_r29_c13_6;
  wire [7:0] t_r29_c13_7;
  wire [7:0] t_r29_c13_8;
  wire [7:0] t_r29_c13_9;
  wire [7:0] t_r29_c13_10;
  wire [7:0] t_r29_c13_11;
  wire [7:0] t_r29_c13_12;
  wire [7:0] t_r29_c14_0;
  wire [7:0] t_r29_c14_1;
  wire [7:0] t_r29_c14_2;
  wire [7:0] t_r29_c14_3;
  wire [7:0] t_r29_c14_4;
  wire [7:0] t_r29_c14_5;
  wire [7:0] t_r29_c14_6;
  wire [7:0] t_r29_c14_7;
  wire [7:0] t_r29_c14_8;
  wire [7:0] t_r29_c14_9;
  wire [7:0] t_r29_c14_10;
  wire [7:0] t_r29_c14_11;
  wire [7:0] t_r29_c14_12;
  wire [7:0] t_r29_c15_0;
  wire [7:0] t_r29_c15_1;
  wire [7:0] t_r29_c15_2;
  wire [7:0] t_r29_c15_3;
  wire [7:0] t_r29_c15_4;
  wire [7:0] t_r29_c15_5;
  wire [7:0] t_r29_c15_6;
  wire [7:0] t_r29_c15_7;
  wire [7:0] t_r29_c15_8;
  wire [7:0] t_r29_c15_9;
  wire [7:0] t_r29_c15_10;
  wire [7:0] t_r29_c15_11;
  wire [7:0] t_r29_c15_12;
  wire [7:0] t_r29_c16_0;
  wire [7:0] t_r29_c16_1;
  wire [7:0] t_r29_c16_2;
  wire [7:0] t_r29_c16_3;
  wire [7:0] t_r29_c16_4;
  wire [7:0] t_r29_c16_5;
  wire [7:0] t_r29_c16_6;
  wire [7:0] t_r29_c16_7;
  wire [7:0] t_r29_c16_8;
  wire [7:0] t_r29_c16_9;
  wire [7:0] t_r29_c16_10;
  wire [7:0] t_r29_c16_11;
  wire [7:0] t_r29_c16_12;
  wire [7:0] t_r29_c17_0;
  wire [7:0] t_r29_c17_1;
  wire [7:0] t_r29_c17_2;
  wire [7:0] t_r29_c17_3;
  wire [7:0] t_r29_c17_4;
  wire [7:0] t_r29_c17_5;
  wire [7:0] t_r29_c17_6;
  wire [7:0] t_r29_c17_7;
  wire [7:0] t_r29_c17_8;
  wire [7:0] t_r29_c17_9;
  wire [7:0] t_r29_c17_10;
  wire [7:0] t_r29_c17_11;
  wire [7:0] t_r29_c17_12;
  wire [7:0] t_r29_c18_0;
  wire [7:0] t_r29_c18_1;
  wire [7:0] t_r29_c18_2;
  wire [7:0] t_r29_c18_3;
  wire [7:0] t_r29_c18_4;
  wire [7:0] t_r29_c18_5;
  wire [7:0] t_r29_c18_6;
  wire [7:0] t_r29_c18_7;
  wire [7:0] t_r29_c18_8;
  wire [7:0] t_r29_c18_9;
  wire [7:0] t_r29_c18_10;
  wire [7:0] t_r29_c18_11;
  wire [7:0] t_r29_c18_12;
  wire [7:0] t_r29_c19_0;
  wire [7:0] t_r29_c19_1;
  wire [7:0] t_r29_c19_2;
  wire [7:0] t_r29_c19_3;
  wire [7:0] t_r29_c19_4;
  wire [7:0] t_r29_c19_5;
  wire [7:0] t_r29_c19_6;
  wire [7:0] t_r29_c19_7;
  wire [7:0] t_r29_c19_8;
  wire [7:0] t_r29_c19_9;
  wire [7:0] t_r29_c19_10;
  wire [7:0] t_r29_c19_11;
  wire [7:0] t_r29_c19_12;
  wire [7:0] t_r29_c20_0;
  wire [7:0] t_r29_c20_1;
  wire [7:0] t_r29_c20_2;
  wire [7:0] t_r29_c20_3;
  wire [7:0] t_r29_c20_4;
  wire [7:0] t_r29_c20_5;
  wire [7:0] t_r29_c20_6;
  wire [7:0] t_r29_c20_7;
  wire [7:0] t_r29_c20_8;
  wire [7:0] t_r29_c20_9;
  wire [7:0] t_r29_c20_10;
  wire [7:0] t_r29_c20_11;
  wire [7:0] t_r29_c20_12;
  wire [7:0] t_r29_c21_0;
  wire [7:0] t_r29_c21_1;
  wire [7:0] t_r29_c21_2;
  wire [7:0] t_r29_c21_3;
  wire [7:0] t_r29_c21_4;
  wire [7:0] t_r29_c21_5;
  wire [7:0] t_r29_c21_6;
  wire [7:0] t_r29_c21_7;
  wire [7:0] t_r29_c21_8;
  wire [7:0] t_r29_c21_9;
  wire [7:0] t_r29_c21_10;
  wire [7:0] t_r29_c21_11;
  wire [7:0] t_r29_c21_12;
  wire [7:0] t_r29_c22_0;
  wire [7:0] t_r29_c22_1;
  wire [7:0] t_r29_c22_2;
  wire [7:0] t_r29_c22_3;
  wire [7:0] t_r29_c22_4;
  wire [7:0] t_r29_c22_5;
  wire [7:0] t_r29_c22_6;
  wire [7:0] t_r29_c22_7;
  wire [7:0] t_r29_c22_8;
  wire [7:0] t_r29_c22_9;
  wire [7:0] t_r29_c22_10;
  wire [7:0] t_r29_c22_11;
  wire [7:0] t_r29_c22_12;
  wire [7:0] t_r29_c23_0;
  wire [7:0] t_r29_c23_1;
  wire [7:0] t_r29_c23_2;
  wire [7:0] t_r29_c23_3;
  wire [7:0] t_r29_c23_4;
  wire [7:0] t_r29_c23_5;
  wire [7:0] t_r29_c23_6;
  wire [7:0] t_r29_c23_7;
  wire [7:0] t_r29_c23_8;
  wire [7:0] t_r29_c23_9;
  wire [7:0] t_r29_c23_10;
  wire [7:0] t_r29_c23_11;
  wire [7:0] t_r29_c23_12;
  wire [7:0] t_r29_c24_0;
  wire [7:0] t_r29_c24_1;
  wire [7:0] t_r29_c24_2;
  wire [7:0] t_r29_c24_3;
  wire [7:0] t_r29_c24_4;
  wire [7:0] t_r29_c24_5;
  wire [7:0] t_r29_c24_6;
  wire [7:0] t_r29_c24_7;
  wire [7:0] t_r29_c24_8;
  wire [7:0] t_r29_c24_9;
  wire [7:0] t_r29_c24_10;
  wire [7:0] t_r29_c24_11;
  wire [7:0] t_r29_c24_12;
  wire [7:0] t_r29_c25_0;
  wire [7:0] t_r29_c25_1;
  wire [7:0] t_r29_c25_2;
  wire [7:0] t_r29_c25_3;
  wire [7:0] t_r29_c25_4;
  wire [7:0] t_r29_c25_5;
  wire [7:0] t_r29_c25_6;
  wire [7:0] t_r29_c25_7;
  wire [7:0] t_r29_c25_8;
  wire [7:0] t_r29_c25_9;
  wire [7:0] t_r29_c25_10;
  wire [7:0] t_r29_c25_11;
  wire [7:0] t_r29_c25_12;
  wire [7:0] t_r29_c26_0;
  wire [7:0] t_r29_c26_1;
  wire [7:0] t_r29_c26_2;
  wire [7:0] t_r29_c26_3;
  wire [7:0] t_r29_c26_4;
  wire [7:0] t_r29_c26_5;
  wire [7:0] t_r29_c26_6;
  wire [7:0] t_r29_c26_7;
  wire [7:0] t_r29_c26_8;
  wire [7:0] t_r29_c26_9;
  wire [7:0] t_r29_c26_10;
  wire [7:0] t_r29_c26_11;
  wire [7:0] t_r29_c26_12;
  wire [7:0] t_r29_c27_0;
  wire [7:0] t_r29_c27_1;
  wire [7:0] t_r29_c27_2;
  wire [7:0] t_r29_c27_3;
  wire [7:0] t_r29_c27_4;
  wire [7:0] t_r29_c27_5;
  wire [7:0] t_r29_c27_6;
  wire [7:0] t_r29_c27_7;
  wire [7:0] t_r29_c27_8;
  wire [7:0] t_r29_c27_9;
  wire [7:0] t_r29_c27_10;
  wire [7:0] t_r29_c27_11;
  wire [7:0] t_r29_c27_12;
  wire [7:0] t_r29_c28_0;
  wire [7:0] t_r29_c28_1;
  wire [7:0] t_r29_c28_2;
  wire [7:0] t_r29_c28_3;
  wire [7:0] t_r29_c28_4;
  wire [7:0] t_r29_c28_5;
  wire [7:0] t_r29_c28_6;
  wire [7:0] t_r29_c28_7;
  wire [7:0] t_r29_c28_8;
  wire [7:0] t_r29_c28_9;
  wire [7:0] t_r29_c28_10;
  wire [7:0] t_r29_c28_11;
  wire [7:0] t_r29_c28_12;
  wire [7:0] t_r29_c29_0;
  wire [7:0] t_r29_c29_1;
  wire [7:0] t_r29_c29_2;
  wire [7:0] t_r29_c29_3;
  wire [7:0] t_r29_c29_4;
  wire [7:0] t_r29_c29_5;
  wire [7:0] t_r29_c29_6;
  wire [7:0] t_r29_c29_7;
  wire [7:0] t_r29_c29_8;
  wire [7:0] t_r29_c29_9;
  wire [7:0] t_r29_c29_10;
  wire [7:0] t_r29_c29_11;
  wire [7:0] t_r29_c29_12;
  wire [7:0] t_r29_c30_0;
  wire [7:0] t_r29_c30_1;
  wire [7:0] t_r29_c30_2;
  wire [7:0] t_r29_c30_3;
  wire [7:0] t_r29_c30_4;
  wire [7:0] t_r29_c30_5;
  wire [7:0] t_r29_c30_6;
  wire [7:0] t_r29_c30_7;
  wire [7:0] t_r29_c30_8;
  wire [7:0] t_r29_c30_9;
  wire [7:0] t_r29_c30_10;
  wire [7:0] t_r29_c30_11;
  wire [7:0] t_r29_c30_12;
  wire [7:0] t_r29_c31_0;
  wire [7:0] t_r29_c31_1;
  wire [7:0] t_r29_c31_2;
  wire [7:0] t_r29_c31_3;
  wire [7:0] t_r29_c31_4;
  wire [7:0] t_r29_c31_5;
  wire [7:0] t_r29_c31_6;
  wire [7:0] t_r29_c31_7;
  wire [7:0] t_r29_c31_8;
  wire [7:0] t_r29_c31_9;
  wire [7:0] t_r29_c31_10;
  wire [7:0] t_r29_c31_11;
  wire [7:0] t_r29_c31_12;
  wire [7:0] t_r29_c32_0;
  wire [7:0] t_r29_c32_1;
  wire [7:0] t_r29_c32_2;
  wire [7:0] t_r29_c32_3;
  wire [7:0] t_r29_c32_4;
  wire [7:0] t_r29_c32_5;
  wire [7:0] t_r29_c32_6;
  wire [7:0] t_r29_c32_7;
  wire [7:0] t_r29_c32_8;
  wire [7:0] t_r29_c32_9;
  wire [7:0] t_r29_c32_10;
  wire [7:0] t_r29_c32_11;
  wire [7:0] t_r29_c32_12;
  wire [7:0] t_r29_c33_0;
  wire [7:0] t_r29_c33_1;
  wire [7:0] t_r29_c33_2;
  wire [7:0] t_r29_c33_3;
  wire [7:0] t_r29_c33_4;
  wire [7:0] t_r29_c33_5;
  wire [7:0] t_r29_c33_6;
  wire [7:0] t_r29_c33_7;
  wire [7:0] t_r29_c33_8;
  wire [7:0] t_r29_c33_9;
  wire [7:0] t_r29_c33_10;
  wire [7:0] t_r29_c33_11;
  wire [7:0] t_r29_c33_12;
  wire [7:0] t_r29_c34_0;
  wire [7:0] t_r29_c34_1;
  wire [7:0] t_r29_c34_2;
  wire [7:0] t_r29_c34_3;
  wire [7:0] t_r29_c34_4;
  wire [7:0] t_r29_c34_5;
  wire [7:0] t_r29_c34_6;
  wire [7:0] t_r29_c34_7;
  wire [7:0] t_r29_c34_8;
  wire [7:0] t_r29_c34_9;
  wire [7:0] t_r29_c34_10;
  wire [7:0] t_r29_c34_11;
  wire [7:0] t_r29_c34_12;
  wire [7:0] t_r29_c35_0;
  wire [7:0] t_r29_c35_1;
  wire [7:0] t_r29_c35_2;
  wire [7:0] t_r29_c35_3;
  wire [7:0] t_r29_c35_4;
  wire [7:0] t_r29_c35_5;
  wire [7:0] t_r29_c35_6;
  wire [7:0] t_r29_c35_7;
  wire [7:0] t_r29_c35_8;
  wire [7:0] t_r29_c35_9;
  wire [7:0] t_r29_c35_10;
  wire [7:0] t_r29_c35_11;
  wire [7:0] t_r29_c35_12;
  wire [7:0] t_r29_c36_0;
  wire [7:0] t_r29_c36_1;
  wire [7:0] t_r29_c36_2;
  wire [7:0] t_r29_c36_3;
  wire [7:0] t_r29_c36_4;
  wire [7:0] t_r29_c36_5;
  wire [7:0] t_r29_c36_6;
  wire [7:0] t_r29_c36_7;
  wire [7:0] t_r29_c36_8;
  wire [7:0] t_r29_c36_9;
  wire [7:0] t_r29_c36_10;
  wire [7:0] t_r29_c36_11;
  wire [7:0] t_r29_c36_12;
  wire [7:0] t_r29_c37_0;
  wire [7:0] t_r29_c37_1;
  wire [7:0] t_r29_c37_2;
  wire [7:0] t_r29_c37_3;
  wire [7:0] t_r29_c37_4;
  wire [7:0] t_r29_c37_5;
  wire [7:0] t_r29_c37_6;
  wire [7:0] t_r29_c37_7;
  wire [7:0] t_r29_c37_8;
  wire [7:0] t_r29_c37_9;
  wire [7:0] t_r29_c37_10;
  wire [7:0] t_r29_c37_11;
  wire [7:0] t_r29_c37_12;
  wire [7:0] t_r29_c38_0;
  wire [7:0] t_r29_c38_1;
  wire [7:0] t_r29_c38_2;
  wire [7:0] t_r29_c38_3;
  wire [7:0] t_r29_c38_4;
  wire [7:0] t_r29_c38_5;
  wire [7:0] t_r29_c38_6;
  wire [7:0] t_r29_c38_7;
  wire [7:0] t_r29_c38_8;
  wire [7:0] t_r29_c38_9;
  wire [7:0] t_r29_c38_10;
  wire [7:0] t_r29_c38_11;
  wire [7:0] t_r29_c38_12;
  wire [7:0] t_r29_c39_0;
  wire [7:0] t_r29_c39_1;
  wire [7:0] t_r29_c39_2;
  wire [7:0] t_r29_c39_3;
  wire [7:0] t_r29_c39_4;
  wire [7:0] t_r29_c39_5;
  wire [7:0] t_r29_c39_6;
  wire [7:0] t_r29_c39_7;
  wire [7:0] t_r29_c39_8;
  wire [7:0] t_r29_c39_9;
  wire [7:0] t_r29_c39_10;
  wire [7:0] t_r29_c39_11;
  wire [7:0] t_r29_c39_12;
  wire [7:0] t_r29_c40_0;
  wire [7:0] t_r29_c40_1;
  wire [7:0] t_r29_c40_2;
  wire [7:0] t_r29_c40_3;
  wire [7:0] t_r29_c40_4;
  wire [7:0] t_r29_c40_5;
  wire [7:0] t_r29_c40_6;
  wire [7:0] t_r29_c40_7;
  wire [7:0] t_r29_c40_8;
  wire [7:0] t_r29_c40_9;
  wire [7:0] t_r29_c40_10;
  wire [7:0] t_r29_c40_11;
  wire [7:0] t_r29_c40_12;
  wire [7:0] t_r29_c41_0;
  wire [7:0] t_r29_c41_1;
  wire [7:0] t_r29_c41_2;
  wire [7:0] t_r29_c41_3;
  wire [7:0] t_r29_c41_4;
  wire [7:0] t_r29_c41_5;
  wire [7:0] t_r29_c41_6;
  wire [7:0] t_r29_c41_7;
  wire [7:0] t_r29_c41_8;
  wire [7:0] t_r29_c41_9;
  wire [7:0] t_r29_c41_10;
  wire [7:0] t_r29_c41_11;
  wire [7:0] t_r29_c41_12;
  wire [7:0] t_r29_c42_0;
  wire [7:0] t_r29_c42_1;
  wire [7:0] t_r29_c42_2;
  wire [7:0] t_r29_c42_3;
  wire [7:0] t_r29_c42_4;
  wire [7:0] t_r29_c42_5;
  wire [7:0] t_r29_c42_6;
  wire [7:0] t_r29_c42_7;
  wire [7:0] t_r29_c42_8;
  wire [7:0] t_r29_c42_9;
  wire [7:0] t_r29_c42_10;
  wire [7:0] t_r29_c42_11;
  wire [7:0] t_r29_c42_12;
  wire [7:0] t_r29_c43_0;
  wire [7:0] t_r29_c43_1;
  wire [7:0] t_r29_c43_2;
  wire [7:0] t_r29_c43_3;
  wire [7:0] t_r29_c43_4;
  wire [7:0] t_r29_c43_5;
  wire [7:0] t_r29_c43_6;
  wire [7:0] t_r29_c43_7;
  wire [7:0] t_r29_c43_8;
  wire [7:0] t_r29_c43_9;
  wire [7:0] t_r29_c43_10;
  wire [7:0] t_r29_c43_11;
  wire [7:0] t_r29_c43_12;
  wire [7:0] t_r29_c44_0;
  wire [7:0] t_r29_c44_1;
  wire [7:0] t_r29_c44_2;
  wire [7:0] t_r29_c44_3;
  wire [7:0] t_r29_c44_4;
  wire [7:0] t_r29_c44_5;
  wire [7:0] t_r29_c44_6;
  wire [7:0] t_r29_c44_7;
  wire [7:0] t_r29_c44_8;
  wire [7:0] t_r29_c44_9;
  wire [7:0] t_r29_c44_10;
  wire [7:0] t_r29_c44_11;
  wire [7:0] t_r29_c44_12;
  wire [7:0] t_r29_c45_0;
  wire [7:0] t_r29_c45_1;
  wire [7:0] t_r29_c45_2;
  wire [7:0] t_r29_c45_3;
  wire [7:0] t_r29_c45_4;
  wire [7:0] t_r29_c45_5;
  wire [7:0] t_r29_c45_6;
  wire [7:0] t_r29_c45_7;
  wire [7:0] t_r29_c45_8;
  wire [7:0] t_r29_c45_9;
  wire [7:0] t_r29_c45_10;
  wire [7:0] t_r29_c45_11;
  wire [7:0] t_r29_c45_12;
  wire [7:0] t_r29_c46_0;
  wire [7:0] t_r29_c46_1;
  wire [7:0] t_r29_c46_2;
  wire [7:0] t_r29_c46_3;
  wire [7:0] t_r29_c46_4;
  wire [7:0] t_r29_c46_5;
  wire [7:0] t_r29_c46_6;
  wire [7:0] t_r29_c46_7;
  wire [7:0] t_r29_c46_8;
  wire [7:0] t_r29_c46_9;
  wire [7:0] t_r29_c46_10;
  wire [7:0] t_r29_c46_11;
  wire [7:0] t_r29_c46_12;
  wire [7:0] t_r29_c47_0;
  wire [7:0] t_r29_c47_1;
  wire [7:0] t_r29_c47_2;
  wire [7:0] t_r29_c47_3;
  wire [7:0] t_r29_c47_4;
  wire [7:0] t_r29_c47_5;
  wire [7:0] t_r29_c47_6;
  wire [7:0] t_r29_c47_7;
  wire [7:0] t_r29_c47_8;
  wire [7:0] t_r29_c47_9;
  wire [7:0] t_r29_c47_10;
  wire [7:0] t_r29_c47_11;
  wire [7:0] t_r29_c47_12;
  wire [7:0] t_r29_c48_0;
  wire [7:0] t_r29_c48_1;
  wire [7:0] t_r29_c48_2;
  wire [7:0] t_r29_c48_3;
  wire [7:0] t_r29_c48_4;
  wire [7:0] t_r29_c48_5;
  wire [7:0] t_r29_c48_6;
  wire [7:0] t_r29_c48_7;
  wire [7:0] t_r29_c48_8;
  wire [7:0] t_r29_c48_9;
  wire [7:0] t_r29_c48_10;
  wire [7:0] t_r29_c48_11;
  wire [7:0] t_r29_c48_12;
  wire [7:0] t_r29_c49_0;
  wire [7:0] t_r29_c49_1;
  wire [7:0] t_r29_c49_2;
  wire [7:0] t_r29_c49_3;
  wire [7:0] t_r29_c49_4;
  wire [7:0] t_r29_c49_5;
  wire [7:0] t_r29_c49_6;
  wire [7:0] t_r29_c49_7;
  wire [7:0] t_r29_c49_8;
  wire [7:0] t_r29_c49_9;
  wire [7:0] t_r29_c49_10;
  wire [7:0] t_r29_c49_11;
  wire [7:0] t_r29_c49_12;
  wire [7:0] t_r29_c50_0;
  wire [7:0] t_r29_c50_1;
  wire [7:0] t_r29_c50_2;
  wire [7:0] t_r29_c50_3;
  wire [7:0] t_r29_c50_4;
  wire [7:0] t_r29_c50_5;
  wire [7:0] t_r29_c50_6;
  wire [7:0] t_r29_c50_7;
  wire [7:0] t_r29_c50_8;
  wire [7:0] t_r29_c50_9;
  wire [7:0] t_r29_c50_10;
  wire [7:0] t_r29_c50_11;
  wire [7:0] t_r29_c50_12;
  wire [7:0] t_r29_c51_0;
  wire [7:0] t_r29_c51_1;
  wire [7:0] t_r29_c51_2;
  wire [7:0] t_r29_c51_3;
  wire [7:0] t_r29_c51_4;
  wire [7:0] t_r29_c51_5;
  wire [7:0] t_r29_c51_6;
  wire [7:0] t_r29_c51_7;
  wire [7:0] t_r29_c51_8;
  wire [7:0] t_r29_c51_9;
  wire [7:0] t_r29_c51_10;
  wire [7:0] t_r29_c51_11;
  wire [7:0] t_r29_c51_12;
  wire [7:0] t_r29_c52_0;
  wire [7:0] t_r29_c52_1;
  wire [7:0] t_r29_c52_2;
  wire [7:0] t_r29_c52_3;
  wire [7:0] t_r29_c52_4;
  wire [7:0] t_r29_c52_5;
  wire [7:0] t_r29_c52_6;
  wire [7:0] t_r29_c52_7;
  wire [7:0] t_r29_c52_8;
  wire [7:0] t_r29_c52_9;
  wire [7:0] t_r29_c52_10;
  wire [7:0] t_r29_c52_11;
  wire [7:0] t_r29_c52_12;
  wire [7:0] t_r29_c53_0;
  wire [7:0] t_r29_c53_1;
  wire [7:0] t_r29_c53_2;
  wire [7:0] t_r29_c53_3;
  wire [7:0] t_r29_c53_4;
  wire [7:0] t_r29_c53_5;
  wire [7:0] t_r29_c53_6;
  wire [7:0] t_r29_c53_7;
  wire [7:0] t_r29_c53_8;
  wire [7:0] t_r29_c53_9;
  wire [7:0] t_r29_c53_10;
  wire [7:0] t_r29_c53_11;
  wire [7:0] t_r29_c53_12;
  wire [7:0] t_r29_c54_0;
  wire [7:0] t_r29_c54_1;
  wire [7:0] t_r29_c54_2;
  wire [7:0] t_r29_c54_3;
  wire [7:0] t_r29_c54_4;
  wire [7:0] t_r29_c54_5;
  wire [7:0] t_r29_c54_6;
  wire [7:0] t_r29_c54_7;
  wire [7:0] t_r29_c54_8;
  wire [7:0] t_r29_c54_9;
  wire [7:0] t_r29_c54_10;
  wire [7:0] t_r29_c54_11;
  wire [7:0] t_r29_c54_12;
  wire [7:0] t_r29_c55_0;
  wire [7:0] t_r29_c55_1;
  wire [7:0] t_r29_c55_2;
  wire [7:0] t_r29_c55_3;
  wire [7:0] t_r29_c55_4;
  wire [7:0] t_r29_c55_5;
  wire [7:0] t_r29_c55_6;
  wire [7:0] t_r29_c55_7;
  wire [7:0] t_r29_c55_8;
  wire [7:0] t_r29_c55_9;
  wire [7:0] t_r29_c55_10;
  wire [7:0] t_r29_c55_11;
  wire [7:0] t_r29_c55_12;
  wire [7:0] t_r29_c56_0;
  wire [7:0] t_r29_c56_1;
  wire [7:0] t_r29_c56_2;
  wire [7:0] t_r29_c56_3;
  wire [7:0] t_r29_c56_4;
  wire [7:0] t_r29_c56_5;
  wire [7:0] t_r29_c56_6;
  wire [7:0] t_r29_c56_7;
  wire [7:0] t_r29_c56_8;
  wire [7:0] t_r29_c56_9;
  wire [7:0] t_r29_c56_10;
  wire [7:0] t_r29_c56_11;
  wire [7:0] t_r29_c56_12;
  wire [7:0] t_r29_c57_0;
  wire [7:0] t_r29_c57_1;
  wire [7:0] t_r29_c57_2;
  wire [7:0] t_r29_c57_3;
  wire [7:0] t_r29_c57_4;
  wire [7:0] t_r29_c57_5;
  wire [7:0] t_r29_c57_6;
  wire [7:0] t_r29_c57_7;
  wire [7:0] t_r29_c57_8;
  wire [7:0] t_r29_c57_9;
  wire [7:0] t_r29_c57_10;
  wire [7:0] t_r29_c57_11;
  wire [7:0] t_r29_c57_12;
  wire [7:0] t_r29_c58_0;
  wire [7:0] t_r29_c58_1;
  wire [7:0] t_r29_c58_2;
  wire [7:0] t_r29_c58_3;
  wire [7:0] t_r29_c58_4;
  wire [7:0] t_r29_c58_5;
  wire [7:0] t_r29_c58_6;
  wire [7:0] t_r29_c58_7;
  wire [7:0] t_r29_c58_8;
  wire [7:0] t_r29_c58_9;
  wire [7:0] t_r29_c58_10;
  wire [7:0] t_r29_c58_11;
  wire [7:0] t_r29_c58_12;
  wire [7:0] t_r29_c59_0;
  wire [7:0] t_r29_c59_1;
  wire [7:0] t_r29_c59_2;
  wire [7:0] t_r29_c59_3;
  wire [7:0] t_r29_c59_4;
  wire [7:0] t_r29_c59_5;
  wire [7:0] t_r29_c59_6;
  wire [7:0] t_r29_c59_7;
  wire [7:0] t_r29_c59_8;
  wire [7:0] t_r29_c59_9;
  wire [7:0] t_r29_c59_10;
  wire [7:0] t_r29_c59_11;
  wire [7:0] t_r29_c59_12;
  wire [7:0] t_r29_c60_0;
  wire [7:0] t_r29_c60_1;
  wire [7:0] t_r29_c60_2;
  wire [7:0] t_r29_c60_3;
  wire [7:0] t_r29_c60_4;
  wire [7:0] t_r29_c60_5;
  wire [7:0] t_r29_c60_6;
  wire [7:0] t_r29_c60_7;
  wire [7:0] t_r29_c60_8;
  wire [7:0] t_r29_c60_9;
  wire [7:0] t_r29_c60_10;
  wire [7:0] t_r29_c60_11;
  wire [7:0] t_r29_c60_12;
  wire [7:0] t_r29_c61_0;
  wire [7:0] t_r29_c61_1;
  wire [7:0] t_r29_c61_2;
  wire [7:0] t_r29_c61_3;
  wire [7:0] t_r29_c61_4;
  wire [7:0] t_r29_c61_5;
  wire [7:0] t_r29_c61_6;
  wire [7:0] t_r29_c61_7;
  wire [7:0] t_r29_c61_8;
  wire [7:0] t_r29_c61_9;
  wire [7:0] t_r29_c61_10;
  wire [7:0] t_r29_c61_11;
  wire [7:0] t_r29_c61_12;
  wire [7:0] t_r29_c62_0;
  wire [7:0] t_r29_c62_1;
  wire [7:0] t_r29_c62_2;
  wire [7:0] t_r29_c62_3;
  wire [7:0] t_r29_c62_4;
  wire [7:0] t_r29_c62_5;
  wire [7:0] t_r29_c62_6;
  wire [7:0] t_r29_c62_7;
  wire [7:0] t_r29_c62_8;
  wire [7:0] t_r29_c62_9;
  wire [7:0] t_r29_c62_10;
  wire [7:0] t_r29_c62_11;
  wire [7:0] t_r29_c62_12;
  wire [7:0] t_r29_c63_0;
  wire [7:0] t_r29_c63_1;
  wire [7:0] t_r29_c63_2;
  wire [7:0] t_r29_c63_3;
  wire [7:0] t_r29_c63_4;
  wire [7:0] t_r29_c63_5;
  wire [7:0] t_r29_c63_6;
  wire [7:0] t_r29_c63_7;
  wire [7:0] t_r29_c63_8;
  wire [7:0] t_r29_c63_9;
  wire [7:0] t_r29_c63_10;
  wire [7:0] t_r29_c63_11;
  wire [7:0] t_r29_c63_12;
  wire [7:0] t_r29_c64_0;
  wire [7:0] t_r29_c64_1;
  wire [7:0] t_r29_c64_2;
  wire [7:0] t_r29_c64_3;
  wire [7:0] t_r29_c64_4;
  wire [7:0] t_r29_c64_5;
  wire [7:0] t_r29_c64_6;
  wire [7:0] t_r29_c64_7;
  wire [7:0] t_r29_c64_8;
  wire [7:0] t_r29_c64_9;
  wire [7:0] t_r29_c64_10;
  wire [7:0] t_r29_c64_11;
  wire [7:0] t_r29_c64_12;
  wire [7:0] t_r29_c65_0;
  wire [7:0] t_r29_c65_1;
  wire [7:0] t_r29_c65_2;
  wire [7:0] t_r29_c65_3;
  wire [7:0] t_r29_c65_4;
  wire [7:0] t_r29_c65_5;
  wire [7:0] t_r29_c65_6;
  wire [7:0] t_r29_c65_7;
  wire [7:0] t_r29_c65_8;
  wire [7:0] t_r29_c65_9;
  wire [7:0] t_r29_c65_10;
  wire [7:0] t_r29_c65_11;
  wire [7:0] t_r29_c65_12;
  wire [7:0] t_r30_c0_0;
  wire [7:0] t_r30_c0_1;
  wire [7:0] t_r30_c0_2;
  wire [7:0] t_r30_c0_3;
  wire [7:0] t_r30_c0_4;
  wire [7:0] t_r30_c0_5;
  wire [7:0] t_r30_c0_6;
  wire [7:0] t_r30_c0_7;
  wire [7:0] t_r30_c0_8;
  wire [7:0] t_r30_c0_9;
  wire [7:0] t_r30_c0_10;
  wire [7:0] t_r30_c0_11;
  wire [7:0] t_r30_c0_12;
  wire [7:0] t_r30_c1_0;
  wire [7:0] t_r30_c1_1;
  wire [7:0] t_r30_c1_2;
  wire [7:0] t_r30_c1_3;
  wire [7:0] t_r30_c1_4;
  wire [7:0] t_r30_c1_5;
  wire [7:0] t_r30_c1_6;
  wire [7:0] t_r30_c1_7;
  wire [7:0] t_r30_c1_8;
  wire [7:0] t_r30_c1_9;
  wire [7:0] t_r30_c1_10;
  wire [7:0] t_r30_c1_11;
  wire [7:0] t_r30_c1_12;
  wire [7:0] t_r30_c2_0;
  wire [7:0] t_r30_c2_1;
  wire [7:0] t_r30_c2_2;
  wire [7:0] t_r30_c2_3;
  wire [7:0] t_r30_c2_4;
  wire [7:0] t_r30_c2_5;
  wire [7:0] t_r30_c2_6;
  wire [7:0] t_r30_c2_7;
  wire [7:0] t_r30_c2_8;
  wire [7:0] t_r30_c2_9;
  wire [7:0] t_r30_c2_10;
  wire [7:0] t_r30_c2_11;
  wire [7:0] t_r30_c2_12;
  wire [7:0] t_r30_c3_0;
  wire [7:0] t_r30_c3_1;
  wire [7:0] t_r30_c3_2;
  wire [7:0] t_r30_c3_3;
  wire [7:0] t_r30_c3_4;
  wire [7:0] t_r30_c3_5;
  wire [7:0] t_r30_c3_6;
  wire [7:0] t_r30_c3_7;
  wire [7:0] t_r30_c3_8;
  wire [7:0] t_r30_c3_9;
  wire [7:0] t_r30_c3_10;
  wire [7:0] t_r30_c3_11;
  wire [7:0] t_r30_c3_12;
  wire [7:0] t_r30_c4_0;
  wire [7:0] t_r30_c4_1;
  wire [7:0] t_r30_c4_2;
  wire [7:0] t_r30_c4_3;
  wire [7:0] t_r30_c4_4;
  wire [7:0] t_r30_c4_5;
  wire [7:0] t_r30_c4_6;
  wire [7:0] t_r30_c4_7;
  wire [7:0] t_r30_c4_8;
  wire [7:0] t_r30_c4_9;
  wire [7:0] t_r30_c4_10;
  wire [7:0] t_r30_c4_11;
  wire [7:0] t_r30_c4_12;
  wire [7:0] t_r30_c5_0;
  wire [7:0] t_r30_c5_1;
  wire [7:0] t_r30_c5_2;
  wire [7:0] t_r30_c5_3;
  wire [7:0] t_r30_c5_4;
  wire [7:0] t_r30_c5_5;
  wire [7:0] t_r30_c5_6;
  wire [7:0] t_r30_c5_7;
  wire [7:0] t_r30_c5_8;
  wire [7:0] t_r30_c5_9;
  wire [7:0] t_r30_c5_10;
  wire [7:0] t_r30_c5_11;
  wire [7:0] t_r30_c5_12;
  wire [7:0] t_r30_c6_0;
  wire [7:0] t_r30_c6_1;
  wire [7:0] t_r30_c6_2;
  wire [7:0] t_r30_c6_3;
  wire [7:0] t_r30_c6_4;
  wire [7:0] t_r30_c6_5;
  wire [7:0] t_r30_c6_6;
  wire [7:0] t_r30_c6_7;
  wire [7:0] t_r30_c6_8;
  wire [7:0] t_r30_c6_9;
  wire [7:0] t_r30_c6_10;
  wire [7:0] t_r30_c6_11;
  wire [7:0] t_r30_c6_12;
  wire [7:0] t_r30_c7_0;
  wire [7:0] t_r30_c7_1;
  wire [7:0] t_r30_c7_2;
  wire [7:0] t_r30_c7_3;
  wire [7:0] t_r30_c7_4;
  wire [7:0] t_r30_c7_5;
  wire [7:0] t_r30_c7_6;
  wire [7:0] t_r30_c7_7;
  wire [7:0] t_r30_c7_8;
  wire [7:0] t_r30_c7_9;
  wire [7:0] t_r30_c7_10;
  wire [7:0] t_r30_c7_11;
  wire [7:0] t_r30_c7_12;
  wire [7:0] t_r30_c8_0;
  wire [7:0] t_r30_c8_1;
  wire [7:0] t_r30_c8_2;
  wire [7:0] t_r30_c8_3;
  wire [7:0] t_r30_c8_4;
  wire [7:0] t_r30_c8_5;
  wire [7:0] t_r30_c8_6;
  wire [7:0] t_r30_c8_7;
  wire [7:0] t_r30_c8_8;
  wire [7:0] t_r30_c8_9;
  wire [7:0] t_r30_c8_10;
  wire [7:0] t_r30_c8_11;
  wire [7:0] t_r30_c8_12;
  wire [7:0] t_r30_c9_0;
  wire [7:0] t_r30_c9_1;
  wire [7:0] t_r30_c9_2;
  wire [7:0] t_r30_c9_3;
  wire [7:0] t_r30_c9_4;
  wire [7:0] t_r30_c9_5;
  wire [7:0] t_r30_c9_6;
  wire [7:0] t_r30_c9_7;
  wire [7:0] t_r30_c9_8;
  wire [7:0] t_r30_c9_9;
  wire [7:0] t_r30_c9_10;
  wire [7:0] t_r30_c9_11;
  wire [7:0] t_r30_c9_12;
  wire [7:0] t_r30_c10_0;
  wire [7:0] t_r30_c10_1;
  wire [7:0] t_r30_c10_2;
  wire [7:0] t_r30_c10_3;
  wire [7:0] t_r30_c10_4;
  wire [7:0] t_r30_c10_5;
  wire [7:0] t_r30_c10_6;
  wire [7:0] t_r30_c10_7;
  wire [7:0] t_r30_c10_8;
  wire [7:0] t_r30_c10_9;
  wire [7:0] t_r30_c10_10;
  wire [7:0] t_r30_c10_11;
  wire [7:0] t_r30_c10_12;
  wire [7:0] t_r30_c11_0;
  wire [7:0] t_r30_c11_1;
  wire [7:0] t_r30_c11_2;
  wire [7:0] t_r30_c11_3;
  wire [7:0] t_r30_c11_4;
  wire [7:0] t_r30_c11_5;
  wire [7:0] t_r30_c11_6;
  wire [7:0] t_r30_c11_7;
  wire [7:0] t_r30_c11_8;
  wire [7:0] t_r30_c11_9;
  wire [7:0] t_r30_c11_10;
  wire [7:0] t_r30_c11_11;
  wire [7:0] t_r30_c11_12;
  wire [7:0] t_r30_c12_0;
  wire [7:0] t_r30_c12_1;
  wire [7:0] t_r30_c12_2;
  wire [7:0] t_r30_c12_3;
  wire [7:0] t_r30_c12_4;
  wire [7:0] t_r30_c12_5;
  wire [7:0] t_r30_c12_6;
  wire [7:0] t_r30_c12_7;
  wire [7:0] t_r30_c12_8;
  wire [7:0] t_r30_c12_9;
  wire [7:0] t_r30_c12_10;
  wire [7:0] t_r30_c12_11;
  wire [7:0] t_r30_c12_12;
  wire [7:0] t_r30_c13_0;
  wire [7:0] t_r30_c13_1;
  wire [7:0] t_r30_c13_2;
  wire [7:0] t_r30_c13_3;
  wire [7:0] t_r30_c13_4;
  wire [7:0] t_r30_c13_5;
  wire [7:0] t_r30_c13_6;
  wire [7:0] t_r30_c13_7;
  wire [7:0] t_r30_c13_8;
  wire [7:0] t_r30_c13_9;
  wire [7:0] t_r30_c13_10;
  wire [7:0] t_r30_c13_11;
  wire [7:0] t_r30_c13_12;
  wire [7:0] t_r30_c14_0;
  wire [7:0] t_r30_c14_1;
  wire [7:0] t_r30_c14_2;
  wire [7:0] t_r30_c14_3;
  wire [7:0] t_r30_c14_4;
  wire [7:0] t_r30_c14_5;
  wire [7:0] t_r30_c14_6;
  wire [7:0] t_r30_c14_7;
  wire [7:0] t_r30_c14_8;
  wire [7:0] t_r30_c14_9;
  wire [7:0] t_r30_c14_10;
  wire [7:0] t_r30_c14_11;
  wire [7:0] t_r30_c14_12;
  wire [7:0] t_r30_c15_0;
  wire [7:0] t_r30_c15_1;
  wire [7:0] t_r30_c15_2;
  wire [7:0] t_r30_c15_3;
  wire [7:0] t_r30_c15_4;
  wire [7:0] t_r30_c15_5;
  wire [7:0] t_r30_c15_6;
  wire [7:0] t_r30_c15_7;
  wire [7:0] t_r30_c15_8;
  wire [7:0] t_r30_c15_9;
  wire [7:0] t_r30_c15_10;
  wire [7:0] t_r30_c15_11;
  wire [7:0] t_r30_c15_12;
  wire [7:0] t_r30_c16_0;
  wire [7:0] t_r30_c16_1;
  wire [7:0] t_r30_c16_2;
  wire [7:0] t_r30_c16_3;
  wire [7:0] t_r30_c16_4;
  wire [7:0] t_r30_c16_5;
  wire [7:0] t_r30_c16_6;
  wire [7:0] t_r30_c16_7;
  wire [7:0] t_r30_c16_8;
  wire [7:0] t_r30_c16_9;
  wire [7:0] t_r30_c16_10;
  wire [7:0] t_r30_c16_11;
  wire [7:0] t_r30_c16_12;
  wire [7:0] t_r30_c17_0;
  wire [7:0] t_r30_c17_1;
  wire [7:0] t_r30_c17_2;
  wire [7:0] t_r30_c17_3;
  wire [7:0] t_r30_c17_4;
  wire [7:0] t_r30_c17_5;
  wire [7:0] t_r30_c17_6;
  wire [7:0] t_r30_c17_7;
  wire [7:0] t_r30_c17_8;
  wire [7:0] t_r30_c17_9;
  wire [7:0] t_r30_c17_10;
  wire [7:0] t_r30_c17_11;
  wire [7:0] t_r30_c17_12;
  wire [7:0] t_r30_c18_0;
  wire [7:0] t_r30_c18_1;
  wire [7:0] t_r30_c18_2;
  wire [7:0] t_r30_c18_3;
  wire [7:0] t_r30_c18_4;
  wire [7:0] t_r30_c18_5;
  wire [7:0] t_r30_c18_6;
  wire [7:0] t_r30_c18_7;
  wire [7:0] t_r30_c18_8;
  wire [7:0] t_r30_c18_9;
  wire [7:0] t_r30_c18_10;
  wire [7:0] t_r30_c18_11;
  wire [7:0] t_r30_c18_12;
  wire [7:0] t_r30_c19_0;
  wire [7:0] t_r30_c19_1;
  wire [7:0] t_r30_c19_2;
  wire [7:0] t_r30_c19_3;
  wire [7:0] t_r30_c19_4;
  wire [7:0] t_r30_c19_5;
  wire [7:0] t_r30_c19_6;
  wire [7:0] t_r30_c19_7;
  wire [7:0] t_r30_c19_8;
  wire [7:0] t_r30_c19_9;
  wire [7:0] t_r30_c19_10;
  wire [7:0] t_r30_c19_11;
  wire [7:0] t_r30_c19_12;
  wire [7:0] t_r30_c20_0;
  wire [7:0] t_r30_c20_1;
  wire [7:0] t_r30_c20_2;
  wire [7:0] t_r30_c20_3;
  wire [7:0] t_r30_c20_4;
  wire [7:0] t_r30_c20_5;
  wire [7:0] t_r30_c20_6;
  wire [7:0] t_r30_c20_7;
  wire [7:0] t_r30_c20_8;
  wire [7:0] t_r30_c20_9;
  wire [7:0] t_r30_c20_10;
  wire [7:0] t_r30_c20_11;
  wire [7:0] t_r30_c20_12;
  wire [7:0] t_r30_c21_0;
  wire [7:0] t_r30_c21_1;
  wire [7:0] t_r30_c21_2;
  wire [7:0] t_r30_c21_3;
  wire [7:0] t_r30_c21_4;
  wire [7:0] t_r30_c21_5;
  wire [7:0] t_r30_c21_6;
  wire [7:0] t_r30_c21_7;
  wire [7:0] t_r30_c21_8;
  wire [7:0] t_r30_c21_9;
  wire [7:0] t_r30_c21_10;
  wire [7:0] t_r30_c21_11;
  wire [7:0] t_r30_c21_12;
  wire [7:0] t_r30_c22_0;
  wire [7:0] t_r30_c22_1;
  wire [7:0] t_r30_c22_2;
  wire [7:0] t_r30_c22_3;
  wire [7:0] t_r30_c22_4;
  wire [7:0] t_r30_c22_5;
  wire [7:0] t_r30_c22_6;
  wire [7:0] t_r30_c22_7;
  wire [7:0] t_r30_c22_8;
  wire [7:0] t_r30_c22_9;
  wire [7:0] t_r30_c22_10;
  wire [7:0] t_r30_c22_11;
  wire [7:0] t_r30_c22_12;
  wire [7:0] t_r30_c23_0;
  wire [7:0] t_r30_c23_1;
  wire [7:0] t_r30_c23_2;
  wire [7:0] t_r30_c23_3;
  wire [7:0] t_r30_c23_4;
  wire [7:0] t_r30_c23_5;
  wire [7:0] t_r30_c23_6;
  wire [7:0] t_r30_c23_7;
  wire [7:0] t_r30_c23_8;
  wire [7:0] t_r30_c23_9;
  wire [7:0] t_r30_c23_10;
  wire [7:0] t_r30_c23_11;
  wire [7:0] t_r30_c23_12;
  wire [7:0] t_r30_c24_0;
  wire [7:0] t_r30_c24_1;
  wire [7:0] t_r30_c24_2;
  wire [7:0] t_r30_c24_3;
  wire [7:0] t_r30_c24_4;
  wire [7:0] t_r30_c24_5;
  wire [7:0] t_r30_c24_6;
  wire [7:0] t_r30_c24_7;
  wire [7:0] t_r30_c24_8;
  wire [7:0] t_r30_c24_9;
  wire [7:0] t_r30_c24_10;
  wire [7:0] t_r30_c24_11;
  wire [7:0] t_r30_c24_12;
  wire [7:0] t_r30_c25_0;
  wire [7:0] t_r30_c25_1;
  wire [7:0] t_r30_c25_2;
  wire [7:0] t_r30_c25_3;
  wire [7:0] t_r30_c25_4;
  wire [7:0] t_r30_c25_5;
  wire [7:0] t_r30_c25_6;
  wire [7:0] t_r30_c25_7;
  wire [7:0] t_r30_c25_8;
  wire [7:0] t_r30_c25_9;
  wire [7:0] t_r30_c25_10;
  wire [7:0] t_r30_c25_11;
  wire [7:0] t_r30_c25_12;
  wire [7:0] t_r30_c26_0;
  wire [7:0] t_r30_c26_1;
  wire [7:0] t_r30_c26_2;
  wire [7:0] t_r30_c26_3;
  wire [7:0] t_r30_c26_4;
  wire [7:0] t_r30_c26_5;
  wire [7:0] t_r30_c26_6;
  wire [7:0] t_r30_c26_7;
  wire [7:0] t_r30_c26_8;
  wire [7:0] t_r30_c26_9;
  wire [7:0] t_r30_c26_10;
  wire [7:0] t_r30_c26_11;
  wire [7:0] t_r30_c26_12;
  wire [7:0] t_r30_c27_0;
  wire [7:0] t_r30_c27_1;
  wire [7:0] t_r30_c27_2;
  wire [7:0] t_r30_c27_3;
  wire [7:0] t_r30_c27_4;
  wire [7:0] t_r30_c27_5;
  wire [7:0] t_r30_c27_6;
  wire [7:0] t_r30_c27_7;
  wire [7:0] t_r30_c27_8;
  wire [7:0] t_r30_c27_9;
  wire [7:0] t_r30_c27_10;
  wire [7:0] t_r30_c27_11;
  wire [7:0] t_r30_c27_12;
  wire [7:0] t_r30_c28_0;
  wire [7:0] t_r30_c28_1;
  wire [7:0] t_r30_c28_2;
  wire [7:0] t_r30_c28_3;
  wire [7:0] t_r30_c28_4;
  wire [7:0] t_r30_c28_5;
  wire [7:0] t_r30_c28_6;
  wire [7:0] t_r30_c28_7;
  wire [7:0] t_r30_c28_8;
  wire [7:0] t_r30_c28_9;
  wire [7:0] t_r30_c28_10;
  wire [7:0] t_r30_c28_11;
  wire [7:0] t_r30_c28_12;
  wire [7:0] t_r30_c29_0;
  wire [7:0] t_r30_c29_1;
  wire [7:0] t_r30_c29_2;
  wire [7:0] t_r30_c29_3;
  wire [7:0] t_r30_c29_4;
  wire [7:0] t_r30_c29_5;
  wire [7:0] t_r30_c29_6;
  wire [7:0] t_r30_c29_7;
  wire [7:0] t_r30_c29_8;
  wire [7:0] t_r30_c29_9;
  wire [7:0] t_r30_c29_10;
  wire [7:0] t_r30_c29_11;
  wire [7:0] t_r30_c29_12;
  wire [7:0] t_r30_c30_0;
  wire [7:0] t_r30_c30_1;
  wire [7:0] t_r30_c30_2;
  wire [7:0] t_r30_c30_3;
  wire [7:0] t_r30_c30_4;
  wire [7:0] t_r30_c30_5;
  wire [7:0] t_r30_c30_6;
  wire [7:0] t_r30_c30_7;
  wire [7:0] t_r30_c30_8;
  wire [7:0] t_r30_c30_9;
  wire [7:0] t_r30_c30_10;
  wire [7:0] t_r30_c30_11;
  wire [7:0] t_r30_c30_12;
  wire [7:0] t_r30_c31_0;
  wire [7:0] t_r30_c31_1;
  wire [7:0] t_r30_c31_2;
  wire [7:0] t_r30_c31_3;
  wire [7:0] t_r30_c31_4;
  wire [7:0] t_r30_c31_5;
  wire [7:0] t_r30_c31_6;
  wire [7:0] t_r30_c31_7;
  wire [7:0] t_r30_c31_8;
  wire [7:0] t_r30_c31_9;
  wire [7:0] t_r30_c31_10;
  wire [7:0] t_r30_c31_11;
  wire [7:0] t_r30_c31_12;
  wire [7:0] t_r30_c32_0;
  wire [7:0] t_r30_c32_1;
  wire [7:0] t_r30_c32_2;
  wire [7:0] t_r30_c32_3;
  wire [7:0] t_r30_c32_4;
  wire [7:0] t_r30_c32_5;
  wire [7:0] t_r30_c32_6;
  wire [7:0] t_r30_c32_7;
  wire [7:0] t_r30_c32_8;
  wire [7:0] t_r30_c32_9;
  wire [7:0] t_r30_c32_10;
  wire [7:0] t_r30_c32_11;
  wire [7:0] t_r30_c32_12;
  wire [7:0] t_r30_c33_0;
  wire [7:0] t_r30_c33_1;
  wire [7:0] t_r30_c33_2;
  wire [7:0] t_r30_c33_3;
  wire [7:0] t_r30_c33_4;
  wire [7:0] t_r30_c33_5;
  wire [7:0] t_r30_c33_6;
  wire [7:0] t_r30_c33_7;
  wire [7:0] t_r30_c33_8;
  wire [7:0] t_r30_c33_9;
  wire [7:0] t_r30_c33_10;
  wire [7:0] t_r30_c33_11;
  wire [7:0] t_r30_c33_12;
  wire [7:0] t_r30_c34_0;
  wire [7:0] t_r30_c34_1;
  wire [7:0] t_r30_c34_2;
  wire [7:0] t_r30_c34_3;
  wire [7:0] t_r30_c34_4;
  wire [7:0] t_r30_c34_5;
  wire [7:0] t_r30_c34_6;
  wire [7:0] t_r30_c34_7;
  wire [7:0] t_r30_c34_8;
  wire [7:0] t_r30_c34_9;
  wire [7:0] t_r30_c34_10;
  wire [7:0] t_r30_c34_11;
  wire [7:0] t_r30_c34_12;
  wire [7:0] t_r30_c35_0;
  wire [7:0] t_r30_c35_1;
  wire [7:0] t_r30_c35_2;
  wire [7:0] t_r30_c35_3;
  wire [7:0] t_r30_c35_4;
  wire [7:0] t_r30_c35_5;
  wire [7:0] t_r30_c35_6;
  wire [7:0] t_r30_c35_7;
  wire [7:0] t_r30_c35_8;
  wire [7:0] t_r30_c35_9;
  wire [7:0] t_r30_c35_10;
  wire [7:0] t_r30_c35_11;
  wire [7:0] t_r30_c35_12;
  wire [7:0] t_r30_c36_0;
  wire [7:0] t_r30_c36_1;
  wire [7:0] t_r30_c36_2;
  wire [7:0] t_r30_c36_3;
  wire [7:0] t_r30_c36_4;
  wire [7:0] t_r30_c36_5;
  wire [7:0] t_r30_c36_6;
  wire [7:0] t_r30_c36_7;
  wire [7:0] t_r30_c36_8;
  wire [7:0] t_r30_c36_9;
  wire [7:0] t_r30_c36_10;
  wire [7:0] t_r30_c36_11;
  wire [7:0] t_r30_c36_12;
  wire [7:0] t_r30_c37_0;
  wire [7:0] t_r30_c37_1;
  wire [7:0] t_r30_c37_2;
  wire [7:0] t_r30_c37_3;
  wire [7:0] t_r30_c37_4;
  wire [7:0] t_r30_c37_5;
  wire [7:0] t_r30_c37_6;
  wire [7:0] t_r30_c37_7;
  wire [7:0] t_r30_c37_8;
  wire [7:0] t_r30_c37_9;
  wire [7:0] t_r30_c37_10;
  wire [7:0] t_r30_c37_11;
  wire [7:0] t_r30_c37_12;
  wire [7:0] t_r30_c38_0;
  wire [7:0] t_r30_c38_1;
  wire [7:0] t_r30_c38_2;
  wire [7:0] t_r30_c38_3;
  wire [7:0] t_r30_c38_4;
  wire [7:0] t_r30_c38_5;
  wire [7:0] t_r30_c38_6;
  wire [7:0] t_r30_c38_7;
  wire [7:0] t_r30_c38_8;
  wire [7:0] t_r30_c38_9;
  wire [7:0] t_r30_c38_10;
  wire [7:0] t_r30_c38_11;
  wire [7:0] t_r30_c38_12;
  wire [7:0] t_r30_c39_0;
  wire [7:0] t_r30_c39_1;
  wire [7:0] t_r30_c39_2;
  wire [7:0] t_r30_c39_3;
  wire [7:0] t_r30_c39_4;
  wire [7:0] t_r30_c39_5;
  wire [7:0] t_r30_c39_6;
  wire [7:0] t_r30_c39_7;
  wire [7:0] t_r30_c39_8;
  wire [7:0] t_r30_c39_9;
  wire [7:0] t_r30_c39_10;
  wire [7:0] t_r30_c39_11;
  wire [7:0] t_r30_c39_12;
  wire [7:0] t_r30_c40_0;
  wire [7:0] t_r30_c40_1;
  wire [7:0] t_r30_c40_2;
  wire [7:0] t_r30_c40_3;
  wire [7:0] t_r30_c40_4;
  wire [7:0] t_r30_c40_5;
  wire [7:0] t_r30_c40_6;
  wire [7:0] t_r30_c40_7;
  wire [7:0] t_r30_c40_8;
  wire [7:0] t_r30_c40_9;
  wire [7:0] t_r30_c40_10;
  wire [7:0] t_r30_c40_11;
  wire [7:0] t_r30_c40_12;
  wire [7:0] t_r30_c41_0;
  wire [7:0] t_r30_c41_1;
  wire [7:0] t_r30_c41_2;
  wire [7:0] t_r30_c41_3;
  wire [7:0] t_r30_c41_4;
  wire [7:0] t_r30_c41_5;
  wire [7:0] t_r30_c41_6;
  wire [7:0] t_r30_c41_7;
  wire [7:0] t_r30_c41_8;
  wire [7:0] t_r30_c41_9;
  wire [7:0] t_r30_c41_10;
  wire [7:0] t_r30_c41_11;
  wire [7:0] t_r30_c41_12;
  wire [7:0] t_r30_c42_0;
  wire [7:0] t_r30_c42_1;
  wire [7:0] t_r30_c42_2;
  wire [7:0] t_r30_c42_3;
  wire [7:0] t_r30_c42_4;
  wire [7:0] t_r30_c42_5;
  wire [7:0] t_r30_c42_6;
  wire [7:0] t_r30_c42_7;
  wire [7:0] t_r30_c42_8;
  wire [7:0] t_r30_c42_9;
  wire [7:0] t_r30_c42_10;
  wire [7:0] t_r30_c42_11;
  wire [7:0] t_r30_c42_12;
  wire [7:0] t_r30_c43_0;
  wire [7:0] t_r30_c43_1;
  wire [7:0] t_r30_c43_2;
  wire [7:0] t_r30_c43_3;
  wire [7:0] t_r30_c43_4;
  wire [7:0] t_r30_c43_5;
  wire [7:0] t_r30_c43_6;
  wire [7:0] t_r30_c43_7;
  wire [7:0] t_r30_c43_8;
  wire [7:0] t_r30_c43_9;
  wire [7:0] t_r30_c43_10;
  wire [7:0] t_r30_c43_11;
  wire [7:0] t_r30_c43_12;
  wire [7:0] t_r30_c44_0;
  wire [7:0] t_r30_c44_1;
  wire [7:0] t_r30_c44_2;
  wire [7:0] t_r30_c44_3;
  wire [7:0] t_r30_c44_4;
  wire [7:0] t_r30_c44_5;
  wire [7:0] t_r30_c44_6;
  wire [7:0] t_r30_c44_7;
  wire [7:0] t_r30_c44_8;
  wire [7:0] t_r30_c44_9;
  wire [7:0] t_r30_c44_10;
  wire [7:0] t_r30_c44_11;
  wire [7:0] t_r30_c44_12;
  wire [7:0] t_r30_c45_0;
  wire [7:0] t_r30_c45_1;
  wire [7:0] t_r30_c45_2;
  wire [7:0] t_r30_c45_3;
  wire [7:0] t_r30_c45_4;
  wire [7:0] t_r30_c45_5;
  wire [7:0] t_r30_c45_6;
  wire [7:0] t_r30_c45_7;
  wire [7:0] t_r30_c45_8;
  wire [7:0] t_r30_c45_9;
  wire [7:0] t_r30_c45_10;
  wire [7:0] t_r30_c45_11;
  wire [7:0] t_r30_c45_12;
  wire [7:0] t_r30_c46_0;
  wire [7:0] t_r30_c46_1;
  wire [7:0] t_r30_c46_2;
  wire [7:0] t_r30_c46_3;
  wire [7:0] t_r30_c46_4;
  wire [7:0] t_r30_c46_5;
  wire [7:0] t_r30_c46_6;
  wire [7:0] t_r30_c46_7;
  wire [7:0] t_r30_c46_8;
  wire [7:0] t_r30_c46_9;
  wire [7:0] t_r30_c46_10;
  wire [7:0] t_r30_c46_11;
  wire [7:0] t_r30_c46_12;
  wire [7:0] t_r30_c47_0;
  wire [7:0] t_r30_c47_1;
  wire [7:0] t_r30_c47_2;
  wire [7:0] t_r30_c47_3;
  wire [7:0] t_r30_c47_4;
  wire [7:0] t_r30_c47_5;
  wire [7:0] t_r30_c47_6;
  wire [7:0] t_r30_c47_7;
  wire [7:0] t_r30_c47_8;
  wire [7:0] t_r30_c47_9;
  wire [7:0] t_r30_c47_10;
  wire [7:0] t_r30_c47_11;
  wire [7:0] t_r30_c47_12;
  wire [7:0] t_r30_c48_0;
  wire [7:0] t_r30_c48_1;
  wire [7:0] t_r30_c48_2;
  wire [7:0] t_r30_c48_3;
  wire [7:0] t_r30_c48_4;
  wire [7:0] t_r30_c48_5;
  wire [7:0] t_r30_c48_6;
  wire [7:0] t_r30_c48_7;
  wire [7:0] t_r30_c48_8;
  wire [7:0] t_r30_c48_9;
  wire [7:0] t_r30_c48_10;
  wire [7:0] t_r30_c48_11;
  wire [7:0] t_r30_c48_12;
  wire [7:0] t_r30_c49_0;
  wire [7:0] t_r30_c49_1;
  wire [7:0] t_r30_c49_2;
  wire [7:0] t_r30_c49_3;
  wire [7:0] t_r30_c49_4;
  wire [7:0] t_r30_c49_5;
  wire [7:0] t_r30_c49_6;
  wire [7:0] t_r30_c49_7;
  wire [7:0] t_r30_c49_8;
  wire [7:0] t_r30_c49_9;
  wire [7:0] t_r30_c49_10;
  wire [7:0] t_r30_c49_11;
  wire [7:0] t_r30_c49_12;
  wire [7:0] t_r30_c50_0;
  wire [7:0] t_r30_c50_1;
  wire [7:0] t_r30_c50_2;
  wire [7:0] t_r30_c50_3;
  wire [7:0] t_r30_c50_4;
  wire [7:0] t_r30_c50_5;
  wire [7:0] t_r30_c50_6;
  wire [7:0] t_r30_c50_7;
  wire [7:0] t_r30_c50_8;
  wire [7:0] t_r30_c50_9;
  wire [7:0] t_r30_c50_10;
  wire [7:0] t_r30_c50_11;
  wire [7:0] t_r30_c50_12;
  wire [7:0] t_r30_c51_0;
  wire [7:0] t_r30_c51_1;
  wire [7:0] t_r30_c51_2;
  wire [7:0] t_r30_c51_3;
  wire [7:0] t_r30_c51_4;
  wire [7:0] t_r30_c51_5;
  wire [7:0] t_r30_c51_6;
  wire [7:0] t_r30_c51_7;
  wire [7:0] t_r30_c51_8;
  wire [7:0] t_r30_c51_9;
  wire [7:0] t_r30_c51_10;
  wire [7:0] t_r30_c51_11;
  wire [7:0] t_r30_c51_12;
  wire [7:0] t_r30_c52_0;
  wire [7:0] t_r30_c52_1;
  wire [7:0] t_r30_c52_2;
  wire [7:0] t_r30_c52_3;
  wire [7:0] t_r30_c52_4;
  wire [7:0] t_r30_c52_5;
  wire [7:0] t_r30_c52_6;
  wire [7:0] t_r30_c52_7;
  wire [7:0] t_r30_c52_8;
  wire [7:0] t_r30_c52_9;
  wire [7:0] t_r30_c52_10;
  wire [7:0] t_r30_c52_11;
  wire [7:0] t_r30_c52_12;
  wire [7:0] t_r30_c53_0;
  wire [7:0] t_r30_c53_1;
  wire [7:0] t_r30_c53_2;
  wire [7:0] t_r30_c53_3;
  wire [7:0] t_r30_c53_4;
  wire [7:0] t_r30_c53_5;
  wire [7:0] t_r30_c53_6;
  wire [7:0] t_r30_c53_7;
  wire [7:0] t_r30_c53_8;
  wire [7:0] t_r30_c53_9;
  wire [7:0] t_r30_c53_10;
  wire [7:0] t_r30_c53_11;
  wire [7:0] t_r30_c53_12;
  wire [7:0] t_r30_c54_0;
  wire [7:0] t_r30_c54_1;
  wire [7:0] t_r30_c54_2;
  wire [7:0] t_r30_c54_3;
  wire [7:0] t_r30_c54_4;
  wire [7:0] t_r30_c54_5;
  wire [7:0] t_r30_c54_6;
  wire [7:0] t_r30_c54_7;
  wire [7:0] t_r30_c54_8;
  wire [7:0] t_r30_c54_9;
  wire [7:0] t_r30_c54_10;
  wire [7:0] t_r30_c54_11;
  wire [7:0] t_r30_c54_12;
  wire [7:0] t_r30_c55_0;
  wire [7:0] t_r30_c55_1;
  wire [7:0] t_r30_c55_2;
  wire [7:0] t_r30_c55_3;
  wire [7:0] t_r30_c55_4;
  wire [7:0] t_r30_c55_5;
  wire [7:0] t_r30_c55_6;
  wire [7:0] t_r30_c55_7;
  wire [7:0] t_r30_c55_8;
  wire [7:0] t_r30_c55_9;
  wire [7:0] t_r30_c55_10;
  wire [7:0] t_r30_c55_11;
  wire [7:0] t_r30_c55_12;
  wire [7:0] t_r30_c56_0;
  wire [7:0] t_r30_c56_1;
  wire [7:0] t_r30_c56_2;
  wire [7:0] t_r30_c56_3;
  wire [7:0] t_r30_c56_4;
  wire [7:0] t_r30_c56_5;
  wire [7:0] t_r30_c56_6;
  wire [7:0] t_r30_c56_7;
  wire [7:0] t_r30_c56_8;
  wire [7:0] t_r30_c56_9;
  wire [7:0] t_r30_c56_10;
  wire [7:0] t_r30_c56_11;
  wire [7:0] t_r30_c56_12;
  wire [7:0] t_r30_c57_0;
  wire [7:0] t_r30_c57_1;
  wire [7:0] t_r30_c57_2;
  wire [7:0] t_r30_c57_3;
  wire [7:0] t_r30_c57_4;
  wire [7:0] t_r30_c57_5;
  wire [7:0] t_r30_c57_6;
  wire [7:0] t_r30_c57_7;
  wire [7:0] t_r30_c57_8;
  wire [7:0] t_r30_c57_9;
  wire [7:0] t_r30_c57_10;
  wire [7:0] t_r30_c57_11;
  wire [7:0] t_r30_c57_12;
  wire [7:0] t_r30_c58_0;
  wire [7:0] t_r30_c58_1;
  wire [7:0] t_r30_c58_2;
  wire [7:0] t_r30_c58_3;
  wire [7:0] t_r30_c58_4;
  wire [7:0] t_r30_c58_5;
  wire [7:0] t_r30_c58_6;
  wire [7:0] t_r30_c58_7;
  wire [7:0] t_r30_c58_8;
  wire [7:0] t_r30_c58_9;
  wire [7:0] t_r30_c58_10;
  wire [7:0] t_r30_c58_11;
  wire [7:0] t_r30_c58_12;
  wire [7:0] t_r30_c59_0;
  wire [7:0] t_r30_c59_1;
  wire [7:0] t_r30_c59_2;
  wire [7:0] t_r30_c59_3;
  wire [7:0] t_r30_c59_4;
  wire [7:0] t_r30_c59_5;
  wire [7:0] t_r30_c59_6;
  wire [7:0] t_r30_c59_7;
  wire [7:0] t_r30_c59_8;
  wire [7:0] t_r30_c59_9;
  wire [7:0] t_r30_c59_10;
  wire [7:0] t_r30_c59_11;
  wire [7:0] t_r30_c59_12;
  wire [7:0] t_r30_c60_0;
  wire [7:0] t_r30_c60_1;
  wire [7:0] t_r30_c60_2;
  wire [7:0] t_r30_c60_3;
  wire [7:0] t_r30_c60_4;
  wire [7:0] t_r30_c60_5;
  wire [7:0] t_r30_c60_6;
  wire [7:0] t_r30_c60_7;
  wire [7:0] t_r30_c60_8;
  wire [7:0] t_r30_c60_9;
  wire [7:0] t_r30_c60_10;
  wire [7:0] t_r30_c60_11;
  wire [7:0] t_r30_c60_12;
  wire [7:0] t_r30_c61_0;
  wire [7:0] t_r30_c61_1;
  wire [7:0] t_r30_c61_2;
  wire [7:0] t_r30_c61_3;
  wire [7:0] t_r30_c61_4;
  wire [7:0] t_r30_c61_5;
  wire [7:0] t_r30_c61_6;
  wire [7:0] t_r30_c61_7;
  wire [7:0] t_r30_c61_8;
  wire [7:0] t_r30_c61_9;
  wire [7:0] t_r30_c61_10;
  wire [7:0] t_r30_c61_11;
  wire [7:0] t_r30_c61_12;
  wire [7:0] t_r30_c62_0;
  wire [7:0] t_r30_c62_1;
  wire [7:0] t_r30_c62_2;
  wire [7:0] t_r30_c62_3;
  wire [7:0] t_r30_c62_4;
  wire [7:0] t_r30_c62_5;
  wire [7:0] t_r30_c62_6;
  wire [7:0] t_r30_c62_7;
  wire [7:0] t_r30_c62_8;
  wire [7:0] t_r30_c62_9;
  wire [7:0] t_r30_c62_10;
  wire [7:0] t_r30_c62_11;
  wire [7:0] t_r30_c62_12;
  wire [7:0] t_r30_c63_0;
  wire [7:0] t_r30_c63_1;
  wire [7:0] t_r30_c63_2;
  wire [7:0] t_r30_c63_3;
  wire [7:0] t_r30_c63_4;
  wire [7:0] t_r30_c63_5;
  wire [7:0] t_r30_c63_6;
  wire [7:0] t_r30_c63_7;
  wire [7:0] t_r30_c63_8;
  wire [7:0] t_r30_c63_9;
  wire [7:0] t_r30_c63_10;
  wire [7:0] t_r30_c63_11;
  wire [7:0] t_r30_c63_12;
  wire [7:0] t_r30_c64_0;
  wire [7:0] t_r30_c64_1;
  wire [7:0] t_r30_c64_2;
  wire [7:0] t_r30_c64_3;
  wire [7:0] t_r30_c64_4;
  wire [7:0] t_r30_c64_5;
  wire [7:0] t_r30_c64_6;
  wire [7:0] t_r30_c64_7;
  wire [7:0] t_r30_c64_8;
  wire [7:0] t_r30_c64_9;
  wire [7:0] t_r30_c64_10;
  wire [7:0] t_r30_c64_11;
  wire [7:0] t_r30_c64_12;
  wire [7:0] t_r30_c65_0;
  wire [7:0] t_r30_c65_1;
  wire [7:0] t_r30_c65_2;
  wire [7:0] t_r30_c65_3;
  wire [7:0] t_r30_c65_4;
  wire [7:0] t_r30_c65_5;
  wire [7:0] t_r30_c65_6;
  wire [7:0] t_r30_c65_7;
  wire [7:0] t_r30_c65_8;
  wire [7:0] t_r30_c65_9;
  wire [7:0] t_r30_c65_10;
  wire [7:0] t_r30_c65_11;
  wire [7:0] t_r30_c65_12;
  wire [7:0] t_r31_c0_0;
  wire [7:0] t_r31_c0_1;
  wire [7:0] t_r31_c0_2;
  wire [7:0] t_r31_c0_3;
  wire [7:0] t_r31_c0_4;
  wire [7:0] t_r31_c0_5;
  wire [7:0] t_r31_c0_6;
  wire [7:0] t_r31_c0_7;
  wire [7:0] t_r31_c0_8;
  wire [7:0] t_r31_c0_9;
  wire [7:0] t_r31_c0_10;
  wire [7:0] t_r31_c0_11;
  wire [7:0] t_r31_c0_12;
  wire [7:0] t_r31_c1_0;
  wire [7:0] t_r31_c1_1;
  wire [7:0] t_r31_c1_2;
  wire [7:0] t_r31_c1_3;
  wire [7:0] t_r31_c1_4;
  wire [7:0] t_r31_c1_5;
  wire [7:0] t_r31_c1_6;
  wire [7:0] t_r31_c1_7;
  wire [7:0] t_r31_c1_8;
  wire [7:0] t_r31_c1_9;
  wire [7:0] t_r31_c1_10;
  wire [7:0] t_r31_c1_11;
  wire [7:0] t_r31_c1_12;
  wire [7:0] t_r31_c2_0;
  wire [7:0] t_r31_c2_1;
  wire [7:0] t_r31_c2_2;
  wire [7:0] t_r31_c2_3;
  wire [7:0] t_r31_c2_4;
  wire [7:0] t_r31_c2_5;
  wire [7:0] t_r31_c2_6;
  wire [7:0] t_r31_c2_7;
  wire [7:0] t_r31_c2_8;
  wire [7:0] t_r31_c2_9;
  wire [7:0] t_r31_c2_10;
  wire [7:0] t_r31_c2_11;
  wire [7:0] t_r31_c2_12;
  wire [7:0] t_r31_c3_0;
  wire [7:0] t_r31_c3_1;
  wire [7:0] t_r31_c3_2;
  wire [7:0] t_r31_c3_3;
  wire [7:0] t_r31_c3_4;
  wire [7:0] t_r31_c3_5;
  wire [7:0] t_r31_c3_6;
  wire [7:0] t_r31_c3_7;
  wire [7:0] t_r31_c3_8;
  wire [7:0] t_r31_c3_9;
  wire [7:0] t_r31_c3_10;
  wire [7:0] t_r31_c3_11;
  wire [7:0] t_r31_c3_12;
  wire [7:0] t_r31_c4_0;
  wire [7:0] t_r31_c4_1;
  wire [7:0] t_r31_c4_2;
  wire [7:0] t_r31_c4_3;
  wire [7:0] t_r31_c4_4;
  wire [7:0] t_r31_c4_5;
  wire [7:0] t_r31_c4_6;
  wire [7:0] t_r31_c4_7;
  wire [7:0] t_r31_c4_8;
  wire [7:0] t_r31_c4_9;
  wire [7:0] t_r31_c4_10;
  wire [7:0] t_r31_c4_11;
  wire [7:0] t_r31_c4_12;
  wire [7:0] t_r31_c5_0;
  wire [7:0] t_r31_c5_1;
  wire [7:0] t_r31_c5_2;
  wire [7:0] t_r31_c5_3;
  wire [7:0] t_r31_c5_4;
  wire [7:0] t_r31_c5_5;
  wire [7:0] t_r31_c5_6;
  wire [7:0] t_r31_c5_7;
  wire [7:0] t_r31_c5_8;
  wire [7:0] t_r31_c5_9;
  wire [7:0] t_r31_c5_10;
  wire [7:0] t_r31_c5_11;
  wire [7:0] t_r31_c5_12;
  wire [7:0] t_r31_c6_0;
  wire [7:0] t_r31_c6_1;
  wire [7:0] t_r31_c6_2;
  wire [7:0] t_r31_c6_3;
  wire [7:0] t_r31_c6_4;
  wire [7:0] t_r31_c6_5;
  wire [7:0] t_r31_c6_6;
  wire [7:0] t_r31_c6_7;
  wire [7:0] t_r31_c6_8;
  wire [7:0] t_r31_c6_9;
  wire [7:0] t_r31_c6_10;
  wire [7:0] t_r31_c6_11;
  wire [7:0] t_r31_c6_12;
  wire [7:0] t_r31_c7_0;
  wire [7:0] t_r31_c7_1;
  wire [7:0] t_r31_c7_2;
  wire [7:0] t_r31_c7_3;
  wire [7:0] t_r31_c7_4;
  wire [7:0] t_r31_c7_5;
  wire [7:0] t_r31_c7_6;
  wire [7:0] t_r31_c7_7;
  wire [7:0] t_r31_c7_8;
  wire [7:0] t_r31_c7_9;
  wire [7:0] t_r31_c7_10;
  wire [7:0] t_r31_c7_11;
  wire [7:0] t_r31_c7_12;
  wire [7:0] t_r31_c8_0;
  wire [7:0] t_r31_c8_1;
  wire [7:0] t_r31_c8_2;
  wire [7:0] t_r31_c8_3;
  wire [7:0] t_r31_c8_4;
  wire [7:0] t_r31_c8_5;
  wire [7:0] t_r31_c8_6;
  wire [7:0] t_r31_c8_7;
  wire [7:0] t_r31_c8_8;
  wire [7:0] t_r31_c8_9;
  wire [7:0] t_r31_c8_10;
  wire [7:0] t_r31_c8_11;
  wire [7:0] t_r31_c8_12;
  wire [7:0] t_r31_c9_0;
  wire [7:0] t_r31_c9_1;
  wire [7:0] t_r31_c9_2;
  wire [7:0] t_r31_c9_3;
  wire [7:0] t_r31_c9_4;
  wire [7:0] t_r31_c9_5;
  wire [7:0] t_r31_c9_6;
  wire [7:0] t_r31_c9_7;
  wire [7:0] t_r31_c9_8;
  wire [7:0] t_r31_c9_9;
  wire [7:0] t_r31_c9_10;
  wire [7:0] t_r31_c9_11;
  wire [7:0] t_r31_c9_12;
  wire [7:0] t_r31_c10_0;
  wire [7:0] t_r31_c10_1;
  wire [7:0] t_r31_c10_2;
  wire [7:0] t_r31_c10_3;
  wire [7:0] t_r31_c10_4;
  wire [7:0] t_r31_c10_5;
  wire [7:0] t_r31_c10_6;
  wire [7:0] t_r31_c10_7;
  wire [7:0] t_r31_c10_8;
  wire [7:0] t_r31_c10_9;
  wire [7:0] t_r31_c10_10;
  wire [7:0] t_r31_c10_11;
  wire [7:0] t_r31_c10_12;
  wire [7:0] t_r31_c11_0;
  wire [7:0] t_r31_c11_1;
  wire [7:0] t_r31_c11_2;
  wire [7:0] t_r31_c11_3;
  wire [7:0] t_r31_c11_4;
  wire [7:0] t_r31_c11_5;
  wire [7:0] t_r31_c11_6;
  wire [7:0] t_r31_c11_7;
  wire [7:0] t_r31_c11_8;
  wire [7:0] t_r31_c11_9;
  wire [7:0] t_r31_c11_10;
  wire [7:0] t_r31_c11_11;
  wire [7:0] t_r31_c11_12;
  wire [7:0] t_r31_c12_0;
  wire [7:0] t_r31_c12_1;
  wire [7:0] t_r31_c12_2;
  wire [7:0] t_r31_c12_3;
  wire [7:0] t_r31_c12_4;
  wire [7:0] t_r31_c12_5;
  wire [7:0] t_r31_c12_6;
  wire [7:0] t_r31_c12_7;
  wire [7:0] t_r31_c12_8;
  wire [7:0] t_r31_c12_9;
  wire [7:0] t_r31_c12_10;
  wire [7:0] t_r31_c12_11;
  wire [7:0] t_r31_c12_12;
  wire [7:0] t_r31_c13_0;
  wire [7:0] t_r31_c13_1;
  wire [7:0] t_r31_c13_2;
  wire [7:0] t_r31_c13_3;
  wire [7:0] t_r31_c13_4;
  wire [7:0] t_r31_c13_5;
  wire [7:0] t_r31_c13_6;
  wire [7:0] t_r31_c13_7;
  wire [7:0] t_r31_c13_8;
  wire [7:0] t_r31_c13_9;
  wire [7:0] t_r31_c13_10;
  wire [7:0] t_r31_c13_11;
  wire [7:0] t_r31_c13_12;
  wire [7:0] t_r31_c14_0;
  wire [7:0] t_r31_c14_1;
  wire [7:0] t_r31_c14_2;
  wire [7:0] t_r31_c14_3;
  wire [7:0] t_r31_c14_4;
  wire [7:0] t_r31_c14_5;
  wire [7:0] t_r31_c14_6;
  wire [7:0] t_r31_c14_7;
  wire [7:0] t_r31_c14_8;
  wire [7:0] t_r31_c14_9;
  wire [7:0] t_r31_c14_10;
  wire [7:0] t_r31_c14_11;
  wire [7:0] t_r31_c14_12;
  wire [7:0] t_r31_c15_0;
  wire [7:0] t_r31_c15_1;
  wire [7:0] t_r31_c15_2;
  wire [7:0] t_r31_c15_3;
  wire [7:0] t_r31_c15_4;
  wire [7:0] t_r31_c15_5;
  wire [7:0] t_r31_c15_6;
  wire [7:0] t_r31_c15_7;
  wire [7:0] t_r31_c15_8;
  wire [7:0] t_r31_c15_9;
  wire [7:0] t_r31_c15_10;
  wire [7:0] t_r31_c15_11;
  wire [7:0] t_r31_c15_12;
  wire [7:0] t_r31_c16_0;
  wire [7:0] t_r31_c16_1;
  wire [7:0] t_r31_c16_2;
  wire [7:0] t_r31_c16_3;
  wire [7:0] t_r31_c16_4;
  wire [7:0] t_r31_c16_5;
  wire [7:0] t_r31_c16_6;
  wire [7:0] t_r31_c16_7;
  wire [7:0] t_r31_c16_8;
  wire [7:0] t_r31_c16_9;
  wire [7:0] t_r31_c16_10;
  wire [7:0] t_r31_c16_11;
  wire [7:0] t_r31_c16_12;
  wire [7:0] t_r31_c17_0;
  wire [7:0] t_r31_c17_1;
  wire [7:0] t_r31_c17_2;
  wire [7:0] t_r31_c17_3;
  wire [7:0] t_r31_c17_4;
  wire [7:0] t_r31_c17_5;
  wire [7:0] t_r31_c17_6;
  wire [7:0] t_r31_c17_7;
  wire [7:0] t_r31_c17_8;
  wire [7:0] t_r31_c17_9;
  wire [7:0] t_r31_c17_10;
  wire [7:0] t_r31_c17_11;
  wire [7:0] t_r31_c17_12;
  wire [7:0] t_r31_c18_0;
  wire [7:0] t_r31_c18_1;
  wire [7:0] t_r31_c18_2;
  wire [7:0] t_r31_c18_3;
  wire [7:0] t_r31_c18_4;
  wire [7:0] t_r31_c18_5;
  wire [7:0] t_r31_c18_6;
  wire [7:0] t_r31_c18_7;
  wire [7:0] t_r31_c18_8;
  wire [7:0] t_r31_c18_9;
  wire [7:0] t_r31_c18_10;
  wire [7:0] t_r31_c18_11;
  wire [7:0] t_r31_c18_12;
  wire [7:0] t_r31_c19_0;
  wire [7:0] t_r31_c19_1;
  wire [7:0] t_r31_c19_2;
  wire [7:0] t_r31_c19_3;
  wire [7:0] t_r31_c19_4;
  wire [7:0] t_r31_c19_5;
  wire [7:0] t_r31_c19_6;
  wire [7:0] t_r31_c19_7;
  wire [7:0] t_r31_c19_8;
  wire [7:0] t_r31_c19_9;
  wire [7:0] t_r31_c19_10;
  wire [7:0] t_r31_c19_11;
  wire [7:0] t_r31_c19_12;
  wire [7:0] t_r31_c20_0;
  wire [7:0] t_r31_c20_1;
  wire [7:0] t_r31_c20_2;
  wire [7:0] t_r31_c20_3;
  wire [7:0] t_r31_c20_4;
  wire [7:0] t_r31_c20_5;
  wire [7:0] t_r31_c20_6;
  wire [7:0] t_r31_c20_7;
  wire [7:0] t_r31_c20_8;
  wire [7:0] t_r31_c20_9;
  wire [7:0] t_r31_c20_10;
  wire [7:0] t_r31_c20_11;
  wire [7:0] t_r31_c20_12;
  wire [7:0] t_r31_c21_0;
  wire [7:0] t_r31_c21_1;
  wire [7:0] t_r31_c21_2;
  wire [7:0] t_r31_c21_3;
  wire [7:0] t_r31_c21_4;
  wire [7:0] t_r31_c21_5;
  wire [7:0] t_r31_c21_6;
  wire [7:0] t_r31_c21_7;
  wire [7:0] t_r31_c21_8;
  wire [7:0] t_r31_c21_9;
  wire [7:0] t_r31_c21_10;
  wire [7:0] t_r31_c21_11;
  wire [7:0] t_r31_c21_12;
  wire [7:0] t_r31_c22_0;
  wire [7:0] t_r31_c22_1;
  wire [7:0] t_r31_c22_2;
  wire [7:0] t_r31_c22_3;
  wire [7:0] t_r31_c22_4;
  wire [7:0] t_r31_c22_5;
  wire [7:0] t_r31_c22_6;
  wire [7:0] t_r31_c22_7;
  wire [7:0] t_r31_c22_8;
  wire [7:0] t_r31_c22_9;
  wire [7:0] t_r31_c22_10;
  wire [7:0] t_r31_c22_11;
  wire [7:0] t_r31_c22_12;
  wire [7:0] t_r31_c23_0;
  wire [7:0] t_r31_c23_1;
  wire [7:0] t_r31_c23_2;
  wire [7:0] t_r31_c23_3;
  wire [7:0] t_r31_c23_4;
  wire [7:0] t_r31_c23_5;
  wire [7:0] t_r31_c23_6;
  wire [7:0] t_r31_c23_7;
  wire [7:0] t_r31_c23_8;
  wire [7:0] t_r31_c23_9;
  wire [7:0] t_r31_c23_10;
  wire [7:0] t_r31_c23_11;
  wire [7:0] t_r31_c23_12;
  wire [7:0] t_r31_c24_0;
  wire [7:0] t_r31_c24_1;
  wire [7:0] t_r31_c24_2;
  wire [7:0] t_r31_c24_3;
  wire [7:0] t_r31_c24_4;
  wire [7:0] t_r31_c24_5;
  wire [7:0] t_r31_c24_6;
  wire [7:0] t_r31_c24_7;
  wire [7:0] t_r31_c24_8;
  wire [7:0] t_r31_c24_9;
  wire [7:0] t_r31_c24_10;
  wire [7:0] t_r31_c24_11;
  wire [7:0] t_r31_c24_12;
  wire [7:0] t_r31_c25_0;
  wire [7:0] t_r31_c25_1;
  wire [7:0] t_r31_c25_2;
  wire [7:0] t_r31_c25_3;
  wire [7:0] t_r31_c25_4;
  wire [7:0] t_r31_c25_5;
  wire [7:0] t_r31_c25_6;
  wire [7:0] t_r31_c25_7;
  wire [7:0] t_r31_c25_8;
  wire [7:0] t_r31_c25_9;
  wire [7:0] t_r31_c25_10;
  wire [7:0] t_r31_c25_11;
  wire [7:0] t_r31_c25_12;
  wire [7:0] t_r31_c26_0;
  wire [7:0] t_r31_c26_1;
  wire [7:0] t_r31_c26_2;
  wire [7:0] t_r31_c26_3;
  wire [7:0] t_r31_c26_4;
  wire [7:0] t_r31_c26_5;
  wire [7:0] t_r31_c26_6;
  wire [7:0] t_r31_c26_7;
  wire [7:0] t_r31_c26_8;
  wire [7:0] t_r31_c26_9;
  wire [7:0] t_r31_c26_10;
  wire [7:0] t_r31_c26_11;
  wire [7:0] t_r31_c26_12;
  wire [7:0] t_r31_c27_0;
  wire [7:0] t_r31_c27_1;
  wire [7:0] t_r31_c27_2;
  wire [7:0] t_r31_c27_3;
  wire [7:0] t_r31_c27_4;
  wire [7:0] t_r31_c27_5;
  wire [7:0] t_r31_c27_6;
  wire [7:0] t_r31_c27_7;
  wire [7:0] t_r31_c27_8;
  wire [7:0] t_r31_c27_9;
  wire [7:0] t_r31_c27_10;
  wire [7:0] t_r31_c27_11;
  wire [7:0] t_r31_c27_12;
  wire [7:0] t_r31_c28_0;
  wire [7:0] t_r31_c28_1;
  wire [7:0] t_r31_c28_2;
  wire [7:0] t_r31_c28_3;
  wire [7:0] t_r31_c28_4;
  wire [7:0] t_r31_c28_5;
  wire [7:0] t_r31_c28_6;
  wire [7:0] t_r31_c28_7;
  wire [7:0] t_r31_c28_8;
  wire [7:0] t_r31_c28_9;
  wire [7:0] t_r31_c28_10;
  wire [7:0] t_r31_c28_11;
  wire [7:0] t_r31_c28_12;
  wire [7:0] t_r31_c29_0;
  wire [7:0] t_r31_c29_1;
  wire [7:0] t_r31_c29_2;
  wire [7:0] t_r31_c29_3;
  wire [7:0] t_r31_c29_4;
  wire [7:0] t_r31_c29_5;
  wire [7:0] t_r31_c29_6;
  wire [7:0] t_r31_c29_7;
  wire [7:0] t_r31_c29_8;
  wire [7:0] t_r31_c29_9;
  wire [7:0] t_r31_c29_10;
  wire [7:0] t_r31_c29_11;
  wire [7:0] t_r31_c29_12;
  wire [7:0] t_r31_c30_0;
  wire [7:0] t_r31_c30_1;
  wire [7:0] t_r31_c30_2;
  wire [7:0] t_r31_c30_3;
  wire [7:0] t_r31_c30_4;
  wire [7:0] t_r31_c30_5;
  wire [7:0] t_r31_c30_6;
  wire [7:0] t_r31_c30_7;
  wire [7:0] t_r31_c30_8;
  wire [7:0] t_r31_c30_9;
  wire [7:0] t_r31_c30_10;
  wire [7:0] t_r31_c30_11;
  wire [7:0] t_r31_c30_12;
  wire [7:0] t_r31_c31_0;
  wire [7:0] t_r31_c31_1;
  wire [7:0] t_r31_c31_2;
  wire [7:0] t_r31_c31_3;
  wire [7:0] t_r31_c31_4;
  wire [7:0] t_r31_c31_5;
  wire [7:0] t_r31_c31_6;
  wire [7:0] t_r31_c31_7;
  wire [7:0] t_r31_c31_8;
  wire [7:0] t_r31_c31_9;
  wire [7:0] t_r31_c31_10;
  wire [7:0] t_r31_c31_11;
  wire [7:0] t_r31_c31_12;
  wire [7:0] t_r31_c32_0;
  wire [7:0] t_r31_c32_1;
  wire [7:0] t_r31_c32_2;
  wire [7:0] t_r31_c32_3;
  wire [7:0] t_r31_c32_4;
  wire [7:0] t_r31_c32_5;
  wire [7:0] t_r31_c32_6;
  wire [7:0] t_r31_c32_7;
  wire [7:0] t_r31_c32_8;
  wire [7:0] t_r31_c32_9;
  wire [7:0] t_r31_c32_10;
  wire [7:0] t_r31_c32_11;
  wire [7:0] t_r31_c32_12;
  wire [7:0] t_r31_c33_0;
  wire [7:0] t_r31_c33_1;
  wire [7:0] t_r31_c33_2;
  wire [7:0] t_r31_c33_3;
  wire [7:0] t_r31_c33_4;
  wire [7:0] t_r31_c33_5;
  wire [7:0] t_r31_c33_6;
  wire [7:0] t_r31_c33_7;
  wire [7:0] t_r31_c33_8;
  wire [7:0] t_r31_c33_9;
  wire [7:0] t_r31_c33_10;
  wire [7:0] t_r31_c33_11;
  wire [7:0] t_r31_c33_12;
  wire [7:0] t_r31_c34_0;
  wire [7:0] t_r31_c34_1;
  wire [7:0] t_r31_c34_2;
  wire [7:0] t_r31_c34_3;
  wire [7:0] t_r31_c34_4;
  wire [7:0] t_r31_c34_5;
  wire [7:0] t_r31_c34_6;
  wire [7:0] t_r31_c34_7;
  wire [7:0] t_r31_c34_8;
  wire [7:0] t_r31_c34_9;
  wire [7:0] t_r31_c34_10;
  wire [7:0] t_r31_c34_11;
  wire [7:0] t_r31_c34_12;
  wire [7:0] t_r31_c35_0;
  wire [7:0] t_r31_c35_1;
  wire [7:0] t_r31_c35_2;
  wire [7:0] t_r31_c35_3;
  wire [7:0] t_r31_c35_4;
  wire [7:0] t_r31_c35_5;
  wire [7:0] t_r31_c35_6;
  wire [7:0] t_r31_c35_7;
  wire [7:0] t_r31_c35_8;
  wire [7:0] t_r31_c35_9;
  wire [7:0] t_r31_c35_10;
  wire [7:0] t_r31_c35_11;
  wire [7:0] t_r31_c35_12;
  wire [7:0] t_r31_c36_0;
  wire [7:0] t_r31_c36_1;
  wire [7:0] t_r31_c36_2;
  wire [7:0] t_r31_c36_3;
  wire [7:0] t_r31_c36_4;
  wire [7:0] t_r31_c36_5;
  wire [7:0] t_r31_c36_6;
  wire [7:0] t_r31_c36_7;
  wire [7:0] t_r31_c36_8;
  wire [7:0] t_r31_c36_9;
  wire [7:0] t_r31_c36_10;
  wire [7:0] t_r31_c36_11;
  wire [7:0] t_r31_c36_12;
  wire [7:0] t_r31_c37_0;
  wire [7:0] t_r31_c37_1;
  wire [7:0] t_r31_c37_2;
  wire [7:0] t_r31_c37_3;
  wire [7:0] t_r31_c37_4;
  wire [7:0] t_r31_c37_5;
  wire [7:0] t_r31_c37_6;
  wire [7:0] t_r31_c37_7;
  wire [7:0] t_r31_c37_8;
  wire [7:0] t_r31_c37_9;
  wire [7:0] t_r31_c37_10;
  wire [7:0] t_r31_c37_11;
  wire [7:0] t_r31_c37_12;
  wire [7:0] t_r31_c38_0;
  wire [7:0] t_r31_c38_1;
  wire [7:0] t_r31_c38_2;
  wire [7:0] t_r31_c38_3;
  wire [7:0] t_r31_c38_4;
  wire [7:0] t_r31_c38_5;
  wire [7:0] t_r31_c38_6;
  wire [7:0] t_r31_c38_7;
  wire [7:0] t_r31_c38_8;
  wire [7:0] t_r31_c38_9;
  wire [7:0] t_r31_c38_10;
  wire [7:0] t_r31_c38_11;
  wire [7:0] t_r31_c38_12;
  wire [7:0] t_r31_c39_0;
  wire [7:0] t_r31_c39_1;
  wire [7:0] t_r31_c39_2;
  wire [7:0] t_r31_c39_3;
  wire [7:0] t_r31_c39_4;
  wire [7:0] t_r31_c39_5;
  wire [7:0] t_r31_c39_6;
  wire [7:0] t_r31_c39_7;
  wire [7:0] t_r31_c39_8;
  wire [7:0] t_r31_c39_9;
  wire [7:0] t_r31_c39_10;
  wire [7:0] t_r31_c39_11;
  wire [7:0] t_r31_c39_12;
  wire [7:0] t_r31_c40_0;
  wire [7:0] t_r31_c40_1;
  wire [7:0] t_r31_c40_2;
  wire [7:0] t_r31_c40_3;
  wire [7:0] t_r31_c40_4;
  wire [7:0] t_r31_c40_5;
  wire [7:0] t_r31_c40_6;
  wire [7:0] t_r31_c40_7;
  wire [7:0] t_r31_c40_8;
  wire [7:0] t_r31_c40_9;
  wire [7:0] t_r31_c40_10;
  wire [7:0] t_r31_c40_11;
  wire [7:0] t_r31_c40_12;
  wire [7:0] t_r31_c41_0;
  wire [7:0] t_r31_c41_1;
  wire [7:0] t_r31_c41_2;
  wire [7:0] t_r31_c41_3;
  wire [7:0] t_r31_c41_4;
  wire [7:0] t_r31_c41_5;
  wire [7:0] t_r31_c41_6;
  wire [7:0] t_r31_c41_7;
  wire [7:0] t_r31_c41_8;
  wire [7:0] t_r31_c41_9;
  wire [7:0] t_r31_c41_10;
  wire [7:0] t_r31_c41_11;
  wire [7:0] t_r31_c41_12;
  wire [7:0] t_r31_c42_0;
  wire [7:0] t_r31_c42_1;
  wire [7:0] t_r31_c42_2;
  wire [7:0] t_r31_c42_3;
  wire [7:0] t_r31_c42_4;
  wire [7:0] t_r31_c42_5;
  wire [7:0] t_r31_c42_6;
  wire [7:0] t_r31_c42_7;
  wire [7:0] t_r31_c42_8;
  wire [7:0] t_r31_c42_9;
  wire [7:0] t_r31_c42_10;
  wire [7:0] t_r31_c42_11;
  wire [7:0] t_r31_c42_12;
  wire [7:0] t_r31_c43_0;
  wire [7:0] t_r31_c43_1;
  wire [7:0] t_r31_c43_2;
  wire [7:0] t_r31_c43_3;
  wire [7:0] t_r31_c43_4;
  wire [7:0] t_r31_c43_5;
  wire [7:0] t_r31_c43_6;
  wire [7:0] t_r31_c43_7;
  wire [7:0] t_r31_c43_8;
  wire [7:0] t_r31_c43_9;
  wire [7:0] t_r31_c43_10;
  wire [7:0] t_r31_c43_11;
  wire [7:0] t_r31_c43_12;
  wire [7:0] t_r31_c44_0;
  wire [7:0] t_r31_c44_1;
  wire [7:0] t_r31_c44_2;
  wire [7:0] t_r31_c44_3;
  wire [7:0] t_r31_c44_4;
  wire [7:0] t_r31_c44_5;
  wire [7:0] t_r31_c44_6;
  wire [7:0] t_r31_c44_7;
  wire [7:0] t_r31_c44_8;
  wire [7:0] t_r31_c44_9;
  wire [7:0] t_r31_c44_10;
  wire [7:0] t_r31_c44_11;
  wire [7:0] t_r31_c44_12;
  wire [7:0] t_r31_c45_0;
  wire [7:0] t_r31_c45_1;
  wire [7:0] t_r31_c45_2;
  wire [7:0] t_r31_c45_3;
  wire [7:0] t_r31_c45_4;
  wire [7:0] t_r31_c45_5;
  wire [7:0] t_r31_c45_6;
  wire [7:0] t_r31_c45_7;
  wire [7:0] t_r31_c45_8;
  wire [7:0] t_r31_c45_9;
  wire [7:0] t_r31_c45_10;
  wire [7:0] t_r31_c45_11;
  wire [7:0] t_r31_c45_12;
  wire [7:0] t_r31_c46_0;
  wire [7:0] t_r31_c46_1;
  wire [7:0] t_r31_c46_2;
  wire [7:0] t_r31_c46_3;
  wire [7:0] t_r31_c46_4;
  wire [7:0] t_r31_c46_5;
  wire [7:0] t_r31_c46_6;
  wire [7:0] t_r31_c46_7;
  wire [7:0] t_r31_c46_8;
  wire [7:0] t_r31_c46_9;
  wire [7:0] t_r31_c46_10;
  wire [7:0] t_r31_c46_11;
  wire [7:0] t_r31_c46_12;
  wire [7:0] t_r31_c47_0;
  wire [7:0] t_r31_c47_1;
  wire [7:0] t_r31_c47_2;
  wire [7:0] t_r31_c47_3;
  wire [7:0] t_r31_c47_4;
  wire [7:0] t_r31_c47_5;
  wire [7:0] t_r31_c47_6;
  wire [7:0] t_r31_c47_7;
  wire [7:0] t_r31_c47_8;
  wire [7:0] t_r31_c47_9;
  wire [7:0] t_r31_c47_10;
  wire [7:0] t_r31_c47_11;
  wire [7:0] t_r31_c47_12;
  wire [7:0] t_r31_c48_0;
  wire [7:0] t_r31_c48_1;
  wire [7:0] t_r31_c48_2;
  wire [7:0] t_r31_c48_3;
  wire [7:0] t_r31_c48_4;
  wire [7:0] t_r31_c48_5;
  wire [7:0] t_r31_c48_6;
  wire [7:0] t_r31_c48_7;
  wire [7:0] t_r31_c48_8;
  wire [7:0] t_r31_c48_9;
  wire [7:0] t_r31_c48_10;
  wire [7:0] t_r31_c48_11;
  wire [7:0] t_r31_c48_12;
  wire [7:0] t_r31_c49_0;
  wire [7:0] t_r31_c49_1;
  wire [7:0] t_r31_c49_2;
  wire [7:0] t_r31_c49_3;
  wire [7:0] t_r31_c49_4;
  wire [7:0] t_r31_c49_5;
  wire [7:0] t_r31_c49_6;
  wire [7:0] t_r31_c49_7;
  wire [7:0] t_r31_c49_8;
  wire [7:0] t_r31_c49_9;
  wire [7:0] t_r31_c49_10;
  wire [7:0] t_r31_c49_11;
  wire [7:0] t_r31_c49_12;
  wire [7:0] t_r31_c50_0;
  wire [7:0] t_r31_c50_1;
  wire [7:0] t_r31_c50_2;
  wire [7:0] t_r31_c50_3;
  wire [7:0] t_r31_c50_4;
  wire [7:0] t_r31_c50_5;
  wire [7:0] t_r31_c50_6;
  wire [7:0] t_r31_c50_7;
  wire [7:0] t_r31_c50_8;
  wire [7:0] t_r31_c50_9;
  wire [7:0] t_r31_c50_10;
  wire [7:0] t_r31_c50_11;
  wire [7:0] t_r31_c50_12;
  wire [7:0] t_r31_c51_0;
  wire [7:0] t_r31_c51_1;
  wire [7:0] t_r31_c51_2;
  wire [7:0] t_r31_c51_3;
  wire [7:0] t_r31_c51_4;
  wire [7:0] t_r31_c51_5;
  wire [7:0] t_r31_c51_6;
  wire [7:0] t_r31_c51_7;
  wire [7:0] t_r31_c51_8;
  wire [7:0] t_r31_c51_9;
  wire [7:0] t_r31_c51_10;
  wire [7:0] t_r31_c51_11;
  wire [7:0] t_r31_c51_12;
  wire [7:0] t_r31_c52_0;
  wire [7:0] t_r31_c52_1;
  wire [7:0] t_r31_c52_2;
  wire [7:0] t_r31_c52_3;
  wire [7:0] t_r31_c52_4;
  wire [7:0] t_r31_c52_5;
  wire [7:0] t_r31_c52_6;
  wire [7:0] t_r31_c52_7;
  wire [7:0] t_r31_c52_8;
  wire [7:0] t_r31_c52_9;
  wire [7:0] t_r31_c52_10;
  wire [7:0] t_r31_c52_11;
  wire [7:0] t_r31_c52_12;
  wire [7:0] t_r31_c53_0;
  wire [7:0] t_r31_c53_1;
  wire [7:0] t_r31_c53_2;
  wire [7:0] t_r31_c53_3;
  wire [7:0] t_r31_c53_4;
  wire [7:0] t_r31_c53_5;
  wire [7:0] t_r31_c53_6;
  wire [7:0] t_r31_c53_7;
  wire [7:0] t_r31_c53_8;
  wire [7:0] t_r31_c53_9;
  wire [7:0] t_r31_c53_10;
  wire [7:0] t_r31_c53_11;
  wire [7:0] t_r31_c53_12;
  wire [7:0] t_r31_c54_0;
  wire [7:0] t_r31_c54_1;
  wire [7:0] t_r31_c54_2;
  wire [7:0] t_r31_c54_3;
  wire [7:0] t_r31_c54_4;
  wire [7:0] t_r31_c54_5;
  wire [7:0] t_r31_c54_6;
  wire [7:0] t_r31_c54_7;
  wire [7:0] t_r31_c54_8;
  wire [7:0] t_r31_c54_9;
  wire [7:0] t_r31_c54_10;
  wire [7:0] t_r31_c54_11;
  wire [7:0] t_r31_c54_12;
  wire [7:0] t_r31_c55_0;
  wire [7:0] t_r31_c55_1;
  wire [7:0] t_r31_c55_2;
  wire [7:0] t_r31_c55_3;
  wire [7:0] t_r31_c55_4;
  wire [7:0] t_r31_c55_5;
  wire [7:0] t_r31_c55_6;
  wire [7:0] t_r31_c55_7;
  wire [7:0] t_r31_c55_8;
  wire [7:0] t_r31_c55_9;
  wire [7:0] t_r31_c55_10;
  wire [7:0] t_r31_c55_11;
  wire [7:0] t_r31_c55_12;
  wire [7:0] t_r31_c56_0;
  wire [7:0] t_r31_c56_1;
  wire [7:0] t_r31_c56_2;
  wire [7:0] t_r31_c56_3;
  wire [7:0] t_r31_c56_4;
  wire [7:0] t_r31_c56_5;
  wire [7:0] t_r31_c56_6;
  wire [7:0] t_r31_c56_7;
  wire [7:0] t_r31_c56_8;
  wire [7:0] t_r31_c56_9;
  wire [7:0] t_r31_c56_10;
  wire [7:0] t_r31_c56_11;
  wire [7:0] t_r31_c56_12;
  wire [7:0] t_r31_c57_0;
  wire [7:0] t_r31_c57_1;
  wire [7:0] t_r31_c57_2;
  wire [7:0] t_r31_c57_3;
  wire [7:0] t_r31_c57_4;
  wire [7:0] t_r31_c57_5;
  wire [7:0] t_r31_c57_6;
  wire [7:0] t_r31_c57_7;
  wire [7:0] t_r31_c57_8;
  wire [7:0] t_r31_c57_9;
  wire [7:0] t_r31_c57_10;
  wire [7:0] t_r31_c57_11;
  wire [7:0] t_r31_c57_12;
  wire [7:0] t_r31_c58_0;
  wire [7:0] t_r31_c58_1;
  wire [7:0] t_r31_c58_2;
  wire [7:0] t_r31_c58_3;
  wire [7:0] t_r31_c58_4;
  wire [7:0] t_r31_c58_5;
  wire [7:0] t_r31_c58_6;
  wire [7:0] t_r31_c58_7;
  wire [7:0] t_r31_c58_8;
  wire [7:0] t_r31_c58_9;
  wire [7:0] t_r31_c58_10;
  wire [7:0] t_r31_c58_11;
  wire [7:0] t_r31_c58_12;
  wire [7:0] t_r31_c59_0;
  wire [7:0] t_r31_c59_1;
  wire [7:0] t_r31_c59_2;
  wire [7:0] t_r31_c59_3;
  wire [7:0] t_r31_c59_4;
  wire [7:0] t_r31_c59_5;
  wire [7:0] t_r31_c59_6;
  wire [7:0] t_r31_c59_7;
  wire [7:0] t_r31_c59_8;
  wire [7:0] t_r31_c59_9;
  wire [7:0] t_r31_c59_10;
  wire [7:0] t_r31_c59_11;
  wire [7:0] t_r31_c59_12;
  wire [7:0] t_r31_c60_0;
  wire [7:0] t_r31_c60_1;
  wire [7:0] t_r31_c60_2;
  wire [7:0] t_r31_c60_3;
  wire [7:0] t_r31_c60_4;
  wire [7:0] t_r31_c60_5;
  wire [7:0] t_r31_c60_6;
  wire [7:0] t_r31_c60_7;
  wire [7:0] t_r31_c60_8;
  wire [7:0] t_r31_c60_9;
  wire [7:0] t_r31_c60_10;
  wire [7:0] t_r31_c60_11;
  wire [7:0] t_r31_c60_12;
  wire [7:0] t_r31_c61_0;
  wire [7:0] t_r31_c61_1;
  wire [7:0] t_r31_c61_2;
  wire [7:0] t_r31_c61_3;
  wire [7:0] t_r31_c61_4;
  wire [7:0] t_r31_c61_5;
  wire [7:0] t_r31_c61_6;
  wire [7:0] t_r31_c61_7;
  wire [7:0] t_r31_c61_8;
  wire [7:0] t_r31_c61_9;
  wire [7:0] t_r31_c61_10;
  wire [7:0] t_r31_c61_11;
  wire [7:0] t_r31_c61_12;
  wire [7:0] t_r31_c62_0;
  wire [7:0] t_r31_c62_1;
  wire [7:0] t_r31_c62_2;
  wire [7:0] t_r31_c62_3;
  wire [7:0] t_r31_c62_4;
  wire [7:0] t_r31_c62_5;
  wire [7:0] t_r31_c62_6;
  wire [7:0] t_r31_c62_7;
  wire [7:0] t_r31_c62_8;
  wire [7:0] t_r31_c62_9;
  wire [7:0] t_r31_c62_10;
  wire [7:0] t_r31_c62_11;
  wire [7:0] t_r31_c62_12;
  wire [7:0] t_r31_c63_0;
  wire [7:0] t_r31_c63_1;
  wire [7:0] t_r31_c63_2;
  wire [7:0] t_r31_c63_3;
  wire [7:0] t_r31_c63_4;
  wire [7:0] t_r31_c63_5;
  wire [7:0] t_r31_c63_6;
  wire [7:0] t_r31_c63_7;
  wire [7:0] t_r31_c63_8;
  wire [7:0] t_r31_c63_9;
  wire [7:0] t_r31_c63_10;
  wire [7:0] t_r31_c63_11;
  wire [7:0] t_r31_c63_12;
  wire [7:0] t_r31_c64_0;
  wire [7:0] t_r31_c64_1;
  wire [7:0] t_r31_c64_2;
  wire [7:0] t_r31_c64_3;
  wire [7:0] t_r31_c64_4;
  wire [7:0] t_r31_c64_5;
  wire [7:0] t_r31_c64_6;
  wire [7:0] t_r31_c64_7;
  wire [7:0] t_r31_c64_8;
  wire [7:0] t_r31_c64_9;
  wire [7:0] t_r31_c64_10;
  wire [7:0] t_r31_c64_11;
  wire [7:0] t_r31_c64_12;
  wire [7:0] t_r31_c65_0;
  wire [7:0] t_r31_c65_1;
  wire [7:0] t_r31_c65_2;
  wire [7:0] t_r31_c65_3;
  wire [7:0] t_r31_c65_4;
  wire [7:0] t_r31_c65_5;
  wire [7:0] t_r31_c65_6;
  wire [7:0] t_r31_c65_7;
  wire [7:0] t_r31_c65_8;
  wire [7:0] t_r31_c65_9;
  wire [7:0] t_r31_c65_10;
  wire [7:0] t_r31_c65_11;
  wire [7:0] t_r31_c65_12;
  wire [7:0] t_r32_c0_0;
  wire [7:0] t_r32_c0_1;
  wire [7:0] t_r32_c0_2;
  wire [7:0] t_r32_c0_3;
  wire [7:0] t_r32_c0_4;
  wire [7:0] t_r32_c0_5;
  wire [7:0] t_r32_c0_6;
  wire [7:0] t_r32_c0_7;
  wire [7:0] t_r32_c0_8;
  wire [7:0] t_r32_c0_9;
  wire [7:0] t_r32_c0_10;
  wire [7:0] t_r32_c0_11;
  wire [7:0] t_r32_c0_12;
  wire [7:0] t_r32_c1_0;
  wire [7:0] t_r32_c1_1;
  wire [7:0] t_r32_c1_2;
  wire [7:0] t_r32_c1_3;
  wire [7:0] t_r32_c1_4;
  wire [7:0] t_r32_c1_5;
  wire [7:0] t_r32_c1_6;
  wire [7:0] t_r32_c1_7;
  wire [7:0] t_r32_c1_8;
  wire [7:0] t_r32_c1_9;
  wire [7:0] t_r32_c1_10;
  wire [7:0] t_r32_c1_11;
  wire [7:0] t_r32_c1_12;
  wire [7:0] t_r32_c2_0;
  wire [7:0] t_r32_c2_1;
  wire [7:0] t_r32_c2_2;
  wire [7:0] t_r32_c2_3;
  wire [7:0] t_r32_c2_4;
  wire [7:0] t_r32_c2_5;
  wire [7:0] t_r32_c2_6;
  wire [7:0] t_r32_c2_7;
  wire [7:0] t_r32_c2_8;
  wire [7:0] t_r32_c2_9;
  wire [7:0] t_r32_c2_10;
  wire [7:0] t_r32_c2_11;
  wire [7:0] t_r32_c2_12;
  wire [7:0] t_r32_c3_0;
  wire [7:0] t_r32_c3_1;
  wire [7:0] t_r32_c3_2;
  wire [7:0] t_r32_c3_3;
  wire [7:0] t_r32_c3_4;
  wire [7:0] t_r32_c3_5;
  wire [7:0] t_r32_c3_6;
  wire [7:0] t_r32_c3_7;
  wire [7:0] t_r32_c3_8;
  wire [7:0] t_r32_c3_9;
  wire [7:0] t_r32_c3_10;
  wire [7:0] t_r32_c3_11;
  wire [7:0] t_r32_c3_12;
  wire [7:0] t_r32_c4_0;
  wire [7:0] t_r32_c4_1;
  wire [7:0] t_r32_c4_2;
  wire [7:0] t_r32_c4_3;
  wire [7:0] t_r32_c4_4;
  wire [7:0] t_r32_c4_5;
  wire [7:0] t_r32_c4_6;
  wire [7:0] t_r32_c4_7;
  wire [7:0] t_r32_c4_8;
  wire [7:0] t_r32_c4_9;
  wire [7:0] t_r32_c4_10;
  wire [7:0] t_r32_c4_11;
  wire [7:0] t_r32_c4_12;
  wire [7:0] t_r32_c5_0;
  wire [7:0] t_r32_c5_1;
  wire [7:0] t_r32_c5_2;
  wire [7:0] t_r32_c5_3;
  wire [7:0] t_r32_c5_4;
  wire [7:0] t_r32_c5_5;
  wire [7:0] t_r32_c5_6;
  wire [7:0] t_r32_c5_7;
  wire [7:0] t_r32_c5_8;
  wire [7:0] t_r32_c5_9;
  wire [7:0] t_r32_c5_10;
  wire [7:0] t_r32_c5_11;
  wire [7:0] t_r32_c5_12;
  wire [7:0] t_r32_c6_0;
  wire [7:0] t_r32_c6_1;
  wire [7:0] t_r32_c6_2;
  wire [7:0] t_r32_c6_3;
  wire [7:0] t_r32_c6_4;
  wire [7:0] t_r32_c6_5;
  wire [7:0] t_r32_c6_6;
  wire [7:0] t_r32_c6_7;
  wire [7:0] t_r32_c6_8;
  wire [7:0] t_r32_c6_9;
  wire [7:0] t_r32_c6_10;
  wire [7:0] t_r32_c6_11;
  wire [7:0] t_r32_c6_12;
  wire [7:0] t_r32_c7_0;
  wire [7:0] t_r32_c7_1;
  wire [7:0] t_r32_c7_2;
  wire [7:0] t_r32_c7_3;
  wire [7:0] t_r32_c7_4;
  wire [7:0] t_r32_c7_5;
  wire [7:0] t_r32_c7_6;
  wire [7:0] t_r32_c7_7;
  wire [7:0] t_r32_c7_8;
  wire [7:0] t_r32_c7_9;
  wire [7:0] t_r32_c7_10;
  wire [7:0] t_r32_c7_11;
  wire [7:0] t_r32_c7_12;
  wire [7:0] t_r32_c8_0;
  wire [7:0] t_r32_c8_1;
  wire [7:0] t_r32_c8_2;
  wire [7:0] t_r32_c8_3;
  wire [7:0] t_r32_c8_4;
  wire [7:0] t_r32_c8_5;
  wire [7:0] t_r32_c8_6;
  wire [7:0] t_r32_c8_7;
  wire [7:0] t_r32_c8_8;
  wire [7:0] t_r32_c8_9;
  wire [7:0] t_r32_c8_10;
  wire [7:0] t_r32_c8_11;
  wire [7:0] t_r32_c8_12;
  wire [7:0] t_r32_c9_0;
  wire [7:0] t_r32_c9_1;
  wire [7:0] t_r32_c9_2;
  wire [7:0] t_r32_c9_3;
  wire [7:0] t_r32_c9_4;
  wire [7:0] t_r32_c9_5;
  wire [7:0] t_r32_c9_6;
  wire [7:0] t_r32_c9_7;
  wire [7:0] t_r32_c9_8;
  wire [7:0] t_r32_c9_9;
  wire [7:0] t_r32_c9_10;
  wire [7:0] t_r32_c9_11;
  wire [7:0] t_r32_c9_12;
  wire [7:0] t_r32_c10_0;
  wire [7:0] t_r32_c10_1;
  wire [7:0] t_r32_c10_2;
  wire [7:0] t_r32_c10_3;
  wire [7:0] t_r32_c10_4;
  wire [7:0] t_r32_c10_5;
  wire [7:0] t_r32_c10_6;
  wire [7:0] t_r32_c10_7;
  wire [7:0] t_r32_c10_8;
  wire [7:0] t_r32_c10_9;
  wire [7:0] t_r32_c10_10;
  wire [7:0] t_r32_c10_11;
  wire [7:0] t_r32_c10_12;
  wire [7:0] t_r32_c11_0;
  wire [7:0] t_r32_c11_1;
  wire [7:0] t_r32_c11_2;
  wire [7:0] t_r32_c11_3;
  wire [7:0] t_r32_c11_4;
  wire [7:0] t_r32_c11_5;
  wire [7:0] t_r32_c11_6;
  wire [7:0] t_r32_c11_7;
  wire [7:0] t_r32_c11_8;
  wire [7:0] t_r32_c11_9;
  wire [7:0] t_r32_c11_10;
  wire [7:0] t_r32_c11_11;
  wire [7:0] t_r32_c11_12;
  wire [7:0] t_r32_c12_0;
  wire [7:0] t_r32_c12_1;
  wire [7:0] t_r32_c12_2;
  wire [7:0] t_r32_c12_3;
  wire [7:0] t_r32_c12_4;
  wire [7:0] t_r32_c12_5;
  wire [7:0] t_r32_c12_6;
  wire [7:0] t_r32_c12_7;
  wire [7:0] t_r32_c12_8;
  wire [7:0] t_r32_c12_9;
  wire [7:0] t_r32_c12_10;
  wire [7:0] t_r32_c12_11;
  wire [7:0] t_r32_c12_12;
  wire [7:0] t_r32_c13_0;
  wire [7:0] t_r32_c13_1;
  wire [7:0] t_r32_c13_2;
  wire [7:0] t_r32_c13_3;
  wire [7:0] t_r32_c13_4;
  wire [7:0] t_r32_c13_5;
  wire [7:0] t_r32_c13_6;
  wire [7:0] t_r32_c13_7;
  wire [7:0] t_r32_c13_8;
  wire [7:0] t_r32_c13_9;
  wire [7:0] t_r32_c13_10;
  wire [7:0] t_r32_c13_11;
  wire [7:0] t_r32_c13_12;
  wire [7:0] t_r32_c14_0;
  wire [7:0] t_r32_c14_1;
  wire [7:0] t_r32_c14_2;
  wire [7:0] t_r32_c14_3;
  wire [7:0] t_r32_c14_4;
  wire [7:0] t_r32_c14_5;
  wire [7:0] t_r32_c14_6;
  wire [7:0] t_r32_c14_7;
  wire [7:0] t_r32_c14_8;
  wire [7:0] t_r32_c14_9;
  wire [7:0] t_r32_c14_10;
  wire [7:0] t_r32_c14_11;
  wire [7:0] t_r32_c14_12;
  wire [7:0] t_r32_c15_0;
  wire [7:0] t_r32_c15_1;
  wire [7:0] t_r32_c15_2;
  wire [7:0] t_r32_c15_3;
  wire [7:0] t_r32_c15_4;
  wire [7:0] t_r32_c15_5;
  wire [7:0] t_r32_c15_6;
  wire [7:0] t_r32_c15_7;
  wire [7:0] t_r32_c15_8;
  wire [7:0] t_r32_c15_9;
  wire [7:0] t_r32_c15_10;
  wire [7:0] t_r32_c15_11;
  wire [7:0] t_r32_c15_12;
  wire [7:0] t_r32_c16_0;
  wire [7:0] t_r32_c16_1;
  wire [7:0] t_r32_c16_2;
  wire [7:0] t_r32_c16_3;
  wire [7:0] t_r32_c16_4;
  wire [7:0] t_r32_c16_5;
  wire [7:0] t_r32_c16_6;
  wire [7:0] t_r32_c16_7;
  wire [7:0] t_r32_c16_8;
  wire [7:0] t_r32_c16_9;
  wire [7:0] t_r32_c16_10;
  wire [7:0] t_r32_c16_11;
  wire [7:0] t_r32_c16_12;
  wire [7:0] t_r32_c17_0;
  wire [7:0] t_r32_c17_1;
  wire [7:0] t_r32_c17_2;
  wire [7:0] t_r32_c17_3;
  wire [7:0] t_r32_c17_4;
  wire [7:0] t_r32_c17_5;
  wire [7:0] t_r32_c17_6;
  wire [7:0] t_r32_c17_7;
  wire [7:0] t_r32_c17_8;
  wire [7:0] t_r32_c17_9;
  wire [7:0] t_r32_c17_10;
  wire [7:0] t_r32_c17_11;
  wire [7:0] t_r32_c17_12;
  wire [7:0] t_r32_c18_0;
  wire [7:0] t_r32_c18_1;
  wire [7:0] t_r32_c18_2;
  wire [7:0] t_r32_c18_3;
  wire [7:0] t_r32_c18_4;
  wire [7:0] t_r32_c18_5;
  wire [7:0] t_r32_c18_6;
  wire [7:0] t_r32_c18_7;
  wire [7:0] t_r32_c18_8;
  wire [7:0] t_r32_c18_9;
  wire [7:0] t_r32_c18_10;
  wire [7:0] t_r32_c18_11;
  wire [7:0] t_r32_c18_12;
  wire [7:0] t_r32_c19_0;
  wire [7:0] t_r32_c19_1;
  wire [7:0] t_r32_c19_2;
  wire [7:0] t_r32_c19_3;
  wire [7:0] t_r32_c19_4;
  wire [7:0] t_r32_c19_5;
  wire [7:0] t_r32_c19_6;
  wire [7:0] t_r32_c19_7;
  wire [7:0] t_r32_c19_8;
  wire [7:0] t_r32_c19_9;
  wire [7:0] t_r32_c19_10;
  wire [7:0] t_r32_c19_11;
  wire [7:0] t_r32_c19_12;
  wire [7:0] t_r32_c20_0;
  wire [7:0] t_r32_c20_1;
  wire [7:0] t_r32_c20_2;
  wire [7:0] t_r32_c20_3;
  wire [7:0] t_r32_c20_4;
  wire [7:0] t_r32_c20_5;
  wire [7:0] t_r32_c20_6;
  wire [7:0] t_r32_c20_7;
  wire [7:0] t_r32_c20_8;
  wire [7:0] t_r32_c20_9;
  wire [7:0] t_r32_c20_10;
  wire [7:0] t_r32_c20_11;
  wire [7:0] t_r32_c20_12;
  wire [7:0] t_r32_c21_0;
  wire [7:0] t_r32_c21_1;
  wire [7:0] t_r32_c21_2;
  wire [7:0] t_r32_c21_3;
  wire [7:0] t_r32_c21_4;
  wire [7:0] t_r32_c21_5;
  wire [7:0] t_r32_c21_6;
  wire [7:0] t_r32_c21_7;
  wire [7:0] t_r32_c21_8;
  wire [7:0] t_r32_c21_9;
  wire [7:0] t_r32_c21_10;
  wire [7:0] t_r32_c21_11;
  wire [7:0] t_r32_c21_12;
  wire [7:0] t_r32_c22_0;
  wire [7:0] t_r32_c22_1;
  wire [7:0] t_r32_c22_2;
  wire [7:0] t_r32_c22_3;
  wire [7:0] t_r32_c22_4;
  wire [7:0] t_r32_c22_5;
  wire [7:0] t_r32_c22_6;
  wire [7:0] t_r32_c22_7;
  wire [7:0] t_r32_c22_8;
  wire [7:0] t_r32_c22_9;
  wire [7:0] t_r32_c22_10;
  wire [7:0] t_r32_c22_11;
  wire [7:0] t_r32_c22_12;
  wire [7:0] t_r32_c23_0;
  wire [7:0] t_r32_c23_1;
  wire [7:0] t_r32_c23_2;
  wire [7:0] t_r32_c23_3;
  wire [7:0] t_r32_c23_4;
  wire [7:0] t_r32_c23_5;
  wire [7:0] t_r32_c23_6;
  wire [7:0] t_r32_c23_7;
  wire [7:0] t_r32_c23_8;
  wire [7:0] t_r32_c23_9;
  wire [7:0] t_r32_c23_10;
  wire [7:0] t_r32_c23_11;
  wire [7:0] t_r32_c23_12;
  wire [7:0] t_r32_c24_0;
  wire [7:0] t_r32_c24_1;
  wire [7:0] t_r32_c24_2;
  wire [7:0] t_r32_c24_3;
  wire [7:0] t_r32_c24_4;
  wire [7:0] t_r32_c24_5;
  wire [7:0] t_r32_c24_6;
  wire [7:0] t_r32_c24_7;
  wire [7:0] t_r32_c24_8;
  wire [7:0] t_r32_c24_9;
  wire [7:0] t_r32_c24_10;
  wire [7:0] t_r32_c24_11;
  wire [7:0] t_r32_c24_12;
  wire [7:0] t_r32_c25_0;
  wire [7:0] t_r32_c25_1;
  wire [7:0] t_r32_c25_2;
  wire [7:0] t_r32_c25_3;
  wire [7:0] t_r32_c25_4;
  wire [7:0] t_r32_c25_5;
  wire [7:0] t_r32_c25_6;
  wire [7:0] t_r32_c25_7;
  wire [7:0] t_r32_c25_8;
  wire [7:0] t_r32_c25_9;
  wire [7:0] t_r32_c25_10;
  wire [7:0] t_r32_c25_11;
  wire [7:0] t_r32_c25_12;
  wire [7:0] t_r32_c26_0;
  wire [7:0] t_r32_c26_1;
  wire [7:0] t_r32_c26_2;
  wire [7:0] t_r32_c26_3;
  wire [7:0] t_r32_c26_4;
  wire [7:0] t_r32_c26_5;
  wire [7:0] t_r32_c26_6;
  wire [7:0] t_r32_c26_7;
  wire [7:0] t_r32_c26_8;
  wire [7:0] t_r32_c26_9;
  wire [7:0] t_r32_c26_10;
  wire [7:0] t_r32_c26_11;
  wire [7:0] t_r32_c26_12;
  wire [7:0] t_r32_c27_0;
  wire [7:0] t_r32_c27_1;
  wire [7:0] t_r32_c27_2;
  wire [7:0] t_r32_c27_3;
  wire [7:0] t_r32_c27_4;
  wire [7:0] t_r32_c27_5;
  wire [7:0] t_r32_c27_6;
  wire [7:0] t_r32_c27_7;
  wire [7:0] t_r32_c27_8;
  wire [7:0] t_r32_c27_9;
  wire [7:0] t_r32_c27_10;
  wire [7:0] t_r32_c27_11;
  wire [7:0] t_r32_c27_12;
  wire [7:0] t_r32_c28_0;
  wire [7:0] t_r32_c28_1;
  wire [7:0] t_r32_c28_2;
  wire [7:0] t_r32_c28_3;
  wire [7:0] t_r32_c28_4;
  wire [7:0] t_r32_c28_5;
  wire [7:0] t_r32_c28_6;
  wire [7:0] t_r32_c28_7;
  wire [7:0] t_r32_c28_8;
  wire [7:0] t_r32_c28_9;
  wire [7:0] t_r32_c28_10;
  wire [7:0] t_r32_c28_11;
  wire [7:0] t_r32_c28_12;
  wire [7:0] t_r32_c29_0;
  wire [7:0] t_r32_c29_1;
  wire [7:0] t_r32_c29_2;
  wire [7:0] t_r32_c29_3;
  wire [7:0] t_r32_c29_4;
  wire [7:0] t_r32_c29_5;
  wire [7:0] t_r32_c29_6;
  wire [7:0] t_r32_c29_7;
  wire [7:0] t_r32_c29_8;
  wire [7:0] t_r32_c29_9;
  wire [7:0] t_r32_c29_10;
  wire [7:0] t_r32_c29_11;
  wire [7:0] t_r32_c29_12;
  wire [7:0] t_r32_c30_0;
  wire [7:0] t_r32_c30_1;
  wire [7:0] t_r32_c30_2;
  wire [7:0] t_r32_c30_3;
  wire [7:0] t_r32_c30_4;
  wire [7:0] t_r32_c30_5;
  wire [7:0] t_r32_c30_6;
  wire [7:0] t_r32_c30_7;
  wire [7:0] t_r32_c30_8;
  wire [7:0] t_r32_c30_9;
  wire [7:0] t_r32_c30_10;
  wire [7:0] t_r32_c30_11;
  wire [7:0] t_r32_c30_12;
  wire [7:0] t_r32_c31_0;
  wire [7:0] t_r32_c31_1;
  wire [7:0] t_r32_c31_2;
  wire [7:0] t_r32_c31_3;
  wire [7:0] t_r32_c31_4;
  wire [7:0] t_r32_c31_5;
  wire [7:0] t_r32_c31_6;
  wire [7:0] t_r32_c31_7;
  wire [7:0] t_r32_c31_8;
  wire [7:0] t_r32_c31_9;
  wire [7:0] t_r32_c31_10;
  wire [7:0] t_r32_c31_11;
  wire [7:0] t_r32_c31_12;
  wire [7:0] t_r32_c32_0;
  wire [7:0] t_r32_c32_1;
  wire [7:0] t_r32_c32_2;
  wire [7:0] t_r32_c32_3;
  wire [7:0] t_r32_c32_4;
  wire [7:0] t_r32_c32_5;
  wire [7:0] t_r32_c32_6;
  wire [7:0] t_r32_c32_7;
  wire [7:0] t_r32_c32_8;
  wire [7:0] t_r32_c32_9;
  wire [7:0] t_r32_c32_10;
  wire [7:0] t_r32_c32_11;
  wire [7:0] t_r32_c32_12;
  wire [7:0] t_r32_c33_0;
  wire [7:0] t_r32_c33_1;
  wire [7:0] t_r32_c33_2;
  wire [7:0] t_r32_c33_3;
  wire [7:0] t_r32_c33_4;
  wire [7:0] t_r32_c33_5;
  wire [7:0] t_r32_c33_6;
  wire [7:0] t_r32_c33_7;
  wire [7:0] t_r32_c33_8;
  wire [7:0] t_r32_c33_9;
  wire [7:0] t_r32_c33_10;
  wire [7:0] t_r32_c33_11;
  wire [7:0] t_r32_c33_12;
  wire [7:0] t_r32_c34_0;
  wire [7:0] t_r32_c34_1;
  wire [7:0] t_r32_c34_2;
  wire [7:0] t_r32_c34_3;
  wire [7:0] t_r32_c34_4;
  wire [7:0] t_r32_c34_5;
  wire [7:0] t_r32_c34_6;
  wire [7:0] t_r32_c34_7;
  wire [7:0] t_r32_c34_8;
  wire [7:0] t_r32_c34_9;
  wire [7:0] t_r32_c34_10;
  wire [7:0] t_r32_c34_11;
  wire [7:0] t_r32_c34_12;
  wire [7:0] t_r32_c35_0;
  wire [7:0] t_r32_c35_1;
  wire [7:0] t_r32_c35_2;
  wire [7:0] t_r32_c35_3;
  wire [7:0] t_r32_c35_4;
  wire [7:0] t_r32_c35_5;
  wire [7:0] t_r32_c35_6;
  wire [7:0] t_r32_c35_7;
  wire [7:0] t_r32_c35_8;
  wire [7:0] t_r32_c35_9;
  wire [7:0] t_r32_c35_10;
  wire [7:0] t_r32_c35_11;
  wire [7:0] t_r32_c35_12;
  wire [7:0] t_r32_c36_0;
  wire [7:0] t_r32_c36_1;
  wire [7:0] t_r32_c36_2;
  wire [7:0] t_r32_c36_3;
  wire [7:0] t_r32_c36_4;
  wire [7:0] t_r32_c36_5;
  wire [7:0] t_r32_c36_6;
  wire [7:0] t_r32_c36_7;
  wire [7:0] t_r32_c36_8;
  wire [7:0] t_r32_c36_9;
  wire [7:0] t_r32_c36_10;
  wire [7:0] t_r32_c36_11;
  wire [7:0] t_r32_c36_12;
  wire [7:0] t_r32_c37_0;
  wire [7:0] t_r32_c37_1;
  wire [7:0] t_r32_c37_2;
  wire [7:0] t_r32_c37_3;
  wire [7:0] t_r32_c37_4;
  wire [7:0] t_r32_c37_5;
  wire [7:0] t_r32_c37_6;
  wire [7:0] t_r32_c37_7;
  wire [7:0] t_r32_c37_8;
  wire [7:0] t_r32_c37_9;
  wire [7:0] t_r32_c37_10;
  wire [7:0] t_r32_c37_11;
  wire [7:0] t_r32_c37_12;
  wire [7:0] t_r32_c38_0;
  wire [7:0] t_r32_c38_1;
  wire [7:0] t_r32_c38_2;
  wire [7:0] t_r32_c38_3;
  wire [7:0] t_r32_c38_4;
  wire [7:0] t_r32_c38_5;
  wire [7:0] t_r32_c38_6;
  wire [7:0] t_r32_c38_7;
  wire [7:0] t_r32_c38_8;
  wire [7:0] t_r32_c38_9;
  wire [7:0] t_r32_c38_10;
  wire [7:0] t_r32_c38_11;
  wire [7:0] t_r32_c38_12;
  wire [7:0] t_r32_c39_0;
  wire [7:0] t_r32_c39_1;
  wire [7:0] t_r32_c39_2;
  wire [7:0] t_r32_c39_3;
  wire [7:0] t_r32_c39_4;
  wire [7:0] t_r32_c39_5;
  wire [7:0] t_r32_c39_6;
  wire [7:0] t_r32_c39_7;
  wire [7:0] t_r32_c39_8;
  wire [7:0] t_r32_c39_9;
  wire [7:0] t_r32_c39_10;
  wire [7:0] t_r32_c39_11;
  wire [7:0] t_r32_c39_12;
  wire [7:0] t_r32_c40_0;
  wire [7:0] t_r32_c40_1;
  wire [7:0] t_r32_c40_2;
  wire [7:0] t_r32_c40_3;
  wire [7:0] t_r32_c40_4;
  wire [7:0] t_r32_c40_5;
  wire [7:0] t_r32_c40_6;
  wire [7:0] t_r32_c40_7;
  wire [7:0] t_r32_c40_8;
  wire [7:0] t_r32_c40_9;
  wire [7:0] t_r32_c40_10;
  wire [7:0] t_r32_c40_11;
  wire [7:0] t_r32_c40_12;
  wire [7:0] t_r32_c41_0;
  wire [7:0] t_r32_c41_1;
  wire [7:0] t_r32_c41_2;
  wire [7:0] t_r32_c41_3;
  wire [7:0] t_r32_c41_4;
  wire [7:0] t_r32_c41_5;
  wire [7:0] t_r32_c41_6;
  wire [7:0] t_r32_c41_7;
  wire [7:0] t_r32_c41_8;
  wire [7:0] t_r32_c41_9;
  wire [7:0] t_r32_c41_10;
  wire [7:0] t_r32_c41_11;
  wire [7:0] t_r32_c41_12;
  wire [7:0] t_r32_c42_0;
  wire [7:0] t_r32_c42_1;
  wire [7:0] t_r32_c42_2;
  wire [7:0] t_r32_c42_3;
  wire [7:0] t_r32_c42_4;
  wire [7:0] t_r32_c42_5;
  wire [7:0] t_r32_c42_6;
  wire [7:0] t_r32_c42_7;
  wire [7:0] t_r32_c42_8;
  wire [7:0] t_r32_c42_9;
  wire [7:0] t_r32_c42_10;
  wire [7:0] t_r32_c42_11;
  wire [7:0] t_r32_c42_12;
  wire [7:0] t_r32_c43_0;
  wire [7:0] t_r32_c43_1;
  wire [7:0] t_r32_c43_2;
  wire [7:0] t_r32_c43_3;
  wire [7:0] t_r32_c43_4;
  wire [7:0] t_r32_c43_5;
  wire [7:0] t_r32_c43_6;
  wire [7:0] t_r32_c43_7;
  wire [7:0] t_r32_c43_8;
  wire [7:0] t_r32_c43_9;
  wire [7:0] t_r32_c43_10;
  wire [7:0] t_r32_c43_11;
  wire [7:0] t_r32_c43_12;
  wire [7:0] t_r32_c44_0;
  wire [7:0] t_r32_c44_1;
  wire [7:0] t_r32_c44_2;
  wire [7:0] t_r32_c44_3;
  wire [7:0] t_r32_c44_4;
  wire [7:0] t_r32_c44_5;
  wire [7:0] t_r32_c44_6;
  wire [7:0] t_r32_c44_7;
  wire [7:0] t_r32_c44_8;
  wire [7:0] t_r32_c44_9;
  wire [7:0] t_r32_c44_10;
  wire [7:0] t_r32_c44_11;
  wire [7:0] t_r32_c44_12;
  wire [7:0] t_r32_c45_0;
  wire [7:0] t_r32_c45_1;
  wire [7:0] t_r32_c45_2;
  wire [7:0] t_r32_c45_3;
  wire [7:0] t_r32_c45_4;
  wire [7:0] t_r32_c45_5;
  wire [7:0] t_r32_c45_6;
  wire [7:0] t_r32_c45_7;
  wire [7:0] t_r32_c45_8;
  wire [7:0] t_r32_c45_9;
  wire [7:0] t_r32_c45_10;
  wire [7:0] t_r32_c45_11;
  wire [7:0] t_r32_c45_12;
  wire [7:0] t_r32_c46_0;
  wire [7:0] t_r32_c46_1;
  wire [7:0] t_r32_c46_2;
  wire [7:0] t_r32_c46_3;
  wire [7:0] t_r32_c46_4;
  wire [7:0] t_r32_c46_5;
  wire [7:0] t_r32_c46_6;
  wire [7:0] t_r32_c46_7;
  wire [7:0] t_r32_c46_8;
  wire [7:0] t_r32_c46_9;
  wire [7:0] t_r32_c46_10;
  wire [7:0] t_r32_c46_11;
  wire [7:0] t_r32_c46_12;
  wire [7:0] t_r32_c47_0;
  wire [7:0] t_r32_c47_1;
  wire [7:0] t_r32_c47_2;
  wire [7:0] t_r32_c47_3;
  wire [7:0] t_r32_c47_4;
  wire [7:0] t_r32_c47_5;
  wire [7:0] t_r32_c47_6;
  wire [7:0] t_r32_c47_7;
  wire [7:0] t_r32_c47_8;
  wire [7:0] t_r32_c47_9;
  wire [7:0] t_r32_c47_10;
  wire [7:0] t_r32_c47_11;
  wire [7:0] t_r32_c47_12;
  wire [7:0] t_r32_c48_0;
  wire [7:0] t_r32_c48_1;
  wire [7:0] t_r32_c48_2;
  wire [7:0] t_r32_c48_3;
  wire [7:0] t_r32_c48_4;
  wire [7:0] t_r32_c48_5;
  wire [7:0] t_r32_c48_6;
  wire [7:0] t_r32_c48_7;
  wire [7:0] t_r32_c48_8;
  wire [7:0] t_r32_c48_9;
  wire [7:0] t_r32_c48_10;
  wire [7:0] t_r32_c48_11;
  wire [7:0] t_r32_c48_12;
  wire [7:0] t_r32_c49_0;
  wire [7:0] t_r32_c49_1;
  wire [7:0] t_r32_c49_2;
  wire [7:0] t_r32_c49_3;
  wire [7:0] t_r32_c49_4;
  wire [7:0] t_r32_c49_5;
  wire [7:0] t_r32_c49_6;
  wire [7:0] t_r32_c49_7;
  wire [7:0] t_r32_c49_8;
  wire [7:0] t_r32_c49_9;
  wire [7:0] t_r32_c49_10;
  wire [7:0] t_r32_c49_11;
  wire [7:0] t_r32_c49_12;
  wire [7:0] t_r32_c50_0;
  wire [7:0] t_r32_c50_1;
  wire [7:0] t_r32_c50_2;
  wire [7:0] t_r32_c50_3;
  wire [7:0] t_r32_c50_4;
  wire [7:0] t_r32_c50_5;
  wire [7:0] t_r32_c50_6;
  wire [7:0] t_r32_c50_7;
  wire [7:0] t_r32_c50_8;
  wire [7:0] t_r32_c50_9;
  wire [7:0] t_r32_c50_10;
  wire [7:0] t_r32_c50_11;
  wire [7:0] t_r32_c50_12;
  wire [7:0] t_r32_c51_0;
  wire [7:0] t_r32_c51_1;
  wire [7:0] t_r32_c51_2;
  wire [7:0] t_r32_c51_3;
  wire [7:0] t_r32_c51_4;
  wire [7:0] t_r32_c51_5;
  wire [7:0] t_r32_c51_6;
  wire [7:0] t_r32_c51_7;
  wire [7:0] t_r32_c51_8;
  wire [7:0] t_r32_c51_9;
  wire [7:0] t_r32_c51_10;
  wire [7:0] t_r32_c51_11;
  wire [7:0] t_r32_c51_12;
  wire [7:0] t_r32_c52_0;
  wire [7:0] t_r32_c52_1;
  wire [7:0] t_r32_c52_2;
  wire [7:0] t_r32_c52_3;
  wire [7:0] t_r32_c52_4;
  wire [7:0] t_r32_c52_5;
  wire [7:0] t_r32_c52_6;
  wire [7:0] t_r32_c52_7;
  wire [7:0] t_r32_c52_8;
  wire [7:0] t_r32_c52_9;
  wire [7:0] t_r32_c52_10;
  wire [7:0] t_r32_c52_11;
  wire [7:0] t_r32_c52_12;
  wire [7:0] t_r32_c53_0;
  wire [7:0] t_r32_c53_1;
  wire [7:0] t_r32_c53_2;
  wire [7:0] t_r32_c53_3;
  wire [7:0] t_r32_c53_4;
  wire [7:0] t_r32_c53_5;
  wire [7:0] t_r32_c53_6;
  wire [7:0] t_r32_c53_7;
  wire [7:0] t_r32_c53_8;
  wire [7:0] t_r32_c53_9;
  wire [7:0] t_r32_c53_10;
  wire [7:0] t_r32_c53_11;
  wire [7:0] t_r32_c53_12;
  wire [7:0] t_r32_c54_0;
  wire [7:0] t_r32_c54_1;
  wire [7:0] t_r32_c54_2;
  wire [7:0] t_r32_c54_3;
  wire [7:0] t_r32_c54_4;
  wire [7:0] t_r32_c54_5;
  wire [7:0] t_r32_c54_6;
  wire [7:0] t_r32_c54_7;
  wire [7:0] t_r32_c54_8;
  wire [7:0] t_r32_c54_9;
  wire [7:0] t_r32_c54_10;
  wire [7:0] t_r32_c54_11;
  wire [7:0] t_r32_c54_12;
  wire [7:0] t_r32_c55_0;
  wire [7:0] t_r32_c55_1;
  wire [7:0] t_r32_c55_2;
  wire [7:0] t_r32_c55_3;
  wire [7:0] t_r32_c55_4;
  wire [7:0] t_r32_c55_5;
  wire [7:0] t_r32_c55_6;
  wire [7:0] t_r32_c55_7;
  wire [7:0] t_r32_c55_8;
  wire [7:0] t_r32_c55_9;
  wire [7:0] t_r32_c55_10;
  wire [7:0] t_r32_c55_11;
  wire [7:0] t_r32_c55_12;
  wire [7:0] t_r32_c56_0;
  wire [7:0] t_r32_c56_1;
  wire [7:0] t_r32_c56_2;
  wire [7:0] t_r32_c56_3;
  wire [7:0] t_r32_c56_4;
  wire [7:0] t_r32_c56_5;
  wire [7:0] t_r32_c56_6;
  wire [7:0] t_r32_c56_7;
  wire [7:0] t_r32_c56_8;
  wire [7:0] t_r32_c56_9;
  wire [7:0] t_r32_c56_10;
  wire [7:0] t_r32_c56_11;
  wire [7:0] t_r32_c56_12;
  wire [7:0] t_r32_c57_0;
  wire [7:0] t_r32_c57_1;
  wire [7:0] t_r32_c57_2;
  wire [7:0] t_r32_c57_3;
  wire [7:0] t_r32_c57_4;
  wire [7:0] t_r32_c57_5;
  wire [7:0] t_r32_c57_6;
  wire [7:0] t_r32_c57_7;
  wire [7:0] t_r32_c57_8;
  wire [7:0] t_r32_c57_9;
  wire [7:0] t_r32_c57_10;
  wire [7:0] t_r32_c57_11;
  wire [7:0] t_r32_c57_12;
  wire [7:0] t_r32_c58_0;
  wire [7:0] t_r32_c58_1;
  wire [7:0] t_r32_c58_2;
  wire [7:0] t_r32_c58_3;
  wire [7:0] t_r32_c58_4;
  wire [7:0] t_r32_c58_5;
  wire [7:0] t_r32_c58_6;
  wire [7:0] t_r32_c58_7;
  wire [7:0] t_r32_c58_8;
  wire [7:0] t_r32_c58_9;
  wire [7:0] t_r32_c58_10;
  wire [7:0] t_r32_c58_11;
  wire [7:0] t_r32_c58_12;
  wire [7:0] t_r32_c59_0;
  wire [7:0] t_r32_c59_1;
  wire [7:0] t_r32_c59_2;
  wire [7:0] t_r32_c59_3;
  wire [7:0] t_r32_c59_4;
  wire [7:0] t_r32_c59_5;
  wire [7:0] t_r32_c59_6;
  wire [7:0] t_r32_c59_7;
  wire [7:0] t_r32_c59_8;
  wire [7:0] t_r32_c59_9;
  wire [7:0] t_r32_c59_10;
  wire [7:0] t_r32_c59_11;
  wire [7:0] t_r32_c59_12;
  wire [7:0] t_r32_c60_0;
  wire [7:0] t_r32_c60_1;
  wire [7:0] t_r32_c60_2;
  wire [7:0] t_r32_c60_3;
  wire [7:0] t_r32_c60_4;
  wire [7:0] t_r32_c60_5;
  wire [7:0] t_r32_c60_6;
  wire [7:0] t_r32_c60_7;
  wire [7:0] t_r32_c60_8;
  wire [7:0] t_r32_c60_9;
  wire [7:0] t_r32_c60_10;
  wire [7:0] t_r32_c60_11;
  wire [7:0] t_r32_c60_12;
  wire [7:0] t_r32_c61_0;
  wire [7:0] t_r32_c61_1;
  wire [7:0] t_r32_c61_2;
  wire [7:0] t_r32_c61_3;
  wire [7:0] t_r32_c61_4;
  wire [7:0] t_r32_c61_5;
  wire [7:0] t_r32_c61_6;
  wire [7:0] t_r32_c61_7;
  wire [7:0] t_r32_c61_8;
  wire [7:0] t_r32_c61_9;
  wire [7:0] t_r32_c61_10;
  wire [7:0] t_r32_c61_11;
  wire [7:0] t_r32_c61_12;
  wire [7:0] t_r32_c62_0;
  wire [7:0] t_r32_c62_1;
  wire [7:0] t_r32_c62_2;
  wire [7:0] t_r32_c62_3;
  wire [7:0] t_r32_c62_4;
  wire [7:0] t_r32_c62_5;
  wire [7:0] t_r32_c62_6;
  wire [7:0] t_r32_c62_7;
  wire [7:0] t_r32_c62_8;
  wire [7:0] t_r32_c62_9;
  wire [7:0] t_r32_c62_10;
  wire [7:0] t_r32_c62_11;
  wire [7:0] t_r32_c62_12;
  wire [7:0] t_r32_c63_0;
  wire [7:0] t_r32_c63_1;
  wire [7:0] t_r32_c63_2;
  wire [7:0] t_r32_c63_3;
  wire [7:0] t_r32_c63_4;
  wire [7:0] t_r32_c63_5;
  wire [7:0] t_r32_c63_6;
  wire [7:0] t_r32_c63_7;
  wire [7:0] t_r32_c63_8;
  wire [7:0] t_r32_c63_9;
  wire [7:0] t_r32_c63_10;
  wire [7:0] t_r32_c63_11;
  wire [7:0] t_r32_c63_12;
  wire [7:0] t_r32_c64_0;
  wire [7:0] t_r32_c64_1;
  wire [7:0] t_r32_c64_2;
  wire [7:0] t_r32_c64_3;
  wire [7:0] t_r32_c64_4;
  wire [7:0] t_r32_c64_5;
  wire [7:0] t_r32_c64_6;
  wire [7:0] t_r32_c64_7;
  wire [7:0] t_r32_c64_8;
  wire [7:0] t_r32_c64_9;
  wire [7:0] t_r32_c64_10;
  wire [7:0] t_r32_c64_11;
  wire [7:0] t_r32_c64_12;
  wire [7:0] t_r32_c65_0;
  wire [7:0] t_r32_c65_1;
  wire [7:0] t_r32_c65_2;
  wire [7:0] t_r32_c65_3;
  wire [7:0] t_r32_c65_4;
  wire [7:0] t_r32_c65_5;
  wire [7:0] t_r32_c65_6;
  wire [7:0] t_r32_c65_7;
  wire [7:0] t_r32_c65_8;
  wire [7:0] t_r32_c65_9;
  wire [7:0] t_r32_c65_10;
  wire [7:0] t_r32_c65_11;
  wire [7:0] t_r32_c65_12;
  wire [7:0] t_r33_c0_0;
  wire [7:0] t_r33_c0_1;
  wire [7:0] t_r33_c0_2;
  wire [7:0] t_r33_c0_3;
  wire [7:0] t_r33_c0_4;
  wire [7:0] t_r33_c0_5;
  wire [7:0] t_r33_c0_6;
  wire [7:0] t_r33_c0_7;
  wire [7:0] t_r33_c0_8;
  wire [7:0] t_r33_c0_9;
  wire [7:0] t_r33_c0_10;
  wire [7:0] t_r33_c0_11;
  wire [7:0] t_r33_c0_12;
  wire [7:0] t_r33_c1_0;
  wire [7:0] t_r33_c1_1;
  wire [7:0] t_r33_c1_2;
  wire [7:0] t_r33_c1_3;
  wire [7:0] t_r33_c1_4;
  wire [7:0] t_r33_c1_5;
  wire [7:0] t_r33_c1_6;
  wire [7:0] t_r33_c1_7;
  wire [7:0] t_r33_c1_8;
  wire [7:0] t_r33_c1_9;
  wire [7:0] t_r33_c1_10;
  wire [7:0] t_r33_c1_11;
  wire [7:0] t_r33_c1_12;
  wire [7:0] t_r33_c2_0;
  wire [7:0] t_r33_c2_1;
  wire [7:0] t_r33_c2_2;
  wire [7:0] t_r33_c2_3;
  wire [7:0] t_r33_c2_4;
  wire [7:0] t_r33_c2_5;
  wire [7:0] t_r33_c2_6;
  wire [7:0] t_r33_c2_7;
  wire [7:0] t_r33_c2_8;
  wire [7:0] t_r33_c2_9;
  wire [7:0] t_r33_c2_10;
  wire [7:0] t_r33_c2_11;
  wire [7:0] t_r33_c2_12;
  wire [7:0] t_r33_c3_0;
  wire [7:0] t_r33_c3_1;
  wire [7:0] t_r33_c3_2;
  wire [7:0] t_r33_c3_3;
  wire [7:0] t_r33_c3_4;
  wire [7:0] t_r33_c3_5;
  wire [7:0] t_r33_c3_6;
  wire [7:0] t_r33_c3_7;
  wire [7:0] t_r33_c3_8;
  wire [7:0] t_r33_c3_9;
  wire [7:0] t_r33_c3_10;
  wire [7:0] t_r33_c3_11;
  wire [7:0] t_r33_c3_12;
  wire [7:0] t_r33_c4_0;
  wire [7:0] t_r33_c4_1;
  wire [7:0] t_r33_c4_2;
  wire [7:0] t_r33_c4_3;
  wire [7:0] t_r33_c4_4;
  wire [7:0] t_r33_c4_5;
  wire [7:0] t_r33_c4_6;
  wire [7:0] t_r33_c4_7;
  wire [7:0] t_r33_c4_8;
  wire [7:0] t_r33_c4_9;
  wire [7:0] t_r33_c4_10;
  wire [7:0] t_r33_c4_11;
  wire [7:0] t_r33_c4_12;
  wire [7:0] t_r33_c5_0;
  wire [7:0] t_r33_c5_1;
  wire [7:0] t_r33_c5_2;
  wire [7:0] t_r33_c5_3;
  wire [7:0] t_r33_c5_4;
  wire [7:0] t_r33_c5_5;
  wire [7:0] t_r33_c5_6;
  wire [7:0] t_r33_c5_7;
  wire [7:0] t_r33_c5_8;
  wire [7:0] t_r33_c5_9;
  wire [7:0] t_r33_c5_10;
  wire [7:0] t_r33_c5_11;
  wire [7:0] t_r33_c5_12;
  wire [7:0] t_r33_c6_0;
  wire [7:0] t_r33_c6_1;
  wire [7:0] t_r33_c6_2;
  wire [7:0] t_r33_c6_3;
  wire [7:0] t_r33_c6_4;
  wire [7:0] t_r33_c6_5;
  wire [7:0] t_r33_c6_6;
  wire [7:0] t_r33_c6_7;
  wire [7:0] t_r33_c6_8;
  wire [7:0] t_r33_c6_9;
  wire [7:0] t_r33_c6_10;
  wire [7:0] t_r33_c6_11;
  wire [7:0] t_r33_c6_12;
  wire [7:0] t_r33_c7_0;
  wire [7:0] t_r33_c7_1;
  wire [7:0] t_r33_c7_2;
  wire [7:0] t_r33_c7_3;
  wire [7:0] t_r33_c7_4;
  wire [7:0] t_r33_c7_5;
  wire [7:0] t_r33_c7_6;
  wire [7:0] t_r33_c7_7;
  wire [7:0] t_r33_c7_8;
  wire [7:0] t_r33_c7_9;
  wire [7:0] t_r33_c7_10;
  wire [7:0] t_r33_c7_11;
  wire [7:0] t_r33_c7_12;
  wire [7:0] t_r33_c8_0;
  wire [7:0] t_r33_c8_1;
  wire [7:0] t_r33_c8_2;
  wire [7:0] t_r33_c8_3;
  wire [7:0] t_r33_c8_4;
  wire [7:0] t_r33_c8_5;
  wire [7:0] t_r33_c8_6;
  wire [7:0] t_r33_c8_7;
  wire [7:0] t_r33_c8_8;
  wire [7:0] t_r33_c8_9;
  wire [7:0] t_r33_c8_10;
  wire [7:0] t_r33_c8_11;
  wire [7:0] t_r33_c8_12;
  wire [7:0] t_r33_c9_0;
  wire [7:0] t_r33_c9_1;
  wire [7:0] t_r33_c9_2;
  wire [7:0] t_r33_c9_3;
  wire [7:0] t_r33_c9_4;
  wire [7:0] t_r33_c9_5;
  wire [7:0] t_r33_c9_6;
  wire [7:0] t_r33_c9_7;
  wire [7:0] t_r33_c9_8;
  wire [7:0] t_r33_c9_9;
  wire [7:0] t_r33_c9_10;
  wire [7:0] t_r33_c9_11;
  wire [7:0] t_r33_c9_12;
  wire [7:0] t_r33_c10_0;
  wire [7:0] t_r33_c10_1;
  wire [7:0] t_r33_c10_2;
  wire [7:0] t_r33_c10_3;
  wire [7:0] t_r33_c10_4;
  wire [7:0] t_r33_c10_5;
  wire [7:0] t_r33_c10_6;
  wire [7:0] t_r33_c10_7;
  wire [7:0] t_r33_c10_8;
  wire [7:0] t_r33_c10_9;
  wire [7:0] t_r33_c10_10;
  wire [7:0] t_r33_c10_11;
  wire [7:0] t_r33_c10_12;
  wire [7:0] t_r33_c11_0;
  wire [7:0] t_r33_c11_1;
  wire [7:0] t_r33_c11_2;
  wire [7:0] t_r33_c11_3;
  wire [7:0] t_r33_c11_4;
  wire [7:0] t_r33_c11_5;
  wire [7:0] t_r33_c11_6;
  wire [7:0] t_r33_c11_7;
  wire [7:0] t_r33_c11_8;
  wire [7:0] t_r33_c11_9;
  wire [7:0] t_r33_c11_10;
  wire [7:0] t_r33_c11_11;
  wire [7:0] t_r33_c11_12;
  wire [7:0] t_r33_c12_0;
  wire [7:0] t_r33_c12_1;
  wire [7:0] t_r33_c12_2;
  wire [7:0] t_r33_c12_3;
  wire [7:0] t_r33_c12_4;
  wire [7:0] t_r33_c12_5;
  wire [7:0] t_r33_c12_6;
  wire [7:0] t_r33_c12_7;
  wire [7:0] t_r33_c12_8;
  wire [7:0] t_r33_c12_9;
  wire [7:0] t_r33_c12_10;
  wire [7:0] t_r33_c12_11;
  wire [7:0] t_r33_c12_12;
  wire [7:0] t_r33_c13_0;
  wire [7:0] t_r33_c13_1;
  wire [7:0] t_r33_c13_2;
  wire [7:0] t_r33_c13_3;
  wire [7:0] t_r33_c13_4;
  wire [7:0] t_r33_c13_5;
  wire [7:0] t_r33_c13_6;
  wire [7:0] t_r33_c13_7;
  wire [7:0] t_r33_c13_8;
  wire [7:0] t_r33_c13_9;
  wire [7:0] t_r33_c13_10;
  wire [7:0] t_r33_c13_11;
  wire [7:0] t_r33_c13_12;
  wire [7:0] t_r33_c14_0;
  wire [7:0] t_r33_c14_1;
  wire [7:0] t_r33_c14_2;
  wire [7:0] t_r33_c14_3;
  wire [7:0] t_r33_c14_4;
  wire [7:0] t_r33_c14_5;
  wire [7:0] t_r33_c14_6;
  wire [7:0] t_r33_c14_7;
  wire [7:0] t_r33_c14_8;
  wire [7:0] t_r33_c14_9;
  wire [7:0] t_r33_c14_10;
  wire [7:0] t_r33_c14_11;
  wire [7:0] t_r33_c14_12;
  wire [7:0] t_r33_c15_0;
  wire [7:0] t_r33_c15_1;
  wire [7:0] t_r33_c15_2;
  wire [7:0] t_r33_c15_3;
  wire [7:0] t_r33_c15_4;
  wire [7:0] t_r33_c15_5;
  wire [7:0] t_r33_c15_6;
  wire [7:0] t_r33_c15_7;
  wire [7:0] t_r33_c15_8;
  wire [7:0] t_r33_c15_9;
  wire [7:0] t_r33_c15_10;
  wire [7:0] t_r33_c15_11;
  wire [7:0] t_r33_c15_12;
  wire [7:0] t_r33_c16_0;
  wire [7:0] t_r33_c16_1;
  wire [7:0] t_r33_c16_2;
  wire [7:0] t_r33_c16_3;
  wire [7:0] t_r33_c16_4;
  wire [7:0] t_r33_c16_5;
  wire [7:0] t_r33_c16_6;
  wire [7:0] t_r33_c16_7;
  wire [7:0] t_r33_c16_8;
  wire [7:0] t_r33_c16_9;
  wire [7:0] t_r33_c16_10;
  wire [7:0] t_r33_c16_11;
  wire [7:0] t_r33_c16_12;
  wire [7:0] t_r33_c17_0;
  wire [7:0] t_r33_c17_1;
  wire [7:0] t_r33_c17_2;
  wire [7:0] t_r33_c17_3;
  wire [7:0] t_r33_c17_4;
  wire [7:0] t_r33_c17_5;
  wire [7:0] t_r33_c17_6;
  wire [7:0] t_r33_c17_7;
  wire [7:0] t_r33_c17_8;
  wire [7:0] t_r33_c17_9;
  wire [7:0] t_r33_c17_10;
  wire [7:0] t_r33_c17_11;
  wire [7:0] t_r33_c17_12;
  wire [7:0] t_r33_c18_0;
  wire [7:0] t_r33_c18_1;
  wire [7:0] t_r33_c18_2;
  wire [7:0] t_r33_c18_3;
  wire [7:0] t_r33_c18_4;
  wire [7:0] t_r33_c18_5;
  wire [7:0] t_r33_c18_6;
  wire [7:0] t_r33_c18_7;
  wire [7:0] t_r33_c18_8;
  wire [7:0] t_r33_c18_9;
  wire [7:0] t_r33_c18_10;
  wire [7:0] t_r33_c18_11;
  wire [7:0] t_r33_c18_12;
  wire [7:0] t_r33_c19_0;
  wire [7:0] t_r33_c19_1;
  wire [7:0] t_r33_c19_2;
  wire [7:0] t_r33_c19_3;
  wire [7:0] t_r33_c19_4;
  wire [7:0] t_r33_c19_5;
  wire [7:0] t_r33_c19_6;
  wire [7:0] t_r33_c19_7;
  wire [7:0] t_r33_c19_8;
  wire [7:0] t_r33_c19_9;
  wire [7:0] t_r33_c19_10;
  wire [7:0] t_r33_c19_11;
  wire [7:0] t_r33_c19_12;
  wire [7:0] t_r33_c20_0;
  wire [7:0] t_r33_c20_1;
  wire [7:0] t_r33_c20_2;
  wire [7:0] t_r33_c20_3;
  wire [7:0] t_r33_c20_4;
  wire [7:0] t_r33_c20_5;
  wire [7:0] t_r33_c20_6;
  wire [7:0] t_r33_c20_7;
  wire [7:0] t_r33_c20_8;
  wire [7:0] t_r33_c20_9;
  wire [7:0] t_r33_c20_10;
  wire [7:0] t_r33_c20_11;
  wire [7:0] t_r33_c20_12;
  wire [7:0] t_r33_c21_0;
  wire [7:0] t_r33_c21_1;
  wire [7:0] t_r33_c21_2;
  wire [7:0] t_r33_c21_3;
  wire [7:0] t_r33_c21_4;
  wire [7:0] t_r33_c21_5;
  wire [7:0] t_r33_c21_6;
  wire [7:0] t_r33_c21_7;
  wire [7:0] t_r33_c21_8;
  wire [7:0] t_r33_c21_9;
  wire [7:0] t_r33_c21_10;
  wire [7:0] t_r33_c21_11;
  wire [7:0] t_r33_c21_12;
  wire [7:0] t_r33_c22_0;
  wire [7:0] t_r33_c22_1;
  wire [7:0] t_r33_c22_2;
  wire [7:0] t_r33_c22_3;
  wire [7:0] t_r33_c22_4;
  wire [7:0] t_r33_c22_5;
  wire [7:0] t_r33_c22_6;
  wire [7:0] t_r33_c22_7;
  wire [7:0] t_r33_c22_8;
  wire [7:0] t_r33_c22_9;
  wire [7:0] t_r33_c22_10;
  wire [7:0] t_r33_c22_11;
  wire [7:0] t_r33_c22_12;
  wire [7:0] t_r33_c23_0;
  wire [7:0] t_r33_c23_1;
  wire [7:0] t_r33_c23_2;
  wire [7:0] t_r33_c23_3;
  wire [7:0] t_r33_c23_4;
  wire [7:0] t_r33_c23_5;
  wire [7:0] t_r33_c23_6;
  wire [7:0] t_r33_c23_7;
  wire [7:0] t_r33_c23_8;
  wire [7:0] t_r33_c23_9;
  wire [7:0] t_r33_c23_10;
  wire [7:0] t_r33_c23_11;
  wire [7:0] t_r33_c23_12;
  wire [7:0] t_r33_c24_0;
  wire [7:0] t_r33_c24_1;
  wire [7:0] t_r33_c24_2;
  wire [7:0] t_r33_c24_3;
  wire [7:0] t_r33_c24_4;
  wire [7:0] t_r33_c24_5;
  wire [7:0] t_r33_c24_6;
  wire [7:0] t_r33_c24_7;
  wire [7:0] t_r33_c24_8;
  wire [7:0] t_r33_c24_9;
  wire [7:0] t_r33_c24_10;
  wire [7:0] t_r33_c24_11;
  wire [7:0] t_r33_c24_12;
  wire [7:0] t_r33_c25_0;
  wire [7:0] t_r33_c25_1;
  wire [7:0] t_r33_c25_2;
  wire [7:0] t_r33_c25_3;
  wire [7:0] t_r33_c25_4;
  wire [7:0] t_r33_c25_5;
  wire [7:0] t_r33_c25_6;
  wire [7:0] t_r33_c25_7;
  wire [7:0] t_r33_c25_8;
  wire [7:0] t_r33_c25_9;
  wire [7:0] t_r33_c25_10;
  wire [7:0] t_r33_c25_11;
  wire [7:0] t_r33_c25_12;
  wire [7:0] t_r33_c26_0;
  wire [7:0] t_r33_c26_1;
  wire [7:0] t_r33_c26_2;
  wire [7:0] t_r33_c26_3;
  wire [7:0] t_r33_c26_4;
  wire [7:0] t_r33_c26_5;
  wire [7:0] t_r33_c26_6;
  wire [7:0] t_r33_c26_7;
  wire [7:0] t_r33_c26_8;
  wire [7:0] t_r33_c26_9;
  wire [7:0] t_r33_c26_10;
  wire [7:0] t_r33_c26_11;
  wire [7:0] t_r33_c26_12;
  wire [7:0] t_r33_c27_0;
  wire [7:0] t_r33_c27_1;
  wire [7:0] t_r33_c27_2;
  wire [7:0] t_r33_c27_3;
  wire [7:0] t_r33_c27_4;
  wire [7:0] t_r33_c27_5;
  wire [7:0] t_r33_c27_6;
  wire [7:0] t_r33_c27_7;
  wire [7:0] t_r33_c27_8;
  wire [7:0] t_r33_c27_9;
  wire [7:0] t_r33_c27_10;
  wire [7:0] t_r33_c27_11;
  wire [7:0] t_r33_c27_12;
  wire [7:0] t_r33_c28_0;
  wire [7:0] t_r33_c28_1;
  wire [7:0] t_r33_c28_2;
  wire [7:0] t_r33_c28_3;
  wire [7:0] t_r33_c28_4;
  wire [7:0] t_r33_c28_5;
  wire [7:0] t_r33_c28_6;
  wire [7:0] t_r33_c28_7;
  wire [7:0] t_r33_c28_8;
  wire [7:0] t_r33_c28_9;
  wire [7:0] t_r33_c28_10;
  wire [7:0] t_r33_c28_11;
  wire [7:0] t_r33_c28_12;
  wire [7:0] t_r33_c29_0;
  wire [7:0] t_r33_c29_1;
  wire [7:0] t_r33_c29_2;
  wire [7:0] t_r33_c29_3;
  wire [7:0] t_r33_c29_4;
  wire [7:0] t_r33_c29_5;
  wire [7:0] t_r33_c29_6;
  wire [7:0] t_r33_c29_7;
  wire [7:0] t_r33_c29_8;
  wire [7:0] t_r33_c29_9;
  wire [7:0] t_r33_c29_10;
  wire [7:0] t_r33_c29_11;
  wire [7:0] t_r33_c29_12;
  wire [7:0] t_r33_c30_0;
  wire [7:0] t_r33_c30_1;
  wire [7:0] t_r33_c30_2;
  wire [7:0] t_r33_c30_3;
  wire [7:0] t_r33_c30_4;
  wire [7:0] t_r33_c30_5;
  wire [7:0] t_r33_c30_6;
  wire [7:0] t_r33_c30_7;
  wire [7:0] t_r33_c30_8;
  wire [7:0] t_r33_c30_9;
  wire [7:0] t_r33_c30_10;
  wire [7:0] t_r33_c30_11;
  wire [7:0] t_r33_c30_12;
  wire [7:0] t_r33_c31_0;
  wire [7:0] t_r33_c31_1;
  wire [7:0] t_r33_c31_2;
  wire [7:0] t_r33_c31_3;
  wire [7:0] t_r33_c31_4;
  wire [7:0] t_r33_c31_5;
  wire [7:0] t_r33_c31_6;
  wire [7:0] t_r33_c31_7;
  wire [7:0] t_r33_c31_8;
  wire [7:0] t_r33_c31_9;
  wire [7:0] t_r33_c31_10;
  wire [7:0] t_r33_c31_11;
  wire [7:0] t_r33_c31_12;
  wire [7:0] t_r33_c32_0;
  wire [7:0] t_r33_c32_1;
  wire [7:0] t_r33_c32_2;
  wire [7:0] t_r33_c32_3;
  wire [7:0] t_r33_c32_4;
  wire [7:0] t_r33_c32_5;
  wire [7:0] t_r33_c32_6;
  wire [7:0] t_r33_c32_7;
  wire [7:0] t_r33_c32_8;
  wire [7:0] t_r33_c32_9;
  wire [7:0] t_r33_c32_10;
  wire [7:0] t_r33_c32_11;
  wire [7:0] t_r33_c32_12;
  wire [7:0] t_r33_c33_0;
  wire [7:0] t_r33_c33_1;
  wire [7:0] t_r33_c33_2;
  wire [7:0] t_r33_c33_3;
  wire [7:0] t_r33_c33_4;
  wire [7:0] t_r33_c33_5;
  wire [7:0] t_r33_c33_6;
  wire [7:0] t_r33_c33_7;
  wire [7:0] t_r33_c33_8;
  wire [7:0] t_r33_c33_9;
  wire [7:0] t_r33_c33_10;
  wire [7:0] t_r33_c33_11;
  wire [7:0] t_r33_c33_12;
  wire [7:0] t_r33_c34_0;
  wire [7:0] t_r33_c34_1;
  wire [7:0] t_r33_c34_2;
  wire [7:0] t_r33_c34_3;
  wire [7:0] t_r33_c34_4;
  wire [7:0] t_r33_c34_5;
  wire [7:0] t_r33_c34_6;
  wire [7:0] t_r33_c34_7;
  wire [7:0] t_r33_c34_8;
  wire [7:0] t_r33_c34_9;
  wire [7:0] t_r33_c34_10;
  wire [7:0] t_r33_c34_11;
  wire [7:0] t_r33_c34_12;
  wire [7:0] t_r33_c35_0;
  wire [7:0] t_r33_c35_1;
  wire [7:0] t_r33_c35_2;
  wire [7:0] t_r33_c35_3;
  wire [7:0] t_r33_c35_4;
  wire [7:0] t_r33_c35_5;
  wire [7:0] t_r33_c35_6;
  wire [7:0] t_r33_c35_7;
  wire [7:0] t_r33_c35_8;
  wire [7:0] t_r33_c35_9;
  wire [7:0] t_r33_c35_10;
  wire [7:0] t_r33_c35_11;
  wire [7:0] t_r33_c35_12;
  wire [7:0] t_r33_c36_0;
  wire [7:0] t_r33_c36_1;
  wire [7:0] t_r33_c36_2;
  wire [7:0] t_r33_c36_3;
  wire [7:0] t_r33_c36_4;
  wire [7:0] t_r33_c36_5;
  wire [7:0] t_r33_c36_6;
  wire [7:0] t_r33_c36_7;
  wire [7:0] t_r33_c36_8;
  wire [7:0] t_r33_c36_9;
  wire [7:0] t_r33_c36_10;
  wire [7:0] t_r33_c36_11;
  wire [7:0] t_r33_c36_12;
  wire [7:0] t_r33_c37_0;
  wire [7:0] t_r33_c37_1;
  wire [7:0] t_r33_c37_2;
  wire [7:0] t_r33_c37_3;
  wire [7:0] t_r33_c37_4;
  wire [7:0] t_r33_c37_5;
  wire [7:0] t_r33_c37_6;
  wire [7:0] t_r33_c37_7;
  wire [7:0] t_r33_c37_8;
  wire [7:0] t_r33_c37_9;
  wire [7:0] t_r33_c37_10;
  wire [7:0] t_r33_c37_11;
  wire [7:0] t_r33_c37_12;
  wire [7:0] t_r33_c38_0;
  wire [7:0] t_r33_c38_1;
  wire [7:0] t_r33_c38_2;
  wire [7:0] t_r33_c38_3;
  wire [7:0] t_r33_c38_4;
  wire [7:0] t_r33_c38_5;
  wire [7:0] t_r33_c38_6;
  wire [7:0] t_r33_c38_7;
  wire [7:0] t_r33_c38_8;
  wire [7:0] t_r33_c38_9;
  wire [7:0] t_r33_c38_10;
  wire [7:0] t_r33_c38_11;
  wire [7:0] t_r33_c38_12;
  wire [7:0] t_r33_c39_0;
  wire [7:0] t_r33_c39_1;
  wire [7:0] t_r33_c39_2;
  wire [7:0] t_r33_c39_3;
  wire [7:0] t_r33_c39_4;
  wire [7:0] t_r33_c39_5;
  wire [7:0] t_r33_c39_6;
  wire [7:0] t_r33_c39_7;
  wire [7:0] t_r33_c39_8;
  wire [7:0] t_r33_c39_9;
  wire [7:0] t_r33_c39_10;
  wire [7:0] t_r33_c39_11;
  wire [7:0] t_r33_c39_12;
  wire [7:0] t_r33_c40_0;
  wire [7:0] t_r33_c40_1;
  wire [7:0] t_r33_c40_2;
  wire [7:0] t_r33_c40_3;
  wire [7:0] t_r33_c40_4;
  wire [7:0] t_r33_c40_5;
  wire [7:0] t_r33_c40_6;
  wire [7:0] t_r33_c40_7;
  wire [7:0] t_r33_c40_8;
  wire [7:0] t_r33_c40_9;
  wire [7:0] t_r33_c40_10;
  wire [7:0] t_r33_c40_11;
  wire [7:0] t_r33_c40_12;
  wire [7:0] t_r33_c41_0;
  wire [7:0] t_r33_c41_1;
  wire [7:0] t_r33_c41_2;
  wire [7:0] t_r33_c41_3;
  wire [7:0] t_r33_c41_4;
  wire [7:0] t_r33_c41_5;
  wire [7:0] t_r33_c41_6;
  wire [7:0] t_r33_c41_7;
  wire [7:0] t_r33_c41_8;
  wire [7:0] t_r33_c41_9;
  wire [7:0] t_r33_c41_10;
  wire [7:0] t_r33_c41_11;
  wire [7:0] t_r33_c41_12;
  wire [7:0] t_r33_c42_0;
  wire [7:0] t_r33_c42_1;
  wire [7:0] t_r33_c42_2;
  wire [7:0] t_r33_c42_3;
  wire [7:0] t_r33_c42_4;
  wire [7:0] t_r33_c42_5;
  wire [7:0] t_r33_c42_6;
  wire [7:0] t_r33_c42_7;
  wire [7:0] t_r33_c42_8;
  wire [7:0] t_r33_c42_9;
  wire [7:0] t_r33_c42_10;
  wire [7:0] t_r33_c42_11;
  wire [7:0] t_r33_c42_12;
  wire [7:0] t_r33_c43_0;
  wire [7:0] t_r33_c43_1;
  wire [7:0] t_r33_c43_2;
  wire [7:0] t_r33_c43_3;
  wire [7:0] t_r33_c43_4;
  wire [7:0] t_r33_c43_5;
  wire [7:0] t_r33_c43_6;
  wire [7:0] t_r33_c43_7;
  wire [7:0] t_r33_c43_8;
  wire [7:0] t_r33_c43_9;
  wire [7:0] t_r33_c43_10;
  wire [7:0] t_r33_c43_11;
  wire [7:0] t_r33_c43_12;
  wire [7:0] t_r33_c44_0;
  wire [7:0] t_r33_c44_1;
  wire [7:0] t_r33_c44_2;
  wire [7:0] t_r33_c44_3;
  wire [7:0] t_r33_c44_4;
  wire [7:0] t_r33_c44_5;
  wire [7:0] t_r33_c44_6;
  wire [7:0] t_r33_c44_7;
  wire [7:0] t_r33_c44_8;
  wire [7:0] t_r33_c44_9;
  wire [7:0] t_r33_c44_10;
  wire [7:0] t_r33_c44_11;
  wire [7:0] t_r33_c44_12;
  wire [7:0] t_r33_c45_0;
  wire [7:0] t_r33_c45_1;
  wire [7:0] t_r33_c45_2;
  wire [7:0] t_r33_c45_3;
  wire [7:0] t_r33_c45_4;
  wire [7:0] t_r33_c45_5;
  wire [7:0] t_r33_c45_6;
  wire [7:0] t_r33_c45_7;
  wire [7:0] t_r33_c45_8;
  wire [7:0] t_r33_c45_9;
  wire [7:0] t_r33_c45_10;
  wire [7:0] t_r33_c45_11;
  wire [7:0] t_r33_c45_12;
  wire [7:0] t_r33_c46_0;
  wire [7:0] t_r33_c46_1;
  wire [7:0] t_r33_c46_2;
  wire [7:0] t_r33_c46_3;
  wire [7:0] t_r33_c46_4;
  wire [7:0] t_r33_c46_5;
  wire [7:0] t_r33_c46_6;
  wire [7:0] t_r33_c46_7;
  wire [7:0] t_r33_c46_8;
  wire [7:0] t_r33_c46_9;
  wire [7:0] t_r33_c46_10;
  wire [7:0] t_r33_c46_11;
  wire [7:0] t_r33_c46_12;
  wire [7:0] t_r33_c47_0;
  wire [7:0] t_r33_c47_1;
  wire [7:0] t_r33_c47_2;
  wire [7:0] t_r33_c47_3;
  wire [7:0] t_r33_c47_4;
  wire [7:0] t_r33_c47_5;
  wire [7:0] t_r33_c47_6;
  wire [7:0] t_r33_c47_7;
  wire [7:0] t_r33_c47_8;
  wire [7:0] t_r33_c47_9;
  wire [7:0] t_r33_c47_10;
  wire [7:0] t_r33_c47_11;
  wire [7:0] t_r33_c47_12;
  wire [7:0] t_r33_c48_0;
  wire [7:0] t_r33_c48_1;
  wire [7:0] t_r33_c48_2;
  wire [7:0] t_r33_c48_3;
  wire [7:0] t_r33_c48_4;
  wire [7:0] t_r33_c48_5;
  wire [7:0] t_r33_c48_6;
  wire [7:0] t_r33_c48_7;
  wire [7:0] t_r33_c48_8;
  wire [7:0] t_r33_c48_9;
  wire [7:0] t_r33_c48_10;
  wire [7:0] t_r33_c48_11;
  wire [7:0] t_r33_c48_12;
  wire [7:0] t_r33_c49_0;
  wire [7:0] t_r33_c49_1;
  wire [7:0] t_r33_c49_2;
  wire [7:0] t_r33_c49_3;
  wire [7:0] t_r33_c49_4;
  wire [7:0] t_r33_c49_5;
  wire [7:0] t_r33_c49_6;
  wire [7:0] t_r33_c49_7;
  wire [7:0] t_r33_c49_8;
  wire [7:0] t_r33_c49_9;
  wire [7:0] t_r33_c49_10;
  wire [7:0] t_r33_c49_11;
  wire [7:0] t_r33_c49_12;
  wire [7:0] t_r33_c50_0;
  wire [7:0] t_r33_c50_1;
  wire [7:0] t_r33_c50_2;
  wire [7:0] t_r33_c50_3;
  wire [7:0] t_r33_c50_4;
  wire [7:0] t_r33_c50_5;
  wire [7:0] t_r33_c50_6;
  wire [7:0] t_r33_c50_7;
  wire [7:0] t_r33_c50_8;
  wire [7:0] t_r33_c50_9;
  wire [7:0] t_r33_c50_10;
  wire [7:0] t_r33_c50_11;
  wire [7:0] t_r33_c50_12;
  wire [7:0] t_r33_c51_0;
  wire [7:0] t_r33_c51_1;
  wire [7:0] t_r33_c51_2;
  wire [7:0] t_r33_c51_3;
  wire [7:0] t_r33_c51_4;
  wire [7:0] t_r33_c51_5;
  wire [7:0] t_r33_c51_6;
  wire [7:0] t_r33_c51_7;
  wire [7:0] t_r33_c51_8;
  wire [7:0] t_r33_c51_9;
  wire [7:0] t_r33_c51_10;
  wire [7:0] t_r33_c51_11;
  wire [7:0] t_r33_c51_12;
  wire [7:0] t_r33_c52_0;
  wire [7:0] t_r33_c52_1;
  wire [7:0] t_r33_c52_2;
  wire [7:0] t_r33_c52_3;
  wire [7:0] t_r33_c52_4;
  wire [7:0] t_r33_c52_5;
  wire [7:0] t_r33_c52_6;
  wire [7:0] t_r33_c52_7;
  wire [7:0] t_r33_c52_8;
  wire [7:0] t_r33_c52_9;
  wire [7:0] t_r33_c52_10;
  wire [7:0] t_r33_c52_11;
  wire [7:0] t_r33_c52_12;
  wire [7:0] t_r33_c53_0;
  wire [7:0] t_r33_c53_1;
  wire [7:0] t_r33_c53_2;
  wire [7:0] t_r33_c53_3;
  wire [7:0] t_r33_c53_4;
  wire [7:0] t_r33_c53_5;
  wire [7:0] t_r33_c53_6;
  wire [7:0] t_r33_c53_7;
  wire [7:0] t_r33_c53_8;
  wire [7:0] t_r33_c53_9;
  wire [7:0] t_r33_c53_10;
  wire [7:0] t_r33_c53_11;
  wire [7:0] t_r33_c53_12;
  wire [7:0] t_r33_c54_0;
  wire [7:0] t_r33_c54_1;
  wire [7:0] t_r33_c54_2;
  wire [7:0] t_r33_c54_3;
  wire [7:0] t_r33_c54_4;
  wire [7:0] t_r33_c54_5;
  wire [7:0] t_r33_c54_6;
  wire [7:0] t_r33_c54_7;
  wire [7:0] t_r33_c54_8;
  wire [7:0] t_r33_c54_9;
  wire [7:0] t_r33_c54_10;
  wire [7:0] t_r33_c54_11;
  wire [7:0] t_r33_c54_12;
  wire [7:0] t_r33_c55_0;
  wire [7:0] t_r33_c55_1;
  wire [7:0] t_r33_c55_2;
  wire [7:0] t_r33_c55_3;
  wire [7:0] t_r33_c55_4;
  wire [7:0] t_r33_c55_5;
  wire [7:0] t_r33_c55_6;
  wire [7:0] t_r33_c55_7;
  wire [7:0] t_r33_c55_8;
  wire [7:0] t_r33_c55_9;
  wire [7:0] t_r33_c55_10;
  wire [7:0] t_r33_c55_11;
  wire [7:0] t_r33_c55_12;
  wire [7:0] t_r33_c56_0;
  wire [7:0] t_r33_c56_1;
  wire [7:0] t_r33_c56_2;
  wire [7:0] t_r33_c56_3;
  wire [7:0] t_r33_c56_4;
  wire [7:0] t_r33_c56_5;
  wire [7:0] t_r33_c56_6;
  wire [7:0] t_r33_c56_7;
  wire [7:0] t_r33_c56_8;
  wire [7:0] t_r33_c56_9;
  wire [7:0] t_r33_c56_10;
  wire [7:0] t_r33_c56_11;
  wire [7:0] t_r33_c56_12;
  wire [7:0] t_r33_c57_0;
  wire [7:0] t_r33_c57_1;
  wire [7:0] t_r33_c57_2;
  wire [7:0] t_r33_c57_3;
  wire [7:0] t_r33_c57_4;
  wire [7:0] t_r33_c57_5;
  wire [7:0] t_r33_c57_6;
  wire [7:0] t_r33_c57_7;
  wire [7:0] t_r33_c57_8;
  wire [7:0] t_r33_c57_9;
  wire [7:0] t_r33_c57_10;
  wire [7:0] t_r33_c57_11;
  wire [7:0] t_r33_c57_12;
  wire [7:0] t_r33_c58_0;
  wire [7:0] t_r33_c58_1;
  wire [7:0] t_r33_c58_2;
  wire [7:0] t_r33_c58_3;
  wire [7:0] t_r33_c58_4;
  wire [7:0] t_r33_c58_5;
  wire [7:0] t_r33_c58_6;
  wire [7:0] t_r33_c58_7;
  wire [7:0] t_r33_c58_8;
  wire [7:0] t_r33_c58_9;
  wire [7:0] t_r33_c58_10;
  wire [7:0] t_r33_c58_11;
  wire [7:0] t_r33_c58_12;
  wire [7:0] t_r33_c59_0;
  wire [7:0] t_r33_c59_1;
  wire [7:0] t_r33_c59_2;
  wire [7:0] t_r33_c59_3;
  wire [7:0] t_r33_c59_4;
  wire [7:0] t_r33_c59_5;
  wire [7:0] t_r33_c59_6;
  wire [7:0] t_r33_c59_7;
  wire [7:0] t_r33_c59_8;
  wire [7:0] t_r33_c59_9;
  wire [7:0] t_r33_c59_10;
  wire [7:0] t_r33_c59_11;
  wire [7:0] t_r33_c59_12;
  wire [7:0] t_r33_c60_0;
  wire [7:0] t_r33_c60_1;
  wire [7:0] t_r33_c60_2;
  wire [7:0] t_r33_c60_3;
  wire [7:0] t_r33_c60_4;
  wire [7:0] t_r33_c60_5;
  wire [7:0] t_r33_c60_6;
  wire [7:0] t_r33_c60_7;
  wire [7:0] t_r33_c60_8;
  wire [7:0] t_r33_c60_9;
  wire [7:0] t_r33_c60_10;
  wire [7:0] t_r33_c60_11;
  wire [7:0] t_r33_c60_12;
  wire [7:0] t_r33_c61_0;
  wire [7:0] t_r33_c61_1;
  wire [7:0] t_r33_c61_2;
  wire [7:0] t_r33_c61_3;
  wire [7:0] t_r33_c61_4;
  wire [7:0] t_r33_c61_5;
  wire [7:0] t_r33_c61_6;
  wire [7:0] t_r33_c61_7;
  wire [7:0] t_r33_c61_8;
  wire [7:0] t_r33_c61_9;
  wire [7:0] t_r33_c61_10;
  wire [7:0] t_r33_c61_11;
  wire [7:0] t_r33_c61_12;
  wire [7:0] t_r33_c62_0;
  wire [7:0] t_r33_c62_1;
  wire [7:0] t_r33_c62_2;
  wire [7:0] t_r33_c62_3;
  wire [7:0] t_r33_c62_4;
  wire [7:0] t_r33_c62_5;
  wire [7:0] t_r33_c62_6;
  wire [7:0] t_r33_c62_7;
  wire [7:0] t_r33_c62_8;
  wire [7:0] t_r33_c62_9;
  wire [7:0] t_r33_c62_10;
  wire [7:0] t_r33_c62_11;
  wire [7:0] t_r33_c62_12;
  wire [7:0] t_r33_c63_0;
  wire [7:0] t_r33_c63_1;
  wire [7:0] t_r33_c63_2;
  wire [7:0] t_r33_c63_3;
  wire [7:0] t_r33_c63_4;
  wire [7:0] t_r33_c63_5;
  wire [7:0] t_r33_c63_6;
  wire [7:0] t_r33_c63_7;
  wire [7:0] t_r33_c63_8;
  wire [7:0] t_r33_c63_9;
  wire [7:0] t_r33_c63_10;
  wire [7:0] t_r33_c63_11;
  wire [7:0] t_r33_c63_12;
  wire [7:0] t_r33_c64_0;
  wire [7:0] t_r33_c64_1;
  wire [7:0] t_r33_c64_2;
  wire [7:0] t_r33_c64_3;
  wire [7:0] t_r33_c64_4;
  wire [7:0] t_r33_c64_5;
  wire [7:0] t_r33_c64_6;
  wire [7:0] t_r33_c64_7;
  wire [7:0] t_r33_c64_8;
  wire [7:0] t_r33_c64_9;
  wire [7:0] t_r33_c64_10;
  wire [7:0] t_r33_c64_11;
  wire [7:0] t_r33_c64_12;
  wire [7:0] t_r33_c65_0;
  wire [7:0] t_r33_c65_1;
  wire [7:0] t_r33_c65_2;
  wire [7:0] t_r33_c65_3;
  wire [7:0] t_r33_c65_4;
  wire [7:0] t_r33_c65_5;
  wire [7:0] t_r33_c65_6;
  wire [7:0] t_r33_c65_7;
  wire [7:0] t_r33_c65_8;
  wire [7:0] t_r33_c65_9;
  wire [7:0] t_r33_c65_10;
  wire [7:0] t_r33_c65_11;
  wire [7:0] t_r33_c65_12;
  wire [7:0] t_r34_c0_0;
  wire [7:0] t_r34_c0_1;
  wire [7:0] t_r34_c0_2;
  wire [7:0] t_r34_c0_3;
  wire [7:0] t_r34_c0_4;
  wire [7:0] t_r34_c0_5;
  wire [7:0] t_r34_c0_6;
  wire [7:0] t_r34_c0_7;
  wire [7:0] t_r34_c0_8;
  wire [7:0] t_r34_c0_9;
  wire [7:0] t_r34_c0_10;
  wire [7:0] t_r34_c0_11;
  wire [7:0] t_r34_c0_12;
  wire [7:0] t_r34_c1_0;
  wire [7:0] t_r34_c1_1;
  wire [7:0] t_r34_c1_2;
  wire [7:0] t_r34_c1_3;
  wire [7:0] t_r34_c1_4;
  wire [7:0] t_r34_c1_5;
  wire [7:0] t_r34_c1_6;
  wire [7:0] t_r34_c1_7;
  wire [7:0] t_r34_c1_8;
  wire [7:0] t_r34_c1_9;
  wire [7:0] t_r34_c1_10;
  wire [7:0] t_r34_c1_11;
  wire [7:0] t_r34_c1_12;
  wire [7:0] t_r34_c2_0;
  wire [7:0] t_r34_c2_1;
  wire [7:0] t_r34_c2_2;
  wire [7:0] t_r34_c2_3;
  wire [7:0] t_r34_c2_4;
  wire [7:0] t_r34_c2_5;
  wire [7:0] t_r34_c2_6;
  wire [7:0] t_r34_c2_7;
  wire [7:0] t_r34_c2_8;
  wire [7:0] t_r34_c2_9;
  wire [7:0] t_r34_c2_10;
  wire [7:0] t_r34_c2_11;
  wire [7:0] t_r34_c2_12;
  wire [7:0] t_r34_c3_0;
  wire [7:0] t_r34_c3_1;
  wire [7:0] t_r34_c3_2;
  wire [7:0] t_r34_c3_3;
  wire [7:0] t_r34_c3_4;
  wire [7:0] t_r34_c3_5;
  wire [7:0] t_r34_c3_6;
  wire [7:0] t_r34_c3_7;
  wire [7:0] t_r34_c3_8;
  wire [7:0] t_r34_c3_9;
  wire [7:0] t_r34_c3_10;
  wire [7:0] t_r34_c3_11;
  wire [7:0] t_r34_c3_12;
  wire [7:0] t_r34_c4_0;
  wire [7:0] t_r34_c4_1;
  wire [7:0] t_r34_c4_2;
  wire [7:0] t_r34_c4_3;
  wire [7:0] t_r34_c4_4;
  wire [7:0] t_r34_c4_5;
  wire [7:0] t_r34_c4_6;
  wire [7:0] t_r34_c4_7;
  wire [7:0] t_r34_c4_8;
  wire [7:0] t_r34_c4_9;
  wire [7:0] t_r34_c4_10;
  wire [7:0] t_r34_c4_11;
  wire [7:0] t_r34_c4_12;
  wire [7:0] t_r34_c5_0;
  wire [7:0] t_r34_c5_1;
  wire [7:0] t_r34_c5_2;
  wire [7:0] t_r34_c5_3;
  wire [7:0] t_r34_c5_4;
  wire [7:0] t_r34_c5_5;
  wire [7:0] t_r34_c5_6;
  wire [7:0] t_r34_c5_7;
  wire [7:0] t_r34_c5_8;
  wire [7:0] t_r34_c5_9;
  wire [7:0] t_r34_c5_10;
  wire [7:0] t_r34_c5_11;
  wire [7:0] t_r34_c5_12;
  wire [7:0] t_r34_c6_0;
  wire [7:0] t_r34_c6_1;
  wire [7:0] t_r34_c6_2;
  wire [7:0] t_r34_c6_3;
  wire [7:0] t_r34_c6_4;
  wire [7:0] t_r34_c6_5;
  wire [7:0] t_r34_c6_6;
  wire [7:0] t_r34_c6_7;
  wire [7:0] t_r34_c6_8;
  wire [7:0] t_r34_c6_9;
  wire [7:0] t_r34_c6_10;
  wire [7:0] t_r34_c6_11;
  wire [7:0] t_r34_c6_12;
  wire [7:0] t_r34_c7_0;
  wire [7:0] t_r34_c7_1;
  wire [7:0] t_r34_c7_2;
  wire [7:0] t_r34_c7_3;
  wire [7:0] t_r34_c7_4;
  wire [7:0] t_r34_c7_5;
  wire [7:0] t_r34_c7_6;
  wire [7:0] t_r34_c7_7;
  wire [7:0] t_r34_c7_8;
  wire [7:0] t_r34_c7_9;
  wire [7:0] t_r34_c7_10;
  wire [7:0] t_r34_c7_11;
  wire [7:0] t_r34_c7_12;
  wire [7:0] t_r34_c8_0;
  wire [7:0] t_r34_c8_1;
  wire [7:0] t_r34_c8_2;
  wire [7:0] t_r34_c8_3;
  wire [7:0] t_r34_c8_4;
  wire [7:0] t_r34_c8_5;
  wire [7:0] t_r34_c8_6;
  wire [7:0] t_r34_c8_7;
  wire [7:0] t_r34_c8_8;
  wire [7:0] t_r34_c8_9;
  wire [7:0] t_r34_c8_10;
  wire [7:0] t_r34_c8_11;
  wire [7:0] t_r34_c8_12;
  wire [7:0] t_r34_c9_0;
  wire [7:0] t_r34_c9_1;
  wire [7:0] t_r34_c9_2;
  wire [7:0] t_r34_c9_3;
  wire [7:0] t_r34_c9_4;
  wire [7:0] t_r34_c9_5;
  wire [7:0] t_r34_c9_6;
  wire [7:0] t_r34_c9_7;
  wire [7:0] t_r34_c9_8;
  wire [7:0] t_r34_c9_9;
  wire [7:0] t_r34_c9_10;
  wire [7:0] t_r34_c9_11;
  wire [7:0] t_r34_c9_12;
  wire [7:0] t_r34_c10_0;
  wire [7:0] t_r34_c10_1;
  wire [7:0] t_r34_c10_2;
  wire [7:0] t_r34_c10_3;
  wire [7:0] t_r34_c10_4;
  wire [7:0] t_r34_c10_5;
  wire [7:0] t_r34_c10_6;
  wire [7:0] t_r34_c10_7;
  wire [7:0] t_r34_c10_8;
  wire [7:0] t_r34_c10_9;
  wire [7:0] t_r34_c10_10;
  wire [7:0] t_r34_c10_11;
  wire [7:0] t_r34_c10_12;
  wire [7:0] t_r34_c11_0;
  wire [7:0] t_r34_c11_1;
  wire [7:0] t_r34_c11_2;
  wire [7:0] t_r34_c11_3;
  wire [7:0] t_r34_c11_4;
  wire [7:0] t_r34_c11_5;
  wire [7:0] t_r34_c11_6;
  wire [7:0] t_r34_c11_7;
  wire [7:0] t_r34_c11_8;
  wire [7:0] t_r34_c11_9;
  wire [7:0] t_r34_c11_10;
  wire [7:0] t_r34_c11_11;
  wire [7:0] t_r34_c11_12;
  wire [7:0] t_r34_c12_0;
  wire [7:0] t_r34_c12_1;
  wire [7:0] t_r34_c12_2;
  wire [7:0] t_r34_c12_3;
  wire [7:0] t_r34_c12_4;
  wire [7:0] t_r34_c12_5;
  wire [7:0] t_r34_c12_6;
  wire [7:0] t_r34_c12_7;
  wire [7:0] t_r34_c12_8;
  wire [7:0] t_r34_c12_9;
  wire [7:0] t_r34_c12_10;
  wire [7:0] t_r34_c12_11;
  wire [7:0] t_r34_c12_12;
  wire [7:0] t_r34_c13_0;
  wire [7:0] t_r34_c13_1;
  wire [7:0] t_r34_c13_2;
  wire [7:0] t_r34_c13_3;
  wire [7:0] t_r34_c13_4;
  wire [7:0] t_r34_c13_5;
  wire [7:0] t_r34_c13_6;
  wire [7:0] t_r34_c13_7;
  wire [7:0] t_r34_c13_8;
  wire [7:0] t_r34_c13_9;
  wire [7:0] t_r34_c13_10;
  wire [7:0] t_r34_c13_11;
  wire [7:0] t_r34_c13_12;
  wire [7:0] t_r34_c14_0;
  wire [7:0] t_r34_c14_1;
  wire [7:0] t_r34_c14_2;
  wire [7:0] t_r34_c14_3;
  wire [7:0] t_r34_c14_4;
  wire [7:0] t_r34_c14_5;
  wire [7:0] t_r34_c14_6;
  wire [7:0] t_r34_c14_7;
  wire [7:0] t_r34_c14_8;
  wire [7:0] t_r34_c14_9;
  wire [7:0] t_r34_c14_10;
  wire [7:0] t_r34_c14_11;
  wire [7:0] t_r34_c14_12;
  wire [7:0] t_r34_c15_0;
  wire [7:0] t_r34_c15_1;
  wire [7:0] t_r34_c15_2;
  wire [7:0] t_r34_c15_3;
  wire [7:0] t_r34_c15_4;
  wire [7:0] t_r34_c15_5;
  wire [7:0] t_r34_c15_6;
  wire [7:0] t_r34_c15_7;
  wire [7:0] t_r34_c15_8;
  wire [7:0] t_r34_c15_9;
  wire [7:0] t_r34_c15_10;
  wire [7:0] t_r34_c15_11;
  wire [7:0] t_r34_c15_12;
  wire [7:0] t_r34_c16_0;
  wire [7:0] t_r34_c16_1;
  wire [7:0] t_r34_c16_2;
  wire [7:0] t_r34_c16_3;
  wire [7:0] t_r34_c16_4;
  wire [7:0] t_r34_c16_5;
  wire [7:0] t_r34_c16_6;
  wire [7:0] t_r34_c16_7;
  wire [7:0] t_r34_c16_8;
  wire [7:0] t_r34_c16_9;
  wire [7:0] t_r34_c16_10;
  wire [7:0] t_r34_c16_11;
  wire [7:0] t_r34_c16_12;
  wire [7:0] t_r34_c17_0;
  wire [7:0] t_r34_c17_1;
  wire [7:0] t_r34_c17_2;
  wire [7:0] t_r34_c17_3;
  wire [7:0] t_r34_c17_4;
  wire [7:0] t_r34_c17_5;
  wire [7:0] t_r34_c17_6;
  wire [7:0] t_r34_c17_7;
  wire [7:0] t_r34_c17_8;
  wire [7:0] t_r34_c17_9;
  wire [7:0] t_r34_c17_10;
  wire [7:0] t_r34_c17_11;
  wire [7:0] t_r34_c17_12;
  wire [7:0] t_r34_c18_0;
  wire [7:0] t_r34_c18_1;
  wire [7:0] t_r34_c18_2;
  wire [7:0] t_r34_c18_3;
  wire [7:0] t_r34_c18_4;
  wire [7:0] t_r34_c18_5;
  wire [7:0] t_r34_c18_6;
  wire [7:0] t_r34_c18_7;
  wire [7:0] t_r34_c18_8;
  wire [7:0] t_r34_c18_9;
  wire [7:0] t_r34_c18_10;
  wire [7:0] t_r34_c18_11;
  wire [7:0] t_r34_c18_12;
  wire [7:0] t_r34_c19_0;
  wire [7:0] t_r34_c19_1;
  wire [7:0] t_r34_c19_2;
  wire [7:0] t_r34_c19_3;
  wire [7:0] t_r34_c19_4;
  wire [7:0] t_r34_c19_5;
  wire [7:0] t_r34_c19_6;
  wire [7:0] t_r34_c19_7;
  wire [7:0] t_r34_c19_8;
  wire [7:0] t_r34_c19_9;
  wire [7:0] t_r34_c19_10;
  wire [7:0] t_r34_c19_11;
  wire [7:0] t_r34_c19_12;
  wire [7:0] t_r34_c20_0;
  wire [7:0] t_r34_c20_1;
  wire [7:0] t_r34_c20_2;
  wire [7:0] t_r34_c20_3;
  wire [7:0] t_r34_c20_4;
  wire [7:0] t_r34_c20_5;
  wire [7:0] t_r34_c20_6;
  wire [7:0] t_r34_c20_7;
  wire [7:0] t_r34_c20_8;
  wire [7:0] t_r34_c20_9;
  wire [7:0] t_r34_c20_10;
  wire [7:0] t_r34_c20_11;
  wire [7:0] t_r34_c20_12;
  wire [7:0] t_r34_c21_0;
  wire [7:0] t_r34_c21_1;
  wire [7:0] t_r34_c21_2;
  wire [7:0] t_r34_c21_3;
  wire [7:0] t_r34_c21_4;
  wire [7:0] t_r34_c21_5;
  wire [7:0] t_r34_c21_6;
  wire [7:0] t_r34_c21_7;
  wire [7:0] t_r34_c21_8;
  wire [7:0] t_r34_c21_9;
  wire [7:0] t_r34_c21_10;
  wire [7:0] t_r34_c21_11;
  wire [7:0] t_r34_c21_12;
  wire [7:0] t_r34_c22_0;
  wire [7:0] t_r34_c22_1;
  wire [7:0] t_r34_c22_2;
  wire [7:0] t_r34_c22_3;
  wire [7:0] t_r34_c22_4;
  wire [7:0] t_r34_c22_5;
  wire [7:0] t_r34_c22_6;
  wire [7:0] t_r34_c22_7;
  wire [7:0] t_r34_c22_8;
  wire [7:0] t_r34_c22_9;
  wire [7:0] t_r34_c22_10;
  wire [7:0] t_r34_c22_11;
  wire [7:0] t_r34_c22_12;
  wire [7:0] t_r34_c23_0;
  wire [7:0] t_r34_c23_1;
  wire [7:0] t_r34_c23_2;
  wire [7:0] t_r34_c23_3;
  wire [7:0] t_r34_c23_4;
  wire [7:0] t_r34_c23_5;
  wire [7:0] t_r34_c23_6;
  wire [7:0] t_r34_c23_7;
  wire [7:0] t_r34_c23_8;
  wire [7:0] t_r34_c23_9;
  wire [7:0] t_r34_c23_10;
  wire [7:0] t_r34_c23_11;
  wire [7:0] t_r34_c23_12;
  wire [7:0] t_r34_c24_0;
  wire [7:0] t_r34_c24_1;
  wire [7:0] t_r34_c24_2;
  wire [7:0] t_r34_c24_3;
  wire [7:0] t_r34_c24_4;
  wire [7:0] t_r34_c24_5;
  wire [7:0] t_r34_c24_6;
  wire [7:0] t_r34_c24_7;
  wire [7:0] t_r34_c24_8;
  wire [7:0] t_r34_c24_9;
  wire [7:0] t_r34_c24_10;
  wire [7:0] t_r34_c24_11;
  wire [7:0] t_r34_c24_12;
  wire [7:0] t_r34_c25_0;
  wire [7:0] t_r34_c25_1;
  wire [7:0] t_r34_c25_2;
  wire [7:0] t_r34_c25_3;
  wire [7:0] t_r34_c25_4;
  wire [7:0] t_r34_c25_5;
  wire [7:0] t_r34_c25_6;
  wire [7:0] t_r34_c25_7;
  wire [7:0] t_r34_c25_8;
  wire [7:0] t_r34_c25_9;
  wire [7:0] t_r34_c25_10;
  wire [7:0] t_r34_c25_11;
  wire [7:0] t_r34_c25_12;
  wire [7:0] t_r34_c26_0;
  wire [7:0] t_r34_c26_1;
  wire [7:0] t_r34_c26_2;
  wire [7:0] t_r34_c26_3;
  wire [7:0] t_r34_c26_4;
  wire [7:0] t_r34_c26_5;
  wire [7:0] t_r34_c26_6;
  wire [7:0] t_r34_c26_7;
  wire [7:0] t_r34_c26_8;
  wire [7:0] t_r34_c26_9;
  wire [7:0] t_r34_c26_10;
  wire [7:0] t_r34_c26_11;
  wire [7:0] t_r34_c26_12;
  wire [7:0] t_r34_c27_0;
  wire [7:0] t_r34_c27_1;
  wire [7:0] t_r34_c27_2;
  wire [7:0] t_r34_c27_3;
  wire [7:0] t_r34_c27_4;
  wire [7:0] t_r34_c27_5;
  wire [7:0] t_r34_c27_6;
  wire [7:0] t_r34_c27_7;
  wire [7:0] t_r34_c27_8;
  wire [7:0] t_r34_c27_9;
  wire [7:0] t_r34_c27_10;
  wire [7:0] t_r34_c27_11;
  wire [7:0] t_r34_c27_12;
  wire [7:0] t_r34_c28_0;
  wire [7:0] t_r34_c28_1;
  wire [7:0] t_r34_c28_2;
  wire [7:0] t_r34_c28_3;
  wire [7:0] t_r34_c28_4;
  wire [7:0] t_r34_c28_5;
  wire [7:0] t_r34_c28_6;
  wire [7:0] t_r34_c28_7;
  wire [7:0] t_r34_c28_8;
  wire [7:0] t_r34_c28_9;
  wire [7:0] t_r34_c28_10;
  wire [7:0] t_r34_c28_11;
  wire [7:0] t_r34_c28_12;
  wire [7:0] t_r34_c29_0;
  wire [7:0] t_r34_c29_1;
  wire [7:0] t_r34_c29_2;
  wire [7:0] t_r34_c29_3;
  wire [7:0] t_r34_c29_4;
  wire [7:0] t_r34_c29_5;
  wire [7:0] t_r34_c29_6;
  wire [7:0] t_r34_c29_7;
  wire [7:0] t_r34_c29_8;
  wire [7:0] t_r34_c29_9;
  wire [7:0] t_r34_c29_10;
  wire [7:0] t_r34_c29_11;
  wire [7:0] t_r34_c29_12;
  wire [7:0] t_r34_c30_0;
  wire [7:0] t_r34_c30_1;
  wire [7:0] t_r34_c30_2;
  wire [7:0] t_r34_c30_3;
  wire [7:0] t_r34_c30_4;
  wire [7:0] t_r34_c30_5;
  wire [7:0] t_r34_c30_6;
  wire [7:0] t_r34_c30_7;
  wire [7:0] t_r34_c30_8;
  wire [7:0] t_r34_c30_9;
  wire [7:0] t_r34_c30_10;
  wire [7:0] t_r34_c30_11;
  wire [7:0] t_r34_c30_12;
  wire [7:0] t_r34_c31_0;
  wire [7:0] t_r34_c31_1;
  wire [7:0] t_r34_c31_2;
  wire [7:0] t_r34_c31_3;
  wire [7:0] t_r34_c31_4;
  wire [7:0] t_r34_c31_5;
  wire [7:0] t_r34_c31_6;
  wire [7:0] t_r34_c31_7;
  wire [7:0] t_r34_c31_8;
  wire [7:0] t_r34_c31_9;
  wire [7:0] t_r34_c31_10;
  wire [7:0] t_r34_c31_11;
  wire [7:0] t_r34_c31_12;
  wire [7:0] t_r34_c32_0;
  wire [7:0] t_r34_c32_1;
  wire [7:0] t_r34_c32_2;
  wire [7:0] t_r34_c32_3;
  wire [7:0] t_r34_c32_4;
  wire [7:0] t_r34_c32_5;
  wire [7:0] t_r34_c32_6;
  wire [7:0] t_r34_c32_7;
  wire [7:0] t_r34_c32_8;
  wire [7:0] t_r34_c32_9;
  wire [7:0] t_r34_c32_10;
  wire [7:0] t_r34_c32_11;
  wire [7:0] t_r34_c32_12;
  wire [7:0] t_r34_c33_0;
  wire [7:0] t_r34_c33_1;
  wire [7:0] t_r34_c33_2;
  wire [7:0] t_r34_c33_3;
  wire [7:0] t_r34_c33_4;
  wire [7:0] t_r34_c33_5;
  wire [7:0] t_r34_c33_6;
  wire [7:0] t_r34_c33_7;
  wire [7:0] t_r34_c33_8;
  wire [7:0] t_r34_c33_9;
  wire [7:0] t_r34_c33_10;
  wire [7:0] t_r34_c33_11;
  wire [7:0] t_r34_c33_12;
  wire [7:0] t_r34_c34_0;
  wire [7:0] t_r34_c34_1;
  wire [7:0] t_r34_c34_2;
  wire [7:0] t_r34_c34_3;
  wire [7:0] t_r34_c34_4;
  wire [7:0] t_r34_c34_5;
  wire [7:0] t_r34_c34_6;
  wire [7:0] t_r34_c34_7;
  wire [7:0] t_r34_c34_8;
  wire [7:0] t_r34_c34_9;
  wire [7:0] t_r34_c34_10;
  wire [7:0] t_r34_c34_11;
  wire [7:0] t_r34_c34_12;
  wire [7:0] t_r34_c35_0;
  wire [7:0] t_r34_c35_1;
  wire [7:0] t_r34_c35_2;
  wire [7:0] t_r34_c35_3;
  wire [7:0] t_r34_c35_4;
  wire [7:0] t_r34_c35_5;
  wire [7:0] t_r34_c35_6;
  wire [7:0] t_r34_c35_7;
  wire [7:0] t_r34_c35_8;
  wire [7:0] t_r34_c35_9;
  wire [7:0] t_r34_c35_10;
  wire [7:0] t_r34_c35_11;
  wire [7:0] t_r34_c35_12;
  wire [7:0] t_r34_c36_0;
  wire [7:0] t_r34_c36_1;
  wire [7:0] t_r34_c36_2;
  wire [7:0] t_r34_c36_3;
  wire [7:0] t_r34_c36_4;
  wire [7:0] t_r34_c36_5;
  wire [7:0] t_r34_c36_6;
  wire [7:0] t_r34_c36_7;
  wire [7:0] t_r34_c36_8;
  wire [7:0] t_r34_c36_9;
  wire [7:0] t_r34_c36_10;
  wire [7:0] t_r34_c36_11;
  wire [7:0] t_r34_c36_12;
  wire [7:0] t_r34_c37_0;
  wire [7:0] t_r34_c37_1;
  wire [7:0] t_r34_c37_2;
  wire [7:0] t_r34_c37_3;
  wire [7:0] t_r34_c37_4;
  wire [7:0] t_r34_c37_5;
  wire [7:0] t_r34_c37_6;
  wire [7:0] t_r34_c37_7;
  wire [7:0] t_r34_c37_8;
  wire [7:0] t_r34_c37_9;
  wire [7:0] t_r34_c37_10;
  wire [7:0] t_r34_c37_11;
  wire [7:0] t_r34_c37_12;
  wire [7:0] t_r34_c38_0;
  wire [7:0] t_r34_c38_1;
  wire [7:0] t_r34_c38_2;
  wire [7:0] t_r34_c38_3;
  wire [7:0] t_r34_c38_4;
  wire [7:0] t_r34_c38_5;
  wire [7:0] t_r34_c38_6;
  wire [7:0] t_r34_c38_7;
  wire [7:0] t_r34_c38_8;
  wire [7:0] t_r34_c38_9;
  wire [7:0] t_r34_c38_10;
  wire [7:0] t_r34_c38_11;
  wire [7:0] t_r34_c38_12;
  wire [7:0] t_r34_c39_0;
  wire [7:0] t_r34_c39_1;
  wire [7:0] t_r34_c39_2;
  wire [7:0] t_r34_c39_3;
  wire [7:0] t_r34_c39_4;
  wire [7:0] t_r34_c39_5;
  wire [7:0] t_r34_c39_6;
  wire [7:0] t_r34_c39_7;
  wire [7:0] t_r34_c39_8;
  wire [7:0] t_r34_c39_9;
  wire [7:0] t_r34_c39_10;
  wire [7:0] t_r34_c39_11;
  wire [7:0] t_r34_c39_12;
  wire [7:0] t_r34_c40_0;
  wire [7:0] t_r34_c40_1;
  wire [7:0] t_r34_c40_2;
  wire [7:0] t_r34_c40_3;
  wire [7:0] t_r34_c40_4;
  wire [7:0] t_r34_c40_5;
  wire [7:0] t_r34_c40_6;
  wire [7:0] t_r34_c40_7;
  wire [7:0] t_r34_c40_8;
  wire [7:0] t_r34_c40_9;
  wire [7:0] t_r34_c40_10;
  wire [7:0] t_r34_c40_11;
  wire [7:0] t_r34_c40_12;
  wire [7:0] t_r34_c41_0;
  wire [7:0] t_r34_c41_1;
  wire [7:0] t_r34_c41_2;
  wire [7:0] t_r34_c41_3;
  wire [7:0] t_r34_c41_4;
  wire [7:0] t_r34_c41_5;
  wire [7:0] t_r34_c41_6;
  wire [7:0] t_r34_c41_7;
  wire [7:0] t_r34_c41_8;
  wire [7:0] t_r34_c41_9;
  wire [7:0] t_r34_c41_10;
  wire [7:0] t_r34_c41_11;
  wire [7:0] t_r34_c41_12;
  wire [7:0] t_r34_c42_0;
  wire [7:0] t_r34_c42_1;
  wire [7:0] t_r34_c42_2;
  wire [7:0] t_r34_c42_3;
  wire [7:0] t_r34_c42_4;
  wire [7:0] t_r34_c42_5;
  wire [7:0] t_r34_c42_6;
  wire [7:0] t_r34_c42_7;
  wire [7:0] t_r34_c42_8;
  wire [7:0] t_r34_c42_9;
  wire [7:0] t_r34_c42_10;
  wire [7:0] t_r34_c42_11;
  wire [7:0] t_r34_c42_12;
  wire [7:0] t_r34_c43_0;
  wire [7:0] t_r34_c43_1;
  wire [7:0] t_r34_c43_2;
  wire [7:0] t_r34_c43_3;
  wire [7:0] t_r34_c43_4;
  wire [7:0] t_r34_c43_5;
  wire [7:0] t_r34_c43_6;
  wire [7:0] t_r34_c43_7;
  wire [7:0] t_r34_c43_8;
  wire [7:0] t_r34_c43_9;
  wire [7:0] t_r34_c43_10;
  wire [7:0] t_r34_c43_11;
  wire [7:0] t_r34_c43_12;
  wire [7:0] t_r34_c44_0;
  wire [7:0] t_r34_c44_1;
  wire [7:0] t_r34_c44_2;
  wire [7:0] t_r34_c44_3;
  wire [7:0] t_r34_c44_4;
  wire [7:0] t_r34_c44_5;
  wire [7:0] t_r34_c44_6;
  wire [7:0] t_r34_c44_7;
  wire [7:0] t_r34_c44_8;
  wire [7:0] t_r34_c44_9;
  wire [7:0] t_r34_c44_10;
  wire [7:0] t_r34_c44_11;
  wire [7:0] t_r34_c44_12;
  wire [7:0] t_r34_c45_0;
  wire [7:0] t_r34_c45_1;
  wire [7:0] t_r34_c45_2;
  wire [7:0] t_r34_c45_3;
  wire [7:0] t_r34_c45_4;
  wire [7:0] t_r34_c45_5;
  wire [7:0] t_r34_c45_6;
  wire [7:0] t_r34_c45_7;
  wire [7:0] t_r34_c45_8;
  wire [7:0] t_r34_c45_9;
  wire [7:0] t_r34_c45_10;
  wire [7:0] t_r34_c45_11;
  wire [7:0] t_r34_c45_12;
  wire [7:0] t_r34_c46_0;
  wire [7:0] t_r34_c46_1;
  wire [7:0] t_r34_c46_2;
  wire [7:0] t_r34_c46_3;
  wire [7:0] t_r34_c46_4;
  wire [7:0] t_r34_c46_5;
  wire [7:0] t_r34_c46_6;
  wire [7:0] t_r34_c46_7;
  wire [7:0] t_r34_c46_8;
  wire [7:0] t_r34_c46_9;
  wire [7:0] t_r34_c46_10;
  wire [7:0] t_r34_c46_11;
  wire [7:0] t_r34_c46_12;
  wire [7:0] t_r34_c47_0;
  wire [7:0] t_r34_c47_1;
  wire [7:0] t_r34_c47_2;
  wire [7:0] t_r34_c47_3;
  wire [7:0] t_r34_c47_4;
  wire [7:0] t_r34_c47_5;
  wire [7:0] t_r34_c47_6;
  wire [7:0] t_r34_c47_7;
  wire [7:0] t_r34_c47_8;
  wire [7:0] t_r34_c47_9;
  wire [7:0] t_r34_c47_10;
  wire [7:0] t_r34_c47_11;
  wire [7:0] t_r34_c47_12;
  wire [7:0] t_r34_c48_0;
  wire [7:0] t_r34_c48_1;
  wire [7:0] t_r34_c48_2;
  wire [7:0] t_r34_c48_3;
  wire [7:0] t_r34_c48_4;
  wire [7:0] t_r34_c48_5;
  wire [7:0] t_r34_c48_6;
  wire [7:0] t_r34_c48_7;
  wire [7:0] t_r34_c48_8;
  wire [7:0] t_r34_c48_9;
  wire [7:0] t_r34_c48_10;
  wire [7:0] t_r34_c48_11;
  wire [7:0] t_r34_c48_12;
  wire [7:0] t_r34_c49_0;
  wire [7:0] t_r34_c49_1;
  wire [7:0] t_r34_c49_2;
  wire [7:0] t_r34_c49_3;
  wire [7:0] t_r34_c49_4;
  wire [7:0] t_r34_c49_5;
  wire [7:0] t_r34_c49_6;
  wire [7:0] t_r34_c49_7;
  wire [7:0] t_r34_c49_8;
  wire [7:0] t_r34_c49_9;
  wire [7:0] t_r34_c49_10;
  wire [7:0] t_r34_c49_11;
  wire [7:0] t_r34_c49_12;
  wire [7:0] t_r34_c50_0;
  wire [7:0] t_r34_c50_1;
  wire [7:0] t_r34_c50_2;
  wire [7:0] t_r34_c50_3;
  wire [7:0] t_r34_c50_4;
  wire [7:0] t_r34_c50_5;
  wire [7:0] t_r34_c50_6;
  wire [7:0] t_r34_c50_7;
  wire [7:0] t_r34_c50_8;
  wire [7:0] t_r34_c50_9;
  wire [7:0] t_r34_c50_10;
  wire [7:0] t_r34_c50_11;
  wire [7:0] t_r34_c50_12;
  wire [7:0] t_r34_c51_0;
  wire [7:0] t_r34_c51_1;
  wire [7:0] t_r34_c51_2;
  wire [7:0] t_r34_c51_3;
  wire [7:0] t_r34_c51_4;
  wire [7:0] t_r34_c51_5;
  wire [7:0] t_r34_c51_6;
  wire [7:0] t_r34_c51_7;
  wire [7:0] t_r34_c51_8;
  wire [7:0] t_r34_c51_9;
  wire [7:0] t_r34_c51_10;
  wire [7:0] t_r34_c51_11;
  wire [7:0] t_r34_c51_12;
  wire [7:0] t_r34_c52_0;
  wire [7:0] t_r34_c52_1;
  wire [7:0] t_r34_c52_2;
  wire [7:0] t_r34_c52_3;
  wire [7:0] t_r34_c52_4;
  wire [7:0] t_r34_c52_5;
  wire [7:0] t_r34_c52_6;
  wire [7:0] t_r34_c52_7;
  wire [7:0] t_r34_c52_8;
  wire [7:0] t_r34_c52_9;
  wire [7:0] t_r34_c52_10;
  wire [7:0] t_r34_c52_11;
  wire [7:0] t_r34_c52_12;
  wire [7:0] t_r34_c53_0;
  wire [7:0] t_r34_c53_1;
  wire [7:0] t_r34_c53_2;
  wire [7:0] t_r34_c53_3;
  wire [7:0] t_r34_c53_4;
  wire [7:0] t_r34_c53_5;
  wire [7:0] t_r34_c53_6;
  wire [7:0] t_r34_c53_7;
  wire [7:0] t_r34_c53_8;
  wire [7:0] t_r34_c53_9;
  wire [7:0] t_r34_c53_10;
  wire [7:0] t_r34_c53_11;
  wire [7:0] t_r34_c53_12;
  wire [7:0] t_r34_c54_0;
  wire [7:0] t_r34_c54_1;
  wire [7:0] t_r34_c54_2;
  wire [7:0] t_r34_c54_3;
  wire [7:0] t_r34_c54_4;
  wire [7:0] t_r34_c54_5;
  wire [7:0] t_r34_c54_6;
  wire [7:0] t_r34_c54_7;
  wire [7:0] t_r34_c54_8;
  wire [7:0] t_r34_c54_9;
  wire [7:0] t_r34_c54_10;
  wire [7:0] t_r34_c54_11;
  wire [7:0] t_r34_c54_12;
  wire [7:0] t_r34_c55_0;
  wire [7:0] t_r34_c55_1;
  wire [7:0] t_r34_c55_2;
  wire [7:0] t_r34_c55_3;
  wire [7:0] t_r34_c55_4;
  wire [7:0] t_r34_c55_5;
  wire [7:0] t_r34_c55_6;
  wire [7:0] t_r34_c55_7;
  wire [7:0] t_r34_c55_8;
  wire [7:0] t_r34_c55_9;
  wire [7:0] t_r34_c55_10;
  wire [7:0] t_r34_c55_11;
  wire [7:0] t_r34_c55_12;
  wire [7:0] t_r34_c56_0;
  wire [7:0] t_r34_c56_1;
  wire [7:0] t_r34_c56_2;
  wire [7:0] t_r34_c56_3;
  wire [7:0] t_r34_c56_4;
  wire [7:0] t_r34_c56_5;
  wire [7:0] t_r34_c56_6;
  wire [7:0] t_r34_c56_7;
  wire [7:0] t_r34_c56_8;
  wire [7:0] t_r34_c56_9;
  wire [7:0] t_r34_c56_10;
  wire [7:0] t_r34_c56_11;
  wire [7:0] t_r34_c56_12;
  wire [7:0] t_r34_c57_0;
  wire [7:0] t_r34_c57_1;
  wire [7:0] t_r34_c57_2;
  wire [7:0] t_r34_c57_3;
  wire [7:0] t_r34_c57_4;
  wire [7:0] t_r34_c57_5;
  wire [7:0] t_r34_c57_6;
  wire [7:0] t_r34_c57_7;
  wire [7:0] t_r34_c57_8;
  wire [7:0] t_r34_c57_9;
  wire [7:0] t_r34_c57_10;
  wire [7:0] t_r34_c57_11;
  wire [7:0] t_r34_c57_12;
  wire [7:0] t_r34_c58_0;
  wire [7:0] t_r34_c58_1;
  wire [7:0] t_r34_c58_2;
  wire [7:0] t_r34_c58_3;
  wire [7:0] t_r34_c58_4;
  wire [7:0] t_r34_c58_5;
  wire [7:0] t_r34_c58_6;
  wire [7:0] t_r34_c58_7;
  wire [7:0] t_r34_c58_8;
  wire [7:0] t_r34_c58_9;
  wire [7:0] t_r34_c58_10;
  wire [7:0] t_r34_c58_11;
  wire [7:0] t_r34_c58_12;
  wire [7:0] t_r34_c59_0;
  wire [7:0] t_r34_c59_1;
  wire [7:0] t_r34_c59_2;
  wire [7:0] t_r34_c59_3;
  wire [7:0] t_r34_c59_4;
  wire [7:0] t_r34_c59_5;
  wire [7:0] t_r34_c59_6;
  wire [7:0] t_r34_c59_7;
  wire [7:0] t_r34_c59_8;
  wire [7:0] t_r34_c59_9;
  wire [7:0] t_r34_c59_10;
  wire [7:0] t_r34_c59_11;
  wire [7:0] t_r34_c59_12;
  wire [7:0] t_r34_c60_0;
  wire [7:0] t_r34_c60_1;
  wire [7:0] t_r34_c60_2;
  wire [7:0] t_r34_c60_3;
  wire [7:0] t_r34_c60_4;
  wire [7:0] t_r34_c60_5;
  wire [7:0] t_r34_c60_6;
  wire [7:0] t_r34_c60_7;
  wire [7:0] t_r34_c60_8;
  wire [7:0] t_r34_c60_9;
  wire [7:0] t_r34_c60_10;
  wire [7:0] t_r34_c60_11;
  wire [7:0] t_r34_c60_12;
  wire [7:0] t_r34_c61_0;
  wire [7:0] t_r34_c61_1;
  wire [7:0] t_r34_c61_2;
  wire [7:0] t_r34_c61_3;
  wire [7:0] t_r34_c61_4;
  wire [7:0] t_r34_c61_5;
  wire [7:0] t_r34_c61_6;
  wire [7:0] t_r34_c61_7;
  wire [7:0] t_r34_c61_8;
  wire [7:0] t_r34_c61_9;
  wire [7:0] t_r34_c61_10;
  wire [7:0] t_r34_c61_11;
  wire [7:0] t_r34_c61_12;
  wire [7:0] t_r34_c62_0;
  wire [7:0] t_r34_c62_1;
  wire [7:0] t_r34_c62_2;
  wire [7:0] t_r34_c62_3;
  wire [7:0] t_r34_c62_4;
  wire [7:0] t_r34_c62_5;
  wire [7:0] t_r34_c62_6;
  wire [7:0] t_r34_c62_7;
  wire [7:0] t_r34_c62_8;
  wire [7:0] t_r34_c62_9;
  wire [7:0] t_r34_c62_10;
  wire [7:0] t_r34_c62_11;
  wire [7:0] t_r34_c62_12;
  wire [7:0] t_r34_c63_0;
  wire [7:0] t_r34_c63_1;
  wire [7:0] t_r34_c63_2;
  wire [7:0] t_r34_c63_3;
  wire [7:0] t_r34_c63_4;
  wire [7:0] t_r34_c63_5;
  wire [7:0] t_r34_c63_6;
  wire [7:0] t_r34_c63_7;
  wire [7:0] t_r34_c63_8;
  wire [7:0] t_r34_c63_9;
  wire [7:0] t_r34_c63_10;
  wire [7:0] t_r34_c63_11;
  wire [7:0] t_r34_c63_12;
  wire [7:0] t_r34_c64_0;
  wire [7:0] t_r34_c64_1;
  wire [7:0] t_r34_c64_2;
  wire [7:0] t_r34_c64_3;
  wire [7:0] t_r34_c64_4;
  wire [7:0] t_r34_c64_5;
  wire [7:0] t_r34_c64_6;
  wire [7:0] t_r34_c64_7;
  wire [7:0] t_r34_c64_8;
  wire [7:0] t_r34_c64_9;
  wire [7:0] t_r34_c64_10;
  wire [7:0] t_r34_c64_11;
  wire [7:0] t_r34_c64_12;
  wire [7:0] t_r34_c65_0;
  wire [7:0] t_r34_c65_1;
  wire [7:0] t_r34_c65_2;
  wire [7:0] t_r34_c65_3;
  wire [7:0] t_r34_c65_4;
  wire [7:0] t_r34_c65_5;
  wire [7:0] t_r34_c65_6;
  wire [7:0] t_r34_c65_7;
  wire [7:0] t_r34_c65_8;
  wire [7:0] t_r34_c65_9;
  wire [7:0] t_r34_c65_10;
  wire [7:0] t_r34_c65_11;
  wire [7:0] t_r34_c65_12;
  wire [7:0] t_r35_c0_0;
  wire [7:0] t_r35_c0_1;
  wire [7:0] t_r35_c0_2;
  wire [7:0] t_r35_c0_3;
  wire [7:0] t_r35_c0_4;
  wire [7:0] t_r35_c0_5;
  wire [7:0] t_r35_c0_6;
  wire [7:0] t_r35_c0_7;
  wire [7:0] t_r35_c0_8;
  wire [7:0] t_r35_c0_9;
  wire [7:0] t_r35_c0_10;
  wire [7:0] t_r35_c0_11;
  wire [7:0] t_r35_c0_12;
  wire [7:0] t_r35_c1_0;
  wire [7:0] t_r35_c1_1;
  wire [7:0] t_r35_c1_2;
  wire [7:0] t_r35_c1_3;
  wire [7:0] t_r35_c1_4;
  wire [7:0] t_r35_c1_5;
  wire [7:0] t_r35_c1_6;
  wire [7:0] t_r35_c1_7;
  wire [7:0] t_r35_c1_8;
  wire [7:0] t_r35_c1_9;
  wire [7:0] t_r35_c1_10;
  wire [7:0] t_r35_c1_11;
  wire [7:0] t_r35_c1_12;
  wire [7:0] t_r35_c2_0;
  wire [7:0] t_r35_c2_1;
  wire [7:0] t_r35_c2_2;
  wire [7:0] t_r35_c2_3;
  wire [7:0] t_r35_c2_4;
  wire [7:0] t_r35_c2_5;
  wire [7:0] t_r35_c2_6;
  wire [7:0] t_r35_c2_7;
  wire [7:0] t_r35_c2_8;
  wire [7:0] t_r35_c2_9;
  wire [7:0] t_r35_c2_10;
  wire [7:0] t_r35_c2_11;
  wire [7:0] t_r35_c2_12;
  wire [7:0] t_r35_c3_0;
  wire [7:0] t_r35_c3_1;
  wire [7:0] t_r35_c3_2;
  wire [7:0] t_r35_c3_3;
  wire [7:0] t_r35_c3_4;
  wire [7:0] t_r35_c3_5;
  wire [7:0] t_r35_c3_6;
  wire [7:0] t_r35_c3_7;
  wire [7:0] t_r35_c3_8;
  wire [7:0] t_r35_c3_9;
  wire [7:0] t_r35_c3_10;
  wire [7:0] t_r35_c3_11;
  wire [7:0] t_r35_c3_12;
  wire [7:0] t_r35_c4_0;
  wire [7:0] t_r35_c4_1;
  wire [7:0] t_r35_c4_2;
  wire [7:0] t_r35_c4_3;
  wire [7:0] t_r35_c4_4;
  wire [7:0] t_r35_c4_5;
  wire [7:0] t_r35_c4_6;
  wire [7:0] t_r35_c4_7;
  wire [7:0] t_r35_c4_8;
  wire [7:0] t_r35_c4_9;
  wire [7:0] t_r35_c4_10;
  wire [7:0] t_r35_c4_11;
  wire [7:0] t_r35_c4_12;
  wire [7:0] t_r35_c5_0;
  wire [7:0] t_r35_c5_1;
  wire [7:0] t_r35_c5_2;
  wire [7:0] t_r35_c5_3;
  wire [7:0] t_r35_c5_4;
  wire [7:0] t_r35_c5_5;
  wire [7:0] t_r35_c5_6;
  wire [7:0] t_r35_c5_7;
  wire [7:0] t_r35_c5_8;
  wire [7:0] t_r35_c5_9;
  wire [7:0] t_r35_c5_10;
  wire [7:0] t_r35_c5_11;
  wire [7:0] t_r35_c5_12;
  wire [7:0] t_r35_c6_0;
  wire [7:0] t_r35_c6_1;
  wire [7:0] t_r35_c6_2;
  wire [7:0] t_r35_c6_3;
  wire [7:0] t_r35_c6_4;
  wire [7:0] t_r35_c6_5;
  wire [7:0] t_r35_c6_6;
  wire [7:0] t_r35_c6_7;
  wire [7:0] t_r35_c6_8;
  wire [7:0] t_r35_c6_9;
  wire [7:0] t_r35_c6_10;
  wire [7:0] t_r35_c6_11;
  wire [7:0] t_r35_c6_12;
  wire [7:0] t_r35_c7_0;
  wire [7:0] t_r35_c7_1;
  wire [7:0] t_r35_c7_2;
  wire [7:0] t_r35_c7_3;
  wire [7:0] t_r35_c7_4;
  wire [7:0] t_r35_c7_5;
  wire [7:0] t_r35_c7_6;
  wire [7:0] t_r35_c7_7;
  wire [7:0] t_r35_c7_8;
  wire [7:0] t_r35_c7_9;
  wire [7:0] t_r35_c7_10;
  wire [7:0] t_r35_c7_11;
  wire [7:0] t_r35_c7_12;
  wire [7:0] t_r35_c8_0;
  wire [7:0] t_r35_c8_1;
  wire [7:0] t_r35_c8_2;
  wire [7:0] t_r35_c8_3;
  wire [7:0] t_r35_c8_4;
  wire [7:0] t_r35_c8_5;
  wire [7:0] t_r35_c8_6;
  wire [7:0] t_r35_c8_7;
  wire [7:0] t_r35_c8_8;
  wire [7:0] t_r35_c8_9;
  wire [7:0] t_r35_c8_10;
  wire [7:0] t_r35_c8_11;
  wire [7:0] t_r35_c8_12;
  wire [7:0] t_r35_c9_0;
  wire [7:0] t_r35_c9_1;
  wire [7:0] t_r35_c9_2;
  wire [7:0] t_r35_c9_3;
  wire [7:0] t_r35_c9_4;
  wire [7:0] t_r35_c9_5;
  wire [7:0] t_r35_c9_6;
  wire [7:0] t_r35_c9_7;
  wire [7:0] t_r35_c9_8;
  wire [7:0] t_r35_c9_9;
  wire [7:0] t_r35_c9_10;
  wire [7:0] t_r35_c9_11;
  wire [7:0] t_r35_c9_12;
  wire [7:0] t_r35_c10_0;
  wire [7:0] t_r35_c10_1;
  wire [7:0] t_r35_c10_2;
  wire [7:0] t_r35_c10_3;
  wire [7:0] t_r35_c10_4;
  wire [7:0] t_r35_c10_5;
  wire [7:0] t_r35_c10_6;
  wire [7:0] t_r35_c10_7;
  wire [7:0] t_r35_c10_8;
  wire [7:0] t_r35_c10_9;
  wire [7:0] t_r35_c10_10;
  wire [7:0] t_r35_c10_11;
  wire [7:0] t_r35_c10_12;
  wire [7:0] t_r35_c11_0;
  wire [7:0] t_r35_c11_1;
  wire [7:0] t_r35_c11_2;
  wire [7:0] t_r35_c11_3;
  wire [7:0] t_r35_c11_4;
  wire [7:0] t_r35_c11_5;
  wire [7:0] t_r35_c11_6;
  wire [7:0] t_r35_c11_7;
  wire [7:0] t_r35_c11_8;
  wire [7:0] t_r35_c11_9;
  wire [7:0] t_r35_c11_10;
  wire [7:0] t_r35_c11_11;
  wire [7:0] t_r35_c11_12;
  wire [7:0] t_r35_c12_0;
  wire [7:0] t_r35_c12_1;
  wire [7:0] t_r35_c12_2;
  wire [7:0] t_r35_c12_3;
  wire [7:0] t_r35_c12_4;
  wire [7:0] t_r35_c12_5;
  wire [7:0] t_r35_c12_6;
  wire [7:0] t_r35_c12_7;
  wire [7:0] t_r35_c12_8;
  wire [7:0] t_r35_c12_9;
  wire [7:0] t_r35_c12_10;
  wire [7:0] t_r35_c12_11;
  wire [7:0] t_r35_c12_12;
  wire [7:0] t_r35_c13_0;
  wire [7:0] t_r35_c13_1;
  wire [7:0] t_r35_c13_2;
  wire [7:0] t_r35_c13_3;
  wire [7:0] t_r35_c13_4;
  wire [7:0] t_r35_c13_5;
  wire [7:0] t_r35_c13_6;
  wire [7:0] t_r35_c13_7;
  wire [7:0] t_r35_c13_8;
  wire [7:0] t_r35_c13_9;
  wire [7:0] t_r35_c13_10;
  wire [7:0] t_r35_c13_11;
  wire [7:0] t_r35_c13_12;
  wire [7:0] t_r35_c14_0;
  wire [7:0] t_r35_c14_1;
  wire [7:0] t_r35_c14_2;
  wire [7:0] t_r35_c14_3;
  wire [7:0] t_r35_c14_4;
  wire [7:0] t_r35_c14_5;
  wire [7:0] t_r35_c14_6;
  wire [7:0] t_r35_c14_7;
  wire [7:0] t_r35_c14_8;
  wire [7:0] t_r35_c14_9;
  wire [7:0] t_r35_c14_10;
  wire [7:0] t_r35_c14_11;
  wire [7:0] t_r35_c14_12;
  wire [7:0] t_r35_c15_0;
  wire [7:0] t_r35_c15_1;
  wire [7:0] t_r35_c15_2;
  wire [7:0] t_r35_c15_3;
  wire [7:0] t_r35_c15_4;
  wire [7:0] t_r35_c15_5;
  wire [7:0] t_r35_c15_6;
  wire [7:0] t_r35_c15_7;
  wire [7:0] t_r35_c15_8;
  wire [7:0] t_r35_c15_9;
  wire [7:0] t_r35_c15_10;
  wire [7:0] t_r35_c15_11;
  wire [7:0] t_r35_c15_12;
  wire [7:0] t_r35_c16_0;
  wire [7:0] t_r35_c16_1;
  wire [7:0] t_r35_c16_2;
  wire [7:0] t_r35_c16_3;
  wire [7:0] t_r35_c16_4;
  wire [7:0] t_r35_c16_5;
  wire [7:0] t_r35_c16_6;
  wire [7:0] t_r35_c16_7;
  wire [7:0] t_r35_c16_8;
  wire [7:0] t_r35_c16_9;
  wire [7:0] t_r35_c16_10;
  wire [7:0] t_r35_c16_11;
  wire [7:0] t_r35_c16_12;
  wire [7:0] t_r35_c17_0;
  wire [7:0] t_r35_c17_1;
  wire [7:0] t_r35_c17_2;
  wire [7:0] t_r35_c17_3;
  wire [7:0] t_r35_c17_4;
  wire [7:0] t_r35_c17_5;
  wire [7:0] t_r35_c17_6;
  wire [7:0] t_r35_c17_7;
  wire [7:0] t_r35_c17_8;
  wire [7:0] t_r35_c17_9;
  wire [7:0] t_r35_c17_10;
  wire [7:0] t_r35_c17_11;
  wire [7:0] t_r35_c17_12;
  wire [7:0] t_r35_c18_0;
  wire [7:0] t_r35_c18_1;
  wire [7:0] t_r35_c18_2;
  wire [7:0] t_r35_c18_3;
  wire [7:0] t_r35_c18_4;
  wire [7:0] t_r35_c18_5;
  wire [7:0] t_r35_c18_6;
  wire [7:0] t_r35_c18_7;
  wire [7:0] t_r35_c18_8;
  wire [7:0] t_r35_c18_9;
  wire [7:0] t_r35_c18_10;
  wire [7:0] t_r35_c18_11;
  wire [7:0] t_r35_c18_12;
  wire [7:0] t_r35_c19_0;
  wire [7:0] t_r35_c19_1;
  wire [7:0] t_r35_c19_2;
  wire [7:0] t_r35_c19_3;
  wire [7:0] t_r35_c19_4;
  wire [7:0] t_r35_c19_5;
  wire [7:0] t_r35_c19_6;
  wire [7:0] t_r35_c19_7;
  wire [7:0] t_r35_c19_8;
  wire [7:0] t_r35_c19_9;
  wire [7:0] t_r35_c19_10;
  wire [7:0] t_r35_c19_11;
  wire [7:0] t_r35_c19_12;
  wire [7:0] t_r35_c20_0;
  wire [7:0] t_r35_c20_1;
  wire [7:0] t_r35_c20_2;
  wire [7:0] t_r35_c20_3;
  wire [7:0] t_r35_c20_4;
  wire [7:0] t_r35_c20_5;
  wire [7:0] t_r35_c20_6;
  wire [7:0] t_r35_c20_7;
  wire [7:0] t_r35_c20_8;
  wire [7:0] t_r35_c20_9;
  wire [7:0] t_r35_c20_10;
  wire [7:0] t_r35_c20_11;
  wire [7:0] t_r35_c20_12;
  wire [7:0] t_r35_c21_0;
  wire [7:0] t_r35_c21_1;
  wire [7:0] t_r35_c21_2;
  wire [7:0] t_r35_c21_3;
  wire [7:0] t_r35_c21_4;
  wire [7:0] t_r35_c21_5;
  wire [7:0] t_r35_c21_6;
  wire [7:0] t_r35_c21_7;
  wire [7:0] t_r35_c21_8;
  wire [7:0] t_r35_c21_9;
  wire [7:0] t_r35_c21_10;
  wire [7:0] t_r35_c21_11;
  wire [7:0] t_r35_c21_12;
  wire [7:0] t_r35_c22_0;
  wire [7:0] t_r35_c22_1;
  wire [7:0] t_r35_c22_2;
  wire [7:0] t_r35_c22_3;
  wire [7:0] t_r35_c22_4;
  wire [7:0] t_r35_c22_5;
  wire [7:0] t_r35_c22_6;
  wire [7:0] t_r35_c22_7;
  wire [7:0] t_r35_c22_8;
  wire [7:0] t_r35_c22_9;
  wire [7:0] t_r35_c22_10;
  wire [7:0] t_r35_c22_11;
  wire [7:0] t_r35_c22_12;
  wire [7:0] t_r35_c23_0;
  wire [7:0] t_r35_c23_1;
  wire [7:0] t_r35_c23_2;
  wire [7:0] t_r35_c23_3;
  wire [7:0] t_r35_c23_4;
  wire [7:0] t_r35_c23_5;
  wire [7:0] t_r35_c23_6;
  wire [7:0] t_r35_c23_7;
  wire [7:0] t_r35_c23_8;
  wire [7:0] t_r35_c23_9;
  wire [7:0] t_r35_c23_10;
  wire [7:0] t_r35_c23_11;
  wire [7:0] t_r35_c23_12;
  wire [7:0] t_r35_c24_0;
  wire [7:0] t_r35_c24_1;
  wire [7:0] t_r35_c24_2;
  wire [7:0] t_r35_c24_3;
  wire [7:0] t_r35_c24_4;
  wire [7:0] t_r35_c24_5;
  wire [7:0] t_r35_c24_6;
  wire [7:0] t_r35_c24_7;
  wire [7:0] t_r35_c24_8;
  wire [7:0] t_r35_c24_9;
  wire [7:0] t_r35_c24_10;
  wire [7:0] t_r35_c24_11;
  wire [7:0] t_r35_c24_12;
  wire [7:0] t_r35_c25_0;
  wire [7:0] t_r35_c25_1;
  wire [7:0] t_r35_c25_2;
  wire [7:0] t_r35_c25_3;
  wire [7:0] t_r35_c25_4;
  wire [7:0] t_r35_c25_5;
  wire [7:0] t_r35_c25_6;
  wire [7:0] t_r35_c25_7;
  wire [7:0] t_r35_c25_8;
  wire [7:0] t_r35_c25_9;
  wire [7:0] t_r35_c25_10;
  wire [7:0] t_r35_c25_11;
  wire [7:0] t_r35_c25_12;
  wire [7:0] t_r35_c26_0;
  wire [7:0] t_r35_c26_1;
  wire [7:0] t_r35_c26_2;
  wire [7:0] t_r35_c26_3;
  wire [7:0] t_r35_c26_4;
  wire [7:0] t_r35_c26_5;
  wire [7:0] t_r35_c26_6;
  wire [7:0] t_r35_c26_7;
  wire [7:0] t_r35_c26_8;
  wire [7:0] t_r35_c26_9;
  wire [7:0] t_r35_c26_10;
  wire [7:0] t_r35_c26_11;
  wire [7:0] t_r35_c26_12;
  wire [7:0] t_r35_c27_0;
  wire [7:0] t_r35_c27_1;
  wire [7:0] t_r35_c27_2;
  wire [7:0] t_r35_c27_3;
  wire [7:0] t_r35_c27_4;
  wire [7:0] t_r35_c27_5;
  wire [7:0] t_r35_c27_6;
  wire [7:0] t_r35_c27_7;
  wire [7:0] t_r35_c27_8;
  wire [7:0] t_r35_c27_9;
  wire [7:0] t_r35_c27_10;
  wire [7:0] t_r35_c27_11;
  wire [7:0] t_r35_c27_12;
  wire [7:0] t_r35_c28_0;
  wire [7:0] t_r35_c28_1;
  wire [7:0] t_r35_c28_2;
  wire [7:0] t_r35_c28_3;
  wire [7:0] t_r35_c28_4;
  wire [7:0] t_r35_c28_5;
  wire [7:0] t_r35_c28_6;
  wire [7:0] t_r35_c28_7;
  wire [7:0] t_r35_c28_8;
  wire [7:0] t_r35_c28_9;
  wire [7:0] t_r35_c28_10;
  wire [7:0] t_r35_c28_11;
  wire [7:0] t_r35_c28_12;
  wire [7:0] t_r35_c29_0;
  wire [7:0] t_r35_c29_1;
  wire [7:0] t_r35_c29_2;
  wire [7:0] t_r35_c29_3;
  wire [7:0] t_r35_c29_4;
  wire [7:0] t_r35_c29_5;
  wire [7:0] t_r35_c29_6;
  wire [7:0] t_r35_c29_7;
  wire [7:0] t_r35_c29_8;
  wire [7:0] t_r35_c29_9;
  wire [7:0] t_r35_c29_10;
  wire [7:0] t_r35_c29_11;
  wire [7:0] t_r35_c29_12;
  wire [7:0] t_r35_c30_0;
  wire [7:0] t_r35_c30_1;
  wire [7:0] t_r35_c30_2;
  wire [7:0] t_r35_c30_3;
  wire [7:0] t_r35_c30_4;
  wire [7:0] t_r35_c30_5;
  wire [7:0] t_r35_c30_6;
  wire [7:0] t_r35_c30_7;
  wire [7:0] t_r35_c30_8;
  wire [7:0] t_r35_c30_9;
  wire [7:0] t_r35_c30_10;
  wire [7:0] t_r35_c30_11;
  wire [7:0] t_r35_c30_12;
  wire [7:0] t_r35_c31_0;
  wire [7:0] t_r35_c31_1;
  wire [7:0] t_r35_c31_2;
  wire [7:0] t_r35_c31_3;
  wire [7:0] t_r35_c31_4;
  wire [7:0] t_r35_c31_5;
  wire [7:0] t_r35_c31_6;
  wire [7:0] t_r35_c31_7;
  wire [7:0] t_r35_c31_8;
  wire [7:0] t_r35_c31_9;
  wire [7:0] t_r35_c31_10;
  wire [7:0] t_r35_c31_11;
  wire [7:0] t_r35_c31_12;
  wire [7:0] t_r35_c32_0;
  wire [7:0] t_r35_c32_1;
  wire [7:0] t_r35_c32_2;
  wire [7:0] t_r35_c32_3;
  wire [7:0] t_r35_c32_4;
  wire [7:0] t_r35_c32_5;
  wire [7:0] t_r35_c32_6;
  wire [7:0] t_r35_c32_7;
  wire [7:0] t_r35_c32_8;
  wire [7:0] t_r35_c32_9;
  wire [7:0] t_r35_c32_10;
  wire [7:0] t_r35_c32_11;
  wire [7:0] t_r35_c32_12;
  wire [7:0] t_r35_c33_0;
  wire [7:0] t_r35_c33_1;
  wire [7:0] t_r35_c33_2;
  wire [7:0] t_r35_c33_3;
  wire [7:0] t_r35_c33_4;
  wire [7:0] t_r35_c33_5;
  wire [7:0] t_r35_c33_6;
  wire [7:0] t_r35_c33_7;
  wire [7:0] t_r35_c33_8;
  wire [7:0] t_r35_c33_9;
  wire [7:0] t_r35_c33_10;
  wire [7:0] t_r35_c33_11;
  wire [7:0] t_r35_c33_12;
  wire [7:0] t_r35_c34_0;
  wire [7:0] t_r35_c34_1;
  wire [7:0] t_r35_c34_2;
  wire [7:0] t_r35_c34_3;
  wire [7:0] t_r35_c34_4;
  wire [7:0] t_r35_c34_5;
  wire [7:0] t_r35_c34_6;
  wire [7:0] t_r35_c34_7;
  wire [7:0] t_r35_c34_8;
  wire [7:0] t_r35_c34_9;
  wire [7:0] t_r35_c34_10;
  wire [7:0] t_r35_c34_11;
  wire [7:0] t_r35_c34_12;
  wire [7:0] t_r35_c35_0;
  wire [7:0] t_r35_c35_1;
  wire [7:0] t_r35_c35_2;
  wire [7:0] t_r35_c35_3;
  wire [7:0] t_r35_c35_4;
  wire [7:0] t_r35_c35_5;
  wire [7:0] t_r35_c35_6;
  wire [7:0] t_r35_c35_7;
  wire [7:0] t_r35_c35_8;
  wire [7:0] t_r35_c35_9;
  wire [7:0] t_r35_c35_10;
  wire [7:0] t_r35_c35_11;
  wire [7:0] t_r35_c35_12;
  wire [7:0] t_r35_c36_0;
  wire [7:0] t_r35_c36_1;
  wire [7:0] t_r35_c36_2;
  wire [7:0] t_r35_c36_3;
  wire [7:0] t_r35_c36_4;
  wire [7:0] t_r35_c36_5;
  wire [7:0] t_r35_c36_6;
  wire [7:0] t_r35_c36_7;
  wire [7:0] t_r35_c36_8;
  wire [7:0] t_r35_c36_9;
  wire [7:0] t_r35_c36_10;
  wire [7:0] t_r35_c36_11;
  wire [7:0] t_r35_c36_12;
  wire [7:0] t_r35_c37_0;
  wire [7:0] t_r35_c37_1;
  wire [7:0] t_r35_c37_2;
  wire [7:0] t_r35_c37_3;
  wire [7:0] t_r35_c37_4;
  wire [7:0] t_r35_c37_5;
  wire [7:0] t_r35_c37_6;
  wire [7:0] t_r35_c37_7;
  wire [7:0] t_r35_c37_8;
  wire [7:0] t_r35_c37_9;
  wire [7:0] t_r35_c37_10;
  wire [7:0] t_r35_c37_11;
  wire [7:0] t_r35_c37_12;
  wire [7:0] t_r35_c38_0;
  wire [7:0] t_r35_c38_1;
  wire [7:0] t_r35_c38_2;
  wire [7:0] t_r35_c38_3;
  wire [7:0] t_r35_c38_4;
  wire [7:0] t_r35_c38_5;
  wire [7:0] t_r35_c38_6;
  wire [7:0] t_r35_c38_7;
  wire [7:0] t_r35_c38_8;
  wire [7:0] t_r35_c38_9;
  wire [7:0] t_r35_c38_10;
  wire [7:0] t_r35_c38_11;
  wire [7:0] t_r35_c38_12;
  wire [7:0] t_r35_c39_0;
  wire [7:0] t_r35_c39_1;
  wire [7:0] t_r35_c39_2;
  wire [7:0] t_r35_c39_3;
  wire [7:0] t_r35_c39_4;
  wire [7:0] t_r35_c39_5;
  wire [7:0] t_r35_c39_6;
  wire [7:0] t_r35_c39_7;
  wire [7:0] t_r35_c39_8;
  wire [7:0] t_r35_c39_9;
  wire [7:0] t_r35_c39_10;
  wire [7:0] t_r35_c39_11;
  wire [7:0] t_r35_c39_12;
  wire [7:0] t_r35_c40_0;
  wire [7:0] t_r35_c40_1;
  wire [7:0] t_r35_c40_2;
  wire [7:0] t_r35_c40_3;
  wire [7:0] t_r35_c40_4;
  wire [7:0] t_r35_c40_5;
  wire [7:0] t_r35_c40_6;
  wire [7:0] t_r35_c40_7;
  wire [7:0] t_r35_c40_8;
  wire [7:0] t_r35_c40_9;
  wire [7:0] t_r35_c40_10;
  wire [7:0] t_r35_c40_11;
  wire [7:0] t_r35_c40_12;
  wire [7:0] t_r35_c41_0;
  wire [7:0] t_r35_c41_1;
  wire [7:0] t_r35_c41_2;
  wire [7:0] t_r35_c41_3;
  wire [7:0] t_r35_c41_4;
  wire [7:0] t_r35_c41_5;
  wire [7:0] t_r35_c41_6;
  wire [7:0] t_r35_c41_7;
  wire [7:0] t_r35_c41_8;
  wire [7:0] t_r35_c41_9;
  wire [7:0] t_r35_c41_10;
  wire [7:0] t_r35_c41_11;
  wire [7:0] t_r35_c41_12;
  wire [7:0] t_r35_c42_0;
  wire [7:0] t_r35_c42_1;
  wire [7:0] t_r35_c42_2;
  wire [7:0] t_r35_c42_3;
  wire [7:0] t_r35_c42_4;
  wire [7:0] t_r35_c42_5;
  wire [7:0] t_r35_c42_6;
  wire [7:0] t_r35_c42_7;
  wire [7:0] t_r35_c42_8;
  wire [7:0] t_r35_c42_9;
  wire [7:0] t_r35_c42_10;
  wire [7:0] t_r35_c42_11;
  wire [7:0] t_r35_c42_12;
  wire [7:0] t_r35_c43_0;
  wire [7:0] t_r35_c43_1;
  wire [7:0] t_r35_c43_2;
  wire [7:0] t_r35_c43_3;
  wire [7:0] t_r35_c43_4;
  wire [7:0] t_r35_c43_5;
  wire [7:0] t_r35_c43_6;
  wire [7:0] t_r35_c43_7;
  wire [7:0] t_r35_c43_8;
  wire [7:0] t_r35_c43_9;
  wire [7:0] t_r35_c43_10;
  wire [7:0] t_r35_c43_11;
  wire [7:0] t_r35_c43_12;
  wire [7:0] t_r35_c44_0;
  wire [7:0] t_r35_c44_1;
  wire [7:0] t_r35_c44_2;
  wire [7:0] t_r35_c44_3;
  wire [7:0] t_r35_c44_4;
  wire [7:0] t_r35_c44_5;
  wire [7:0] t_r35_c44_6;
  wire [7:0] t_r35_c44_7;
  wire [7:0] t_r35_c44_8;
  wire [7:0] t_r35_c44_9;
  wire [7:0] t_r35_c44_10;
  wire [7:0] t_r35_c44_11;
  wire [7:0] t_r35_c44_12;
  wire [7:0] t_r35_c45_0;
  wire [7:0] t_r35_c45_1;
  wire [7:0] t_r35_c45_2;
  wire [7:0] t_r35_c45_3;
  wire [7:0] t_r35_c45_4;
  wire [7:0] t_r35_c45_5;
  wire [7:0] t_r35_c45_6;
  wire [7:0] t_r35_c45_7;
  wire [7:0] t_r35_c45_8;
  wire [7:0] t_r35_c45_9;
  wire [7:0] t_r35_c45_10;
  wire [7:0] t_r35_c45_11;
  wire [7:0] t_r35_c45_12;
  wire [7:0] t_r35_c46_0;
  wire [7:0] t_r35_c46_1;
  wire [7:0] t_r35_c46_2;
  wire [7:0] t_r35_c46_3;
  wire [7:0] t_r35_c46_4;
  wire [7:0] t_r35_c46_5;
  wire [7:0] t_r35_c46_6;
  wire [7:0] t_r35_c46_7;
  wire [7:0] t_r35_c46_8;
  wire [7:0] t_r35_c46_9;
  wire [7:0] t_r35_c46_10;
  wire [7:0] t_r35_c46_11;
  wire [7:0] t_r35_c46_12;
  wire [7:0] t_r35_c47_0;
  wire [7:0] t_r35_c47_1;
  wire [7:0] t_r35_c47_2;
  wire [7:0] t_r35_c47_3;
  wire [7:0] t_r35_c47_4;
  wire [7:0] t_r35_c47_5;
  wire [7:0] t_r35_c47_6;
  wire [7:0] t_r35_c47_7;
  wire [7:0] t_r35_c47_8;
  wire [7:0] t_r35_c47_9;
  wire [7:0] t_r35_c47_10;
  wire [7:0] t_r35_c47_11;
  wire [7:0] t_r35_c47_12;
  wire [7:0] t_r35_c48_0;
  wire [7:0] t_r35_c48_1;
  wire [7:0] t_r35_c48_2;
  wire [7:0] t_r35_c48_3;
  wire [7:0] t_r35_c48_4;
  wire [7:0] t_r35_c48_5;
  wire [7:0] t_r35_c48_6;
  wire [7:0] t_r35_c48_7;
  wire [7:0] t_r35_c48_8;
  wire [7:0] t_r35_c48_9;
  wire [7:0] t_r35_c48_10;
  wire [7:0] t_r35_c48_11;
  wire [7:0] t_r35_c48_12;
  wire [7:0] t_r35_c49_0;
  wire [7:0] t_r35_c49_1;
  wire [7:0] t_r35_c49_2;
  wire [7:0] t_r35_c49_3;
  wire [7:0] t_r35_c49_4;
  wire [7:0] t_r35_c49_5;
  wire [7:0] t_r35_c49_6;
  wire [7:0] t_r35_c49_7;
  wire [7:0] t_r35_c49_8;
  wire [7:0] t_r35_c49_9;
  wire [7:0] t_r35_c49_10;
  wire [7:0] t_r35_c49_11;
  wire [7:0] t_r35_c49_12;
  wire [7:0] t_r35_c50_0;
  wire [7:0] t_r35_c50_1;
  wire [7:0] t_r35_c50_2;
  wire [7:0] t_r35_c50_3;
  wire [7:0] t_r35_c50_4;
  wire [7:0] t_r35_c50_5;
  wire [7:0] t_r35_c50_6;
  wire [7:0] t_r35_c50_7;
  wire [7:0] t_r35_c50_8;
  wire [7:0] t_r35_c50_9;
  wire [7:0] t_r35_c50_10;
  wire [7:0] t_r35_c50_11;
  wire [7:0] t_r35_c50_12;
  wire [7:0] t_r35_c51_0;
  wire [7:0] t_r35_c51_1;
  wire [7:0] t_r35_c51_2;
  wire [7:0] t_r35_c51_3;
  wire [7:0] t_r35_c51_4;
  wire [7:0] t_r35_c51_5;
  wire [7:0] t_r35_c51_6;
  wire [7:0] t_r35_c51_7;
  wire [7:0] t_r35_c51_8;
  wire [7:0] t_r35_c51_9;
  wire [7:0] t_r35_c51_10;
  wire [7:0] t_r35_c51_11;
  wire [7:0] t_r35_c51_12;
  wire [7:0] t_r35_c52_0;
  wire [7:0] t_r35_c52_1;
  wire [7:0] t_r35_c52_2;
  wire [7:0] t_r35_c52_3;
  wire [7:0] t_r35_c52_4;
  wire [7:0] t_r35_c52_5;
  wire [7:0] t_r35_c52_6;
  wire [7:0] t_r35_c52_7;
  wire [7:0] t_r35_c52_8;
  wire [7:0] t_r35_c52_9;
  wire [7:0] t_r35_c52_10;
  wire [7:0] t_r35_c52_11;
  wire [7:0] t_r35_c52_12;
  wire [7:0] t_r35_c53_0;
  wire [7:0] t_r35_c53_1;
  wire [7:0] t_r35_c53_2;
  wire [7:0] t_r35_c53_3;
  wire [7:0] t_r35_c53_4;
  wire [7:0] t_r35_c53_5;
  wire [7:0] t_r35_c53_6;
  wire [7:0] t_r35_c53_7;
  wire [7:0] t_r35_c53_8;
  wire [7:0] t_r35_c53_9;
  wire [7:0] t_r35_c53_10;
  wire [7:0] t_r35_c53_11;
  wire [7:0] t_r35_c53_12;
  wire [7:0] t_r35_c54_0;
  wire [7:0] t_r35_c54_1;
  wire [7:0] t_r35_c54_2;
  wire [7:0] t_r35_c54_3;
  wire [7:0] t_r35_c54_4;
  wire [7:0] t_r35_c54_5;
  wire [7:0] t_r35_c54_6;
  wire [7:0] t_r35_c54_7;
  wire [7:0] t_r35_c54_8;
  wire [7:0] t_r35_c54_9;
  wire [7:0] t_r35_c54_10;
  wire [7:0] t_r35_c54_11;
  wire [7:0] t_r35_c54_12;
  wire [7:0] t_r35_c55_0;
  wire [7:0] t_r35_c55_1;
  wire [7:0] t_r35_c55_2;
  wire [7:0] t_r35_c55_3;
  wire [7:0] t_r35_c55_4;
  wire [7:0] t_r35_c55_5;
  wire [7:0] t_r35_c55_6;
  wire [7:0] t_r35_c55_7;
  wire [7:0] t_r35_c55_8;
  wire [7:0] t_r35_c55_9;
  wire [7:0] t_r35_c55_10;
  wire [7:0] t_r35_c55_11;
  wire [7:0] t_r35_c55_12;
  wire [7:0] t_r35_c56_0;
  wire [7:0] t_r35_c56_1;
  wire [7:0] t_r35_c56_2;
  wire [7:0] t_r35_c56_3;
  wire [7:0] t_r35_c56_4;
  wire [7:0] t_r35_c56_5;
  wire [7:0] t_r35_c56_6;
  wire [7:0] t_r35_c56_7;
  wire [7:0] t_r35_c56_8;
  wire [7:0] t_r35_c56_9;
  wire [7:0] t_r35_c56_10;
  wire [7:0] t_r35_c56_11;
  wire [7:0] t_r35_c56_12;
  wire [7:0] t_r35_c57_0;
  wire [7:0] t_r35_c57_1;
  wire [7:0] t_r35_c57_2;
  wire [7:0] t_r35_c57_3;
  wire [7:0] t_r35_c57_4;
  wire [7:0] t_r35_c57_5;
  wire [7:0] t_r35_c57_6;
  wire [7:0] t_r35_c57_7;
  wire [7:0] t_r35_c57_8;
  wire [7:0] t_r35_c57_9;
  wire [7:0] t_r35_c57_10;
  wire [7:0] t_r35_c57_11;
  wire [7:0] t_r35_c57_12;
  wire [7:0] t_r35_c58_0;
  wire [7:0] t_r35_c58_1;
  wire [7:0] t_r35_c58_2;
  wire [7:0] t_r35_c58_3;
  wire [7:0] t_r35_c58_4;
  wire [7:0] t_r35_c58_5;
  wire [7:0] t_r35_c58_6;
  wire [7:0] t_r35_c58_7;
  wire [7:0] t_r35_c58_8;
  wire [7:0] t_r35_c58_9;
  wire [7:0] t_r35_c58_10;
  wire [7:0] t_r35_c58_11;
  wire [7:0] t_r35_c58_12;
  wire [7:0] t_r35_c59_0;
  wire [7:0] t_r35_c59_1;
  wire [7:0] t_r35_c59_2;
  wire [7:0] t_r35_c59_3;
  wire [7:0] t_r35_c59_4;
  wire [7:0] t_r35_c59_5;
  wire [7:0] t_r35_c59_6;
  wire [7:0] t_r35_c59_7;
  wire [7:0] t_r35_c59_8;
  wire [7:0] t_r35_c59_9;
  wire [7:0] t_r35_c59_10;
  wire [7:0] t_r35_c59_11;
  wire [7:0] t_r35_c59_12;
  wire [7:0] t_r35_c60_0;
  wire [7:0] t_r35_c60_1;
  wire [7:0] t_r35_c60_2;
  wire [7:0] t_r35_c60_3;
  wire [7:0] t_r35_c60_4;
  wire [7:0] t_r35_c60_5;
  wire [7:0] t_r35_c60_6;
  wire [7:0] t_r35_c60_7;
  wire [7:0] t_r35_c60_8;
  wire [7:0] t_r35_c60_9;
  wire [7:0] t_r35_c60_10;
  wire [7:0] t_r35_c60_11;
  wire [7:0] t_r35_c60_12;
  wire [7:0] t_r35_c61_0;
  wire [7:0] t_r35_c61_1;
  wire [7:0] t_r35_c61_2;
  wire [7:0] t_r35_c61_3;
  wire [7:0] t_r35_c61_4;
  wire [7:0] t_r35_c61_5;
  wire [7:0] t_r35_c61_6;
  wire [7:0] t_r35_c61_7;
  wire [7:0] t_r35_c61_8;
  wire [7:0] t_r35_c61_9;
  wire [7:0] t_r35_c61_10;
  wire [7:0] t_r35_c61_11;
  wire [7:0] t_r35_c61_12;
  wire [7:0] t_r35_c62_0;
  wire [7:0] t_r35_c62_1;
  wire [7:0] t_r35_c62_2;
  wire [7:0] t_r35_c62_3;
  wire [7:0] t_r35_c62_4;
  wire [7:0] t_r35_c62_5;
  wire [7:0] t_r35_c62_6;
  wire [7:0] t_r35_c62_7;
  wire [7:0] t_r35_c62_8;
  wire [7:0] t_r35_c62_9;
  wire [7:0] t_r35_c62_10;
  wire [7:0] t_r35_c62_11;
  wire [7:0] t_r35_c62_12;
  wire [7:0] t_r35_c63_0;
  wire [7:0] t_r35_c63_1;
  wire [7:0] t_r35_c63_2;
  wire [7:0] t_r35_c63_3;
  wire [7:0] t_r35_c63_4;
  wire [7:0] t_r35_c63_5;
  wire [7:0] t_r35_c63_6;
  wire [7:0] t_r35_c63_7;
  wire [7:0] t_r35_c63_8;
  wire [7:0] t_r35_c63_9;
  wire [7:0] t_r35_c63_10;
  wire [7:0] t_r35_c63_11;
  wire [7:0] t_r35_c63_12;
  wire [7:0] t_r35_c64_0;
  wire [7:0] t_r35_c64_1;
  wire [7:0] t_r35_c64_2;
  wire [7:0] t_r35_c64_3;
  wire [7:0] t_r35_c64_4;
  wire [7:0] t_r35_c64_5;
  wire [7:0] t_r35_c64_6;
  wire [7:0] t_r35_c64_7;
  wire [7:0] t_r35_c64_8;
  wire [7:0] t_r35_c64_9;
  wire [7:0] t_r35_c64_10;
  wire [7:0] t_r35_c64_11;
  wire [7:0] t_r35_c64_12;
  wire [7:0] t_r35_c65_0;
  wire [7:0] t_r35_c65_1;
  wire [7:0] t_r35_c65_2;
  wire [7:0] t_r35_c65_3;
  wire [7:0] t_r35_c65_4;
  wire [7:0] t_r35_c65_5;
  wire [7:0] t_r35_c65_6;
  wire [7:0] t_r35_c65_7;
  wire [7:0] t_r35_c65_8;
  wire [7:0] t_r35_c65_9;
  wire [7:0] t_r35_c65_10;
  wire [7:0] t_r35_c65_11;
  wire [7:0] t_r35_c65_12;
  wire [7:0] t_r36_c0_0;
  wire [7:0] t_r36_c0_1;
  wire [7:0] t_r36_c0_2;
  wire [7:0] t_r36_c0_3;
  wire [7:0] t_r36_c0_4;
  wire [7:0] t_r36_c0_5;
  wire [7:0] t_r36_c0_6;
  wire [7:0] t_r36_c0_7;
  wire [7:0] t_r36_c0_8;
  wire [7:0] t_r36_c0_9;
  wire [7:0] t_r36_c0_10;
  wire [7:0] t_r36_c0_11;
  wire [7:0] t_r36_c0_12;
  wire [7:0] t_r36_c1_0;
  wire [7:0] t_r36_c1_1;
  wire [7:0] t_r36_c1_2;
  wire [7:0] t_r36_c1_3;
  wire [7:0] t_r36_c1_4;
  wire [7:0] t_r36_c1_5;
  wire [7:0] t_r36_c1_6;
  wire [7:0] t_r36_c1_7;
  wire [7:0] t_r36_c1_8;
  wire [7:0] t_r36_c1_9;
  wire [7:0] t_r36_c1_10;
  wire [7:0] t_r36_c1_11;
  wire [7:0] t_r36_c1_12;
  wire [7:0] t_r36_c2_0;
  wire [7:0] t_r36_c2_1;
  wire [7:0] t_r36_c2_2;
  wire [7:0] t_r36_c2_3;
  wire [7:0] t_r36_c2_4;
  wire [7:0] t_r36_c2_5;
  wire [7:0] t_r36_c2_6;
  wire [7:0] t_r36_c2_7;
  wire [7:0] t_r36_c2_8;
  wire [7:0] t_r36_c2_9;
  wire [7:0] t_r36_c2_10;
  wire [7:0] t_r36_c2_11;
  wire [7:0] t_r36_c2_12;
  wire [7:0] t_r36_c3_0;
  wire [7:0] t_r36_c3_1;
  wire [7:0] t_r36_c3_2;
  wire [7:0] t_r36_c3_3;
  wire [7:0] t_r36_c3_4;
  wire [7:0] t_r36_c3_5;
  wire [7:0] t_r36_c3_6;
  wire [7:0] t_r36_c3_7;
  wire [7:0] t_r36_c3_8;
  wire [7:0] t_r36_c3_9;
  wire [7:0] t_r36_c3_10;
  wire [7:0] t_r36_c3_11;
  wire [7:0] t_r36_c3_12;
  wire [7:0] t_r36_c4_0;
  wire [7:0] t_r36_c4_1;
  wire [7:0] t_r36_c4_2;
  wire [7:0] t_r36_c4_3;
  wire [7:0] t_r36_c4_4;
  wire [7:0] t_r36_c4_5;
  wire [7:0] t_r36_c4_6;
  wire [7:0] t_r36_c4_7;
  wire [7:0] t_r36_c4_8;
  wire [7:0] t_r36_c4_9;
  wire [7:0] t_r36_c4_10;
  wire [7:0] t_r36_c4_11;
  wire [7:0] t_r36_c4_12;
  wire [7:0] t_r36_c5_0;
  wire [7:0] t_r36_c5_1;
  wire [7:0] t_r36_c5_2;
  wire [7:0] t_r36_c5_3;
  wire [7:0] t_r36_c5_4;
  wire [7:0] t_r36_c5_5;
  wire [7:0] t_r36_c5_6;
  wire [7:0] t_r36_c5_7;
  wire [7:0] t_r36_c5_8;
  wire [7:0] t_r36_c5_9;
  wire [7:0] t_r36_c5_10;
  wire [7:0] t_r36_c5_11;
  wire [7:0] t_r36_c5_12;
  wire [7:0] t_r36_c6_0;
  wire [7:0] t_r36_c6_1;
  wire [7:0] t_r36_c6_2;
  wire [7:0] t_r36_c6_3;
  wire [7:0] t_r36_c6_4;
  wire [7:0] t_r36_c6_5;
  wire [7:0] t_r36_c6_6;
  wire [7:0] t_r36_c6_7;
  wire [7:0] t_r36_c6_8;
  wire [7:0] t_r36_c6_9;
  wire [7:0] t_r36_c6_10;
  wire [7:0] t_r36_c6_11;
  wire [7:0] t_r36_c6_12;
  wire [7:0] t_r36_c7_0;
  wire [7:0] t_r36_c7_1;
  wire [7:0] t_r36_c7_2;
  wire [7:0] t_r36_c7_3;
  wire [7:0] t_r36_c7_4;
  wire [7:0] t_r36_c7_5;
  wire [7:0] t_r36_c7_6;
  wire [7:0] t_r36_c7_7;
  wire [7:0] t_r36_c7_8;
  wire [7:0] t_r36_c7_9;
  wire [7:0] t_r36_c7_10;
  wire [7:0] t_r36_c7_11;
  wire [7:0] t_r36_c7_12;
  wire [7:0] t_r36_c8_0;
  wire [7:0] t_r36_c8_1;
  wire [7:0] t_r36_c8_2;
  wire [7:0] t_r36_c8_3;
  wire [7:0] t_r36_c8_4;
  wire [7:0] t_r36_c8_5;
  wire [7:0] t_r36_c8_6;
  wire [7:0] t_r36_c8_7;
  wire [7:0] t_r36_c8_8;
  wire [7:0] t_r36_c8_9;
  wire [7:0] t_r36_c8_10;
  wire [7:0] t_r36_c8_11;
  wire [7:0] t_r36_c8_12;
  wire [7:0] t_r36_c9_0;
  wire [7:0] t_r36_c9_1;
  wire [7:0] t_r36_c9_2;
  wire [7:0] t_r36_c9_3;
  wire [7:0] t_r36_c9_4;
  wire [7:0] t_r36_c9_5;
  wire [7:0] t_r36_c9_6;
  wire [7:0] t_r36_c9_7;
  wire [7:0] t_r36_c9_8;
  wire [7:0] t_r36_c9_9;
  wire [7:0] t_r36_c9_10;
  wire [7:0] t_r36_c9_11;
  wire [7:0] t_r36_c9_12;
  wire [7:0] t_r36_c10_0;
  wire [7:0] t_r36_c10_1;
  wire [7:0] t_r36_c10_2;
  wire [7:0] t_r36_c10_3;
  wire [7:0] t_r36_c10_4;
  wire [7:0] t_r36_c10_5;
  wire [7:0] t_r36_c10_6;
  wire [7:0] t_r36_c10_7;
  wire [7:0] t_r36_c10_8;
  wire [7:0] t_r36_c10_9;
  wire [7:0] t_r36_c10_10;
  wire [7:0] t_r36_c10_11;
  wire [7:0] t_r36_c10_12;
  wire [7:0] t_r36_c11_0;
  wire [7:0] t_r36_c11_1;
  wire [7:0] t_r36_c11_2;
  wire [7:0] t_r36_c11_3;
  wire [7:0] t_r36_c11_4;
  wire [7:0] t_r36_c11_5;
  wire [7:0] t_r36_c11_6;
  wire [7:0] t_r36_c11_7;
  wire [7:0] t_r36_c11_8;
  wire [7:0] t_r36_c11_9;
  wire [7:0] t_r36_c11_10;
  wire [7:0] t_r36_c11_11;
  wire [7:0] t_r36_c11_12;
  wire [7:0] t_r36_c12_0;
  wire [7:0] t_r36_c12_1;
  wire [7:0] t_r36_c12_2;
  wire [7:0] t_r36_c12_3;
  wire [7:0] t_r36_c12_4;
  wire [7:0] t_r36_c12_5;
  wire [7:0] t_r36_c12_6;
  wire [7:0] t_r36_c12_7;
  wire [7:0] t_r36_c12_8;
  wire [7:0] t_r36_c12_9;
  wire [7:0] t_r36_c12_10;
  wire [7:0] t_r36_c12_11;
  wire [7:0] t_r36_c12_12;
  wire [7:0] t_r36_c13_0;
  wire [7:0] t_r36_c13_1;
  wire [7:0] t_r36_c13_2;
  wire [7:0] t_r36_c13_3;
  wire [7:0] t_r36_c13_4;
  wire [7:0] t_r36_c13_5;
  wire [7:0] t_r36_c13_6;
  wire [7:0] t_r36_c13_7;
  wire [7:0] t_r36_c13_8;
  wire [7:0] t_r36_c13_9;
  wire [7:0] t_r36_c13_10;
  wire [7:0] t_r36_c13_11;
  wire [7:0] t_r36_c13_12;
  wire [7:0] t_r36_c14_0;
  wire [7:0] t_r36_c14_1;
  wire [7:0] t_r36_c14_2;
  wire [7:0] t_r36_c14_3;
  wire [7:0] t_r36_c14_4;
  wire [7:0] t_r36_c14_5;
  wire [7:0] t_r36_c14_6;
  wire [7:0] t_r36_c14_7;
  wire [7:0] t_r36_c14_8;
  wire [7:0] t_r36_c14_9;
  wire [7:0] t_r36_c14_10;
  wire [7:0] t_r36_c14_11;
  wire [7:0] t_r36_c14_12;
  wire [7:0] t_r36_c15_0;
  wire [7:0] t_r36_c15_1;
  wire [7:0] t_r36_c15_2;
  wire [7:0] t_r36_c15_3;
  wire [7:0] t_r36_c15_4;
  wire [7:0] t_r36_c15_5;
  wire [7:0] t_r36_c15_6;
  wire [7:0] t_r36_c15_7;
  wire [7:0] t_r36_c15_8;
  wire [7:0] t_r36_c15_9;
  wire [7:0] t_r36_c15_10;
  wire [7:0] t_r36_c15_11;
  wire [7:0] t_r36_c15_12;
  wire [7:0] t_r36_c16_0;
  wire [7:0] t_r36_c16_1;
  wire [7:0] t_r36_c16_2;
  wire [7:0] t_r36_c16_3;
  wire [7:0] t_r36_c16_4;
  wire [7:0] t_r36_c16_5;
  wire [7:0] t_r36_c16_6;
  wire [7:0] t_r36_c16_7;
  wire [7:0] t_r36_c16_8;
  wire [7:0] t_r36_c16_9;
  wire [7:0] t_r36_c16_10;
  wire [7:0] t_r36_c16_11;
  wire [7:0] t_r36_c16_12;
  wire [7:0] t_r36_c17_0;
  wire [7:0] t_r36_c17_1;
  wire [7:0] t_r36_c17_2;
  wire [7:0] t_r36_c17_3;
  wire [7:0] t_r36_c17_4;
  wire [7:0] t_r36_c17_5;
  wire [7:0] t_r36_c17_6;
  wire [7:0] t_r36_c17_7;
  wire [7:0] t_r36_c17_8;
  wire [7:0] t_r36_c17_9;
  wire [7:0] t_r36_c17_10;
  wire [7:0] t_r36_c17_11;
  wire [7:0] t_r36_c17_12;
  wire [7:0] t_r36_c18_0;
  wire [7:0] t_r36_c18_1;
  wire [7:0] t_r36_c18_2;
  wire [7:0] t_r36_c18_3;
  wire [7:0] t_r36_c18_4;
  wire [7:0] t_r36_c18_5;
  wire [7:0] t_r36_c18_6;
  wire [7:0] t_r36_c18_7;
  wire [7:0] t_r36_c18_8;
  wire [7:0] t_r36_c18_9;
  wire [7:0] t_r36_c18_10;
  wire [7:0] t_r36_c18_11;
  wire [7:0] t_r36_c18_12;
  wire [7:0] t_r36_c19_0;
  wire [7:0] t_r36_c19_1;
  wire [7:0] t_r36_c19_2;
  wire [7:0] t_r36_c19_3;
  wire [7:0] t_r36_c19_4;
  wire [7:0] t_r36_c19_5;
  wire [7:0] t_r36_c19_6;
  wire [7:0] t_r36_c19_7;
  wire [7:0] t_r36_c19_8;
  wire [7:0] t_r36_c19_9;
  wire [7:0] t_r36_c19_10;
  wire [7:0] t_r36_c19_11;
  wire [7:0] t_r36_c19_12;
  wire [7:0] t_r36_c20_0;
  wire [7:0] t_r36_c20_1;
  wire [7:0] t_r36_c20_2;
  wire [7:0] t_r36_c20_3;
  wire [7:0] t_r36_c20_4;
  wire [7:0] t_r36_c20_5;
  wire [7:0] t_r36_c20_6;
  wire [7:0] t_r36_c20_7;
  wire [7:0] t_r36_c20_8;
  wire [7:0] t_r36_c20_9;
  wire [7:0] t_r36_c20_10;
  wire [7:0] t_r36_c20_11;
  wire [7:0] t_r36_c20_12;
  wire [7:0] t_r36_c21_0;
  wire [7:0] t_r36_c21_1;
  wire [7:0] t_r36_c21_2;
  wire [7:0] t_r36_c21_3;
  wire [7:0] t_r36_c21_4;
  wire [7:0] t_r36_c21_5;
  wire [7:0] t_r36_c21_6;
  wire [7:0] t_r36_c21_7;
  wire [7:0] t_r36_c21_8;
  wire [7:0] t_r36_c21_9;
  wire [7:0] t_r36_c21_10;
  wire [7:0] t_r36_c21_11;
  wire [7:0] t_r36_c21_12;
  wire [7:0] t_r36_c22_0;
  wire [7:0] t_r36_c22_1;
  wire [7:0] t_r36_c22_2;
  wire [7:0] t_r36_c22_3;
  wire [7:0] t_r36_c22_4;
  wire [7:0] t_r36_c22_5;
  wire [7:0] t_r36_c22_6;
  wire [7:0] t_r36_c22_7;
  wire [7:0] t_r36_c22_8;
  wire [7:0] t_r36_c22_9;
  wire [7:0] t_r36_c22_10;
  wire [7:0] t_r36_c22_11;
  wire [7:0] t_r36_c22_12;
  wire [7:0] t_r36_c23_0;
  wire [7:0] t_r36_c23_1;
  wire [7:0] t_r36_c23_2;
  wire [7:0] t_r36_c23_3;
  wire [7:0] t_r36_c23_4;
  wire [7:0] t_r36_c23_5;
  wire [7:0] t_r36_c23_6;
  wire [7:0] t_r36_c23_7;
  wire [7:0] t_r36_c23_8;
  wire [7:0] t_r36_c23_9;
  wire [7:0] t_r36_c23_10;
  wire [7:0] t_r36_c23_11;
  wire [7:0] t_r36_c23_12;
  wire [7:0] t_r36_c24_0;
  wire [7:0] t_r36_c24_1;
  wire [7:0] t_r36_c24_2;
  wire [7:0] t_r36_c24_3;
  wire [7:0] t_r36_c24_4;
  wire [7:0] t_r36_c24_5;
  wire [7:0] t_r36_c24_6;
  wire [7:0] t_r36_c24_7;
  wire [7:0] t_r36_c24_8;
  wire [7:0] t_r36_c24_9;
  wire [7:0] t_r36_c24_10;
  wire [7:0] t_r36_c24_11;
  wire [7:0] t_r36_c24_12;
  wire [7:0] t_r36_c25_0;
  wire [7:0] t_r36_c25_1;
  wire [7:0] t_r36_c25_2;
  wire [7:0] t_r36_c25_3;
  wire [7:0] t_r36_c25_4;
  wire [7:0] t_r36_c25_5;
  wire [7:0] t_r36_c25_6;
  wire [7:0] t_r36_c25_7;
  wire [7:0] t_r36_c25_8;
  wire [7:0] t_r36_c25_9;
  wire [7:0] t_r36_c25_10;
  wire [7:0] t_r36_c25_11;
  wire [7:0] t_r36_c25_12;
  wire [7:0] t_r36_c26_0;
  wire [7:0] t_r36_c26_1;
  wire [7:0] t_r36_c26_2;
  wire [7:0] t_r36_c26_3;
  wire [7:0] t_r36_c26_4;
  wire [7:0] t_r36_c26_5;
  wire [7:0] t_r36_c26_6;
  wire [7:0] t_r36_c26_7;
  wire [7:0] t_r36_c26_8;
  wire [7:0] t_r36_c26_9;
  wire [7:0] t_r36_c26_10;
  wire [7:0] t_r36_c26_11;
  wire [7:0] t_r36_c26_12;
  wire [7:0] t_r36_c27_0;
  wire [7:0] t_r36_c27_1;
  wire [7:0] t_r36_c27_2;
  wire [7:0] t_r36_c27_3;
  wire [7:0] t_r36_c27_4;
  wire [7:0] t_r36_c27_5;
  wire [7:0] t_r36_c27_6;
  wire [7:0] t_r36_c27_7;
  wire [7:0] t_r36_c27_8;
  wire [7:0] t_r36_c27_9;
  wire [7:0] t_r36_c27_10;
  wire [7:0] t_r36_c27_11;
  wire [7:0] t_r36_c27_12;
  wire [7:0] t_r36_c28_0;
  wire [7:0] t_r36_c28_1;
  wire [7:0] t_r36_c28_2;
  wire [7:0] t_r36_c28_3;
  wire [7:0] t_r36_c28_4;
  wire [7:0] t_r36_c28_5;
  wire [7:0] t_r36_c28_6;
  wire [7:0] t_r36_c28_7;
  wire [7:0] t_r36_c28_8;
  wire [7:0] t_r36_c28_9;
  wire [7:0] t_r36_c28_10;
  wire [7:0] t_r36_c28_11;
  wire [7:0] t_r36_c28_12;
  wire [7:0] t_r36_c29_0;
  wire [7:0] t_r36_c29_1;
  wire [7:0] t_r36_c29_2;
  wire [7:0] t_r36_c29_3;
  wire [7:0] t_r36_c29_4;
  wire [7:0] t_r36_c29_5;
  wire [7:0] t_r36_c29_6;
  wire [7:0] t_r36_c29_7;
  wire [7:0] t_r36_c29_8;
  wire [7:0] t_r36_c29_9;
  wire [7:0] t_r36_c29_10;
  wire [7:0] t_r36_c29_11;
  wire [7:0] t_r36_c29_12;
  wire [7:0] t_r36_c30_0;
  wire [7:0] t_r36_c30_1;
  wire [7:0] t_r36_c30_2;
  wire [7:0] t_r36_c30_3;
  wire [7:0] t_r36_c30_4;
  wire [7:0] t_r36_c30_5;
  wire [7:0] t_r36_c30_6;
  wire [7:0] t_r36_c30_7;
  wire [7:0] t_r36_c30_8;
  wire [7:0] t_r36_c30_9;
  wire [7:0] t_r36_c30_10;
  wire [7:0] t_r36_c30_11;
  wire [7:0] t_r36_c30_12;
  wire [7:0] t_r36_c31_0;
  wire [7:0] t_r36_c31_1;
  wire [7:0] t_r36_c31_2;
  wire [7:0] t_r36_c31_3;
  wire [7:0] t_r36_c31_4;
  wire [7:0] t_r36_c31_5;
  wire [7:0] t_r36_c31_6;
  wire [7:0] t_r36_c31_7;
  wire [7:0] t_r36_c31_8;
  wire [7:0] t_r36_c31_9;
  wire [7:0] t_r36_c31_10;
  wire [7:0] t_r36_c31_11;
  wire [7:0] t_r36_c31_12;
  wire [7:0] t_r36_c32_0;
  wire [7:0] t_r36_c32_1;
  wire [7:0] t_r36_c32_2;
  wire [7:0] t_r36_c32_3;
  wire [7:0] t_r36_c32_4;
  wire [7:0] t_r36_c32_5;
  wire [7:0] t_r36_c32_6;
  wire [7:0] t_r36_c32_7;
  wire [7:0] t_r36_c32_8;
  wire [7:0] t_r36_c32_9;
  wire [7:0] t_r36_c32_10;
  wire [7:0] t_r36_c32_11;
  wire [7:0] t_r36_c32_12;
  wire [7:0] t_r36_c33_0;
  wire [7:0] t_r36_c33_1;
  wire [7:0] t_r36_c33_2;
  wire [7:0] t_r36_c33_3;
  wire [7:0] t_r36_c33_4;
  wire [7:0] t_r36_c33_5;
  wire [7:0] t_r36_c33_6;
  wire [7:0] t_r36_c33_7;
  wire [7:0] t_r36_c33_8;
  wire [7:0] t_r36_c33_9;
  wire [7:0] t_r36_c33_10;
  wire [7:0] t_r36_c33_11;
  wire [7:0] t_r36_c33_12;
  wire [7:0] t_r36_c34_0;
  wire [7:0] t_r36_c34_1;
  wire [7:0] t_r36_c34_2;
  wire [7:0] t_r36_c34_3;
  wire [7:0] t_r36_c34_4;
  wire [7:0] t_r36_c34_5;
  wire [7:0] t_r36_c34_6;
  wire [7:0] t_r36_c34_7;
  wire [7:0] t_r36_c34_8;
  wire [7:0] t_r36_c34_9;
  wire [7:0] t_r36_c34_10;
  wire [7:0] t_r36_c34_11;
  wire [7:0] t_r36_c34_12;
  wire [7:0] t_r36_c35_0;
  wire [7:0] t_r36_c35_1;
  wire [7:0] t_r36_c35_2;
  wire [7:0] t_r36_c35_3;
  wire [7:0] t_r36_c35_4;
  wire [7:0] t_r36_c35_5;
  wire [7:0] t_r36_c35_6;
  wire [7:0] t_r36_c35_7;
  wire [7:0] t_r36_c35_8;
  wire [7:0] t_r36_c35_9;
  wire [7:0] t_r36_c35_10;
  wire [7:0] t_r36_c35_11;
  wire [7:0] t_r36_c35_12;
  wire [7:0] t_r36_c36_0;
  wire [7:0] t_r36_c36_1;
  wire [7:0] t_r36_c36_2;
  wire [7:0] t_r36_c36_3;
  wire [7:0] t_r36_c36_4;
  wire [7:0] t_r36_c36_5;
  wire [7:0] t_r36_c36_6;
  wire [7:0] t_r36_c36_7;
  wire [7:0] t_r36_c36_8;
  wire [7:0] t_r36_c36_9;
  wire [7:0] t_r36_c36_10;
  wire [7:0] t_r36_c36_11;
  wire [7:0] t_r36_c36_12;
  wire [7:0] t_r36_c37_0;
  wire [7:0] t_r36_c37_1;
  wire [7:0] t_r36_c37_2;
  wire [7:0] t_r36_c37_3;
  wire [7:0] t_r36_c37_4;
  wire [7:0] t_r36_c37_5;
  wire [7:0] t_r36_c37_6;
  wire [7:0] t_r36_c37_7;
  wire [7:0] t_r36_c37_8;
  wire [7:0] t_r36_c37_9;
  wire [7:0] t_r36_c37_10;
  wire [7:0] t_r36_c37_11;
  wire [7:0] t_r36_c37_12;
  wire [7:0] t_r36_c38_0;
  wire [7:0] t_r36_c38_1;
  wire [7:0] t_r36_c38_2;
  wire [7:0] t_r36_c38_3;
  wire [7:0] t_r36_c38_4;
  wire [7:0] t_r36_c38_5;
  wire [7:0] t_r36_c38_6;
  wire [7:0] t_r36_c38_7;
  wire [7:0] t_r36_c38_8;
  wire [7:0] t_r36_c38_9;
  wire [7:0] t_r36_c38_10;
  wire [7:0] t_r36_c38_11;
  wire [7:0] t_r36_c38_12;
  wire [7:0] t_r36_c39_0;
  wire [7:0] t_r36_c39_1;
  wire [7:0] t_r36_c39_2;
  wire [7:0] t_r36_c39_3;
  wire [7:0] t_r36_c39_4;
  wire [7:0] t_r36_c39_5;
  wire [7:0] t_r36_c39_6;
  wire [7:0] t_r36_c39_7;
  wire [7:0] t_r36_c39_8;
  wire [7:0] t_r36_c39_9;
  wire [7:0] t_r36_c39_10;
  wire [7:0] t_r36_c39_11;
  wire [7:0] t_r36_c39_12;
  wire [7:0] t_r36_c40_0;
  wire [7:0] t_r36_c40_1;
  wire [7:0] t_r36_c40_2;
  wire [7:0] t_r36_c40_3;
  wire [7:0] t_r36_c40_4;
  wire [7:0] t_r36_c40_5;
  wire [7:0] t_r36_c40_6;
  wire [7:0] t_r36_c40_7;
  wire [7:0] t_r36_c40_8;
  wire [7:0] t_r36_c40_9;
  wire [7:0] t_r36_c40_10;
  wire [7:0] t_r36_c40_11;
  wire [7:0] t_r36_c40_12;
  wire [7:0] t_r36_c41_0;
  wire [7:0] t_r36_c41_1;
  wire [7:0] t_r36_c41_2;
  wire [7:0] t_r36_c41_3;
  wire [7:0] t_r36_c41_4;
  wire [7:0] t_r36_c41_5;
  wire [7:0] t_r36_c41_6;
  wire [7:0] t_r36_c41_7;
  wire [7:0] t_r36_c41_8;
  wire [7:0] t_r36_c41_9;
  wire [7:0] t_r36_c41_10;
  wire [7:0] t_r36_c41_11;
  wire [7:0] t_r36_c41_12;
  wire [7:0] t_r36_c42_0;
  wire [7:0] t_r36_c42_1;
  wire [7:0] t_r36_c42_2;
  wire [7:0] t_r36_c42_3;
  wire [7:0] t_r36_c42_4;
  wire [7:0] t_r36_c42_5;
  wire [7:0] t_r36_c42_6;
  wire [7:0] t_r36_c42_7;
  wire [7:0] t_r36_c42_8;
  wire [7:0] t_r36_c42_9;
  wire [7:0] t_r36_c42_10;
  wire [7:0] t_r36_c42_11;
  wire [7:0] t_r36_c42_12;
  wire [7:0] t_r36_c43_0;
  wire [7:0] t_r36_c43_1;
  wire [7:0] t_r36_c43_2;
  wire [7:0] t_r36_c43_3;
  wire [7:0] t_r36_c43_4;
  wire [7:0] t_r36_c43_5;
  wire [7:0] t_r36_c43_6;
  wire [7:0] t_r36_c43_7;
  wire [7:0] t_r36_c43_8;
  wire [7:0] t_r36_c43_9;
  wire [7:0] t_r36_c43_10;
  wire [7:0] t_r36_c43_11;
  wire [7:0] t_r36_c43_12;
  wire [7:0] t_r36_c44_0;
  wire [7:0] t_r36_c44_1;
  wire [7:0] t_r36_c44_2;
  wire [7:0] t_r36_c44_3;
  wire [7:0] t_r36_c44_4;
  wire [7:0] t_r36_c44_5;
  wire [7:0] t_r36_c44_6;
  wire [7:0] t_r36_c44_7;
  wire [7:0] t_r36_c44_8;
  wire [7:0] t_r36_c44_9;
  wire [7:0] t_r36_c44_10;
  wire [7:0] t_r36_c44_11;
  wire [7:0] t_r36_c44_12;
  wire [7:0] t_r36_c45_0;
  wire [7:0] t_r36_c45_1;
  wire [7:0] t_r36_c45_2;
  wire [7:0] t_r36_c45_3;
  wire [7:0] t_r36_c45_4;
  wire [7:0] t_r36_c45_5;
  wire [7:0] t_r36_c45_6;
  wire [7:0] t_r36_c45_7;
  wire [7:0] t_r36_c45_8;
  wire [7:0] t_r36_c45_9;
  wire [7:0] t_r36_c45_10;
  wire [7:0] t_r36_c45_11;
  wire [7:0] t_r36_c45_12;
  wire [7:0] t_r36_c46_0;
  wire [7:0] t_r36_c46_1;
  wire [7:0] t_r36_c46_2;
  wire [7:0] t_r36_c46_3;
  wire [7:0] t_r36_c46_4;
  wire [7:0] t_r36_c46_5;
  wire [7:0] t_r36_c46_6;
  wire [7:0] t_r36_c46_7;
  wire [7:0] t_r36_c46_8;
  wire [7:0] t_r36_c46_9;
  wire [7:0] t_r36_c46_10;
  wire [7:0] t_r36_c46_11;
  wire [7:0] t_r36_c46_12;
  wire [7:0] t_r36_c47_0;
  wire [7:0] t_r36_c47_1;
  wire [7:0] t_r36_c47_2;
  wire [7:0] t_r36_c47_3;
  wire [7:0] t_r36_c47_4;
  wire [7:0] t_r36_c47_5;
  wire [7:0] t_r36_c47_6;
  wire [7:0] t_r36_c47_7;
  wire [7:0] t_r36_c47_8;
  wire [7:0] t_r36_c47_9;
  wire [7:0] t_r36_c47_10;
  wire [7:0] t_r36_c47_11;
  wire [7:0] t_r36_c47_12;
  wire [7:0] t_r36_c48_0;
  wire [7:0] t_r36_c48_1;
  wire [7:0] t_r36_c48_2;
  wire [7:0] t_r36_c48_3;
  wire [7:0] t_r36_c48_4;
  wire [7:0] t_r36_c48_5;
  wire [7:0] t_r36_c48_6;
  wire [7:0] t_r36_c48_7;
  wire [7:0] t_r36_c48_8;
  wire [7:0] t_r36_c48_9;
  wire [7:0] t_r36_c48_10;
  wire [7:0] t_r36_c48_11;
  wire [7:0] t_r36_c48_12;
  wire [7:0] t_r36_c49_0;
  wire [7:0] t_r36_c49_1;
  wire [7:0] t_r36_c49_2;
  wire [7:0] t_r36_c49_3;
  wire [7:0] t_r36_c49_4;
  wire [7:0] t_r36_c49_5;
  wire [7:0] t_r36_c49_6;
  wire [7:0] t_r36_c49_7;
  wire [7:0] t_r36_c49_8;
  wire [7:0] t_r36_c49_9;
  wire [7:0] t_r36_c49_10;
  wire [7:0] t_r36_c49_11;
  wire [7:0] t_r36_c49_12;
  wire [7:0] t_r36_c50_0;
  wire [7:0] t_r36_c50_1;
  wire [7:0] t_r36_c50_2;
  wire [7:0] t_r36_c50_3;
  wire [7:0] t_r36_c50_4;
  wire [7:0] t_r36_c50_5;
  wire [7:0] t_r36_c50_6;
  wire [7:0] t_r36_c50_7;
  wire [7:0] t_r36_c50_8;
  wire [7:0] t_r36_c50_9;
  wire [7:0] t_r36_c50_10;
  wire [7:0] t_r36_c50_11;
  wire [7:0] t_r36_c50_12;
  wire [7:0] t_r36_c51_0;
  wire [7:0] t_r36_c51_1;
  wire [7:0] t_r36_c51_2;
  wire [7:0] t_r36_c51_3;
  wire [7:0] t_r36_c51_4;
  wire [7:0] t_r36_c51_5;
  wire [7:0] t_r36_c51_6;
  wire [7:0] t_r36_c51_7;
  wire [7:0] t_r36_c51_8;
  wire [7:0] t_r36_c51_9;
  wire [7:0] t_r36_c51_10;
  wire [7:0] t_r36_c51_11;
  wire [7:0] t_r36_c51_12;
  wire [7:0] t_r36_c52_0;
  wire [7:0] t_r36_c52_1;
  wire [7:0] t_r36_c52_2;
  wire [7:0] t_r36_c52_3;
  wire [7:0] t_r36_c52_4;
  wire [7:0] t_r36_c52_5;
  wire [7:0] t_r36_c52_6;
  wire [7:0] t_r36_c52_7;
  wire [7:0] t_r36_c52_8;
  wire [7:0] t_r36_c52_9;
  wire [7:0] t_r36_c52_10;
  wire [7:0] t_r36_c52_11;
  wire [7:0] t_r36_c52_12;
  wire [7:0] t_r36_c53_0;
  wire [7:0] t_r36_c53_1;
  wire [7:0] t_r36_c53_2;
  wire [7:0] t_r36_c53_3;
  wire [7:0] t_r36_c53_4;
  wire [7:0] t_r36_c53_5;
  wire [7:0] t_r36_c53_6;
  wire [7:0] t_r36_c53_7;
  wire [7:0] t_r36_c53_8;
  wire [7:0] t_r36_c53_9;
  wire [7:0] t_r36_c53_10;
  wire [7:0] t_r36_c53_11;
  wire [7:0] t_r36_c53_12;
  wire [7:0] t_r36_c54_0;
  wire [7:0] t_r36_c54_1;
  wire [7:0] t_r36_c54_2;
  wire [7:0] t_r36_c54_3;
  wire [7:0] t_r36_c54_4;
  wire [7:0] t_r36_c54_5;
  wire [7:0] t_r36_c54_6;
  wire [7:0] t_r36_c54_7;
  wire [7:0] t_r36_c54_8;
  wire [7:0] t_r36_c54_9;
  wire [7:0] t_r36_c54_10;
  wire [7:0] t_r36_c54_11;
  wire [7:0] t_r36_c54_12;
  wire [7:0] t_r36_c55_0;
  wire [7:0] t_r36_c55_1;
  wire [7:0] t_r36_c55_2;
  wire [7:0] t_r36_c55_3;
  wire [7:0] t_r36_c55_4;
  wire [7:0] t_r36_c55_5;
  wire [7:0] t_r36_c55_6;
  wire [7:0] t_r36_c55_7;
  wire [7:0] t_r36_c55_8;
  wire [7:0] t_r36_c55_9;
  wire [7:0] t_r36_c55_10;
  wire [7:0] t_r36_c55_11;
  wire [7:0] t_r36_c55_12;
  wire [7:0] t_r36_c56_0;
  wire [7:0] t_r36_c56_1;
  wire [7:0] t_r36_c56_2;
  wire [7:0] t_r36_c56_3;
  wire [7:0] t_r36_c56_4;
  wire [7:0] t_r36_c56_5;
  wire [7:0] t_r36_c56_6;
  wire [7:0] t_r36_c56_7;
  wire [7:0] t_r36_c56_8;
  wire [7:0] t_r36_c56_9;
  wire [7:0] t_r36_c56_10;
  wire [7:0] t_r36_c56_11;
  wire [7:0] t_r36_c56_12;
  wire [7:0] t_r36_c57_0;
  wire [7:0] t_r36_c57_1;
  wire [7:0] t_r36_c57_2;
  wire [7:0] t_r36_c57_3;
  wire [7:0] t_r36_c57_4;
  wire [7:0] t_r36_c57_5;
  wire [7:0] t_r36_c57_6;
  wire [7:0] t_r36_c57_7;
  wire [7:0] t_r36_c57_8;
  wire [7:0] t_r36_c57_9;
  wire [7:0] t_r36_c57_10;
  wire [7:0] t_r36_c57_11;
  wire [7:0] t_r36_c57_12;
  wire [7:0] t_r36_c58_0;
  wire [7:0] t_r36_c58_1;
  wire [7:0] t_r36_c58_2;
  wire [7:0] t_r36_c58_3;
  wire [7:0] t_r36_c58_4;
  wire [7:0] t_r36_c58_5;
  wire [7:0] t_r36_c58_6;
  wire [7:0] t_r36_c58_7;
  wire [7:0] t_r36_c58_8;
  wire [7:0] t_r36_c58_9;
  wire [7:0] t_r36_c58_10;
  wire [7:0] t_r36_c58_11;
  wire [7:0] t_r36_c58_12;
  wire [7:0] t_r36_c59_0;
  wire [7:0] t_r36_c59_1;
  wire [7:0] t_r36_c59_2;
  wire [7:0] t_r36_c59_3;
  wire [7:0] t_r36_c59_4;
  wire [7:0] t_r36_c59_5;
  wire [7:0] t_r36_c59_6;
  wire [7:0] t_r36_c59_7;
  wire [7:0] t_r36_c59_8;
  wire [7:0] t_r36_c59_9;
  wire [7:0] t_r36_c59_10;
  wire [7:0] t_r36_c59_11;
  wire [7:0] t_r36_c59_12;
  wire [7:0] t_r36_c60_0;
  wire [7:0] t_r36_c60_1;
  wire [7:0] t_r36_c60_2;
  wire [7:0] t_r36_c60_3;
  wire [7:0] t_r36_c60_4;
  wire [7:0] t_r36_c60_5;
  wire [7:0] t_r36_c60_6;
  wire [7:0] t_r36_c60_7;
  wire [7:0] t_r36_c60_8;
  wire [7:0] t_r36_c60_9;
  wire [7:0] t_r36_c60_10;
  wire [7:0] t_r36_c60_11;
  wire [7:0] t_r36_c60_12;
  wire [7:0] t_r36_c61_0;
  wire [7:0] t_r36_c61_1;
  wire [7:0] t_r36_c61_2;
  wire [7:0] t_r36_c61_3;
  wire [7:0] t_r36_c61_4;
  wire [7:0] t_r36_c61_5;
  wire [7:0] t_r36_c61_6;
  wire [7:0] t_r36_c61_7;
  wire [7:0] t_r36_c61_8;
  wire [7:0] t_r36_c61_9;
  wire [7:0] t_r36_c61_10;
  wire [7:0] t_r36_c61_11;
  wire [7:0] t_r36_c61_12;
  wire [7:0] t_r36_c62_0;
  wire [7:0] t_r36_c62_1;
  wire [7:0] t_r36_c62_2;
  wire [7:0] t_r36_c62_3;
  wire [7:0] t_r36_c62_4;
  wire [7:0] t_r36_c62_5;
  wire [7:0] t_r36_c62_6;
  wire [7:0] t_r36_c62_7;
  wire [7:0] t_r36_c62_8;
  wire [7:0] t_r36_c62_9;
  wire [7:0] t_r36_c62_10;
  wire [7:0] t_r36_c62_11;
  wire [7:0] t_r36_c62_12;
  wire [7:0] t_r36_c63_0;
  wire [7:0] t_r36_c63_1;
  wire [7:0] t_r36_c63_2;
  wire [7:0] t_r36_c63_3;
  wire [7:0] t_r36_c63_4;
  wire [7:0] t_r36_c63_5;
  wire [7:0] t_r36_c63_6;
  wire [7:0] t_r36_c63_7;
  wire [7:0] t_r36_c63_8;
  wire [7:0] t_r36_c63_9;
  wire [7:0] t_r36_c63_10;
  wire [7:0] t_r36_c63_11;
  wire [7:0] t_r36_c63_12;
  wire [7:0] t_r36_c64_0;
  wire [7:0] t_r36_c64_1;
  wire [7:0] t_r36_c64_2;
  wire [7:0] t_r36_c64_3;
  wire [7:0] t_r36_c64_4;
  wire [7:0] t_r36_c64_5;
  wire [7:0] t_r36_c64_6;
  wire [7:0] t_r36_c64_7;
  wire [7:0] t_r36_c64_8;
  wire [7:0] t_r36_c64_9;
  wire [7:0] t_r36_c64_10;
  wire [7:0] t_r36_c64_11;
  wire [7:0] t_r36_c64_12;
  wire [7:0] t_r36_c65_0;
  wire [7:0] t_r36_c65_1;
  wire [7:0] t_r36_c65_2;
  wire [7:0] t_r36_c65_3;
  wire [7:0] t_r36_c65_4;
  wire [7:0] t_r36_c65_5;
  wire [7:0] t_r36_c65_6;
  wire [7:0] t_r36_c65_7;
  wire [7:0] t_r36_c65_8;
  wire [7:0] t_r36_c65_9;
  wire [7:0] t_r36_c65_10;
  wire [7:0] t_r36_c65_11;
  wire [7:0] t_r36_c65_12;
  wire [7:0] t_r37_c0_0;
  wire [7:0] t_r37_c0_1;
  wire [7:0] t_r37_c0_2;
  wire [7:0] t_r37_c0_3;
  wire [7:0] t_r37_c0_4;
  wire [7:0] t_r37_c0_5;
  wire [7:0] t_r37_c0_6;
  wire [7:0] t_r37_c0_7;
  wire [7:0] t_r37_c0_8;
  wire [7:0] t_r37_c0_9;
  wire [7:0] t_r37_c0_10;
  wire [7:0] t_r37_c0_11;
  wire [7:0] t_r37_c0_12;
  wire [7:0] t_r37_c1_0;
  wire [7:0] t_r37_c1_1;
  wire [7:0] t_r37_c1_2;
  wire [7:0] t_r37_c1_3;
  wire [7:0] t_r37_c1_4;
  wire [7:0] t_r37_c1_5;
  wire [7:0] t_r37_c1_6;
  wire [7:0] t_r37_c1_7;
  wire [7:0] t_r37_c1_8;
  wire [7:0] t_r37_c1_9;
  wire [7:0] t_r37_c1_10;
  wire [7:0] t_r37_c1_11;
  wire [7:0] t_r37_c1_12;
  wire [7:0] t_r37_c2_0;
  wire [7:0] t_r37_c2_1;
  wire [7:0] t_r37_c2_2;
  wire [7:0] t_r37_c2_3;
  wire [7:0] t_r37_c2_4;
  wire [7:0] t_r37_c2_5;
  wire [7:0] t_r37_c2_6;
  wire [7:0] t_r37_c2_7;
  wire [7:0] t_r37_c2_8;
  wire [7:0] t_r37_c2_9;
  wire [7:0] t_r37_c2_10;
  wire [7:0] t_r37_c2_11;
  wire [7:0] t_r37_c2_12;
  wire [7:0] t_r37_c3_0;
  wire [7:0] t_r37_c3_1;
  wire [7:0] t_r37_c3_2;
  wire [7:0] t_r37_c3_3;
  wire [7:0] t_r37_c3_4;
  wire [7:0] t_r37_c3_5;
  wire [7:0] t_r37_c3_6;
  wire [7:0] t_r37_c3_7;
  wire [7:0] t_r37_c3_8;
  wire [7:0] t_r37_c3_9;
  wire [7:0] t_r37_c3_10;
  wire [7:0] t_r37_c3_11;
  wire [7:0] t_r37_c3_12;
  wire [7:0] t_r37_c4_0;
  wire [7:0] t_r37_c4_1;
  wire [7:0] t_r37_c4_2;
  wire [7:0] t_r37_c4_3;
  wire [7:0] t_r37_c4_4;
  wire [7:0] t_r37_c4_5;
  wire [7:0] t_r37_c4_6;
  wire [7:0] t_r37_c4_7;
  wire [7:0] t_r37_c4_8;
  wire [7:0] t_r37_c4_9;
  wire [7:0] t_r37_c4_10;
  wire [7:0] t_r37_c4_11;
  wire [7:0] t_r37_c4_12;
  wire [7:0] t_r37_c5_0;
  wire [7:0] t_r37_c5_1;
  wire [7:0] t_r37_c5_2;
  wire [7:0] t_r37_c5_3;
  wire [7:0] t_r37_c5_4;
  wire [7:0] t_r37_c5_5;
  wire [7:0] t_r37_c5_6;
  wire [7:0] t_r37_c5_7;
  wire [7:0] t_r37_c5_8;
  wire [7:0] t_r37_c5_9;
  wire [7:0] t_r37_c5_10;
  wire [7:0] t_r37_c5_11;
  wire [7:0] t_r37_c5_12;
  wire [7:0] t_r37_c6_0;
  wire [7:0] t_r37_c6_1;
  wire [7:0] t_r37_c6_2;
  wire [7:0] t_r37_c6_3;
  wire [7:0] t_r37_c6_4;
  wire [7:0] t_r37_c6_5;
  wire [7:0] t_r37_c6_6;
  wire [7:0] t_r37_c6_7;
  wire [7:0] t_r37_c6_8;
  wire [7:0] t_r37_c6_9;
  wire [7:0] t_r37_c6_10;
  wire [7:0] t_r37_c6_11;
  wire [7:0] t_r37_c6_12;
  wire [7:0] t_r37_c7_0;
  wire [7:0] t_r37_c7_1;
  wire [7:0] t_r37_c7_2;
  wire [7:0] t_r37_c7_3;
  wire [7:0] t_r37_c7_4;
  wire [7:0] t_r37_c7_5;
  wire [7:0] t_r37_c7_6;
  wire [7:0] t_r37_c7_7;
  wire [7:0] t_r37_c7_8;
  wire [7:0] t_r37_c7_9;
  wire [7:0] t_r37_c7_10;
  wire [7:0] t_r37_c7_11;
  wire [7:0] t_r37_c7_12;
  wire [7:0] t_r37_c8_0;
  wire [7:0] t_r37_c8_1;
  wire [7:0] t_r37_c8_2;
  wire [7:0] t_r37_c8_3;
  wire [7:0] t_r37_c8_4;
  wire [7:0] t_r37_c8_5;
  wire [7:0] t_r37_c8_6;
  wire [7:0] t_r37_c8_7;
  wire [7:0] t_r37_c8_8;
  wire [7:0] t_r37_c8_9;
  wire [7:0] t_r37_c8_10;
  wire [7:0] t_r37_c8_11;
  wire [7:0] t_r37_c8_12;
  wire [7:0] t_r37_c9_0;
  wire [7:0] t_r37_c9_1;
  wire [7:0] t_r37_c9_2;
  wire [7:0] t_r37_c9_3;
  wire [7:0] t_r37_c9_4;
  wire [7:0] t_r37_c9_5;
  wire [7:0] t_r37_c9_6;
  wire [7:0] t_r37_c9_7;
  wire [7:0] t_r37_c9_8;
  wire [7:0] t_r37_c9_9;
  wire [7:0] t_r37_c9_10;
  wire [7:0] t_r37_c9_11;
  wire [7:0] t_r37_c9_12;
  wire [7:0] t_r37_c10_0;
  wire [7:0] t_r37_c10_1;
  wire [7:0] t_r37_c10_2;
  wire [7:0] t_r37_c10_3;
  wire [7:0] t_r37_c10_4;
  wire [7:0] t_r37_c10_5;
  wire [7:0] t_r37_c10_6;
  wire [7:0] t_r37_c10_7;
  wire [7:0] t_r37_c10_8;
  wire [7:0] t_r37_c10_9;
  wire [7:0] t_r37_c10_10;
  wire [7:0] t_r37_c10_11;
  wire [7:0] t_r37_c10_12;
  wire [7:0] t_r37_c11_0;
  wire [7:0] t_r37_c11_1;
  wire [7:0] t_r37_c11_2;
  wire [7:0] t_r37_c11_3;
  wire [7:0] t_r37_c11_4;
  wire [7:0] t_r37_c11_5;
  wire [7:0] t_r37_c11_6;
  wire [7:0] t_r37_c11_7;
  wire [7:0] t_r37_c11_8;
  wire [7:0] t_r37_c11_9;
  wire [7:0] t_r37_c11_10;
  wire [7:0] t_r37_c11_11;
  wire [7:0] t_r37_c11_12;
  wire [7:0] t_r37_c12_0;
  wire [7:0] t_r37_c12_1;
  wire [7:0] t_r37_c12_2;
  wire [7:0] t_r37_c12_3;
  wire [7:0] t_r37_c12_4;
  wire [7:0] t_r37_c12_5;
  wire [7:0] t_r37_c12_6;
  wire [7:0] t_r37_c12_7;
  wire [7:0] t_r37_c12_8;
  wire [7:0] t_r37_c12_9;
  wire [7:0] t_r37_c12_10;
  wire [7:0] t_r37_c12_11;
  wire [7:0] t_r37_c12_12;
  wire [7:0] t_r37_c13_0;
  wire [7:0] t_r37_c13_1;
  wire [7:0] t_r37_c13_2;
  wire [7:0] t_r37_c13_3;
  wire [7:0] t_r37_c13_4;
  wire [7:0] t_r37_c13_5;
  wire [7:0] t_r37_c13_6;
  wire [7:0] t_r37_c13_7;
  wire [7:0] t_r37_c13_8;
  wire [7:0] t_r37_c13_9;
  wire [7:0] t_r37_c13_10;
  wire [7:0] t_r37_c13_11;
  wire [7:0] t_r37_c13_12;
  wire [7:0] t_r37_c14_0;
  wire [7:0] t_r37_c14_1;
  wire [7:0] t_r37_c14_2;
  wire [7:0] t_r37_c14_3;
  wire [7:0] t_r37_c14_4;
  wire [7:0] t_r37_c14_5;
  wire [7:0] t_r37_c14_6;
  wire [7:0] t_r37_c14_7;
  wire [7:0] t_r37_c14_8;
  wire [7:0] t_r37_c14_9;
  wire [7:0] t_r37_c14_10;
  wire [7:0] t_r37_c14_11;
  wire [7:0] t_r37_c14_12;
  wire [7:0] t_r37_c15_0;
  wire [7:0] t_r37_c15_1;
  wire [7:0] t_r37_c15_2;
  wire [7:0] t_r37_c15_3;
  wire [7:0] t_r37_c15_4;
  wire [7:0] t_r37_c15_5;
  wire [7:0] t_r37_c15_6;
  wire [7:0] t_r37_c15_7;
  wire [7:0] t_r37_c15_8;
  wire [7:0] t_r37_c15_9;
  wire [7:0] t_r37_c15_10;
  wire [7:0] t_r37_c15_11;
  wire [7:0] t_r37_c15_12;
  wire [7:0] t_r37_c16_0;
  wire [7:0] t_r37_c16_1;
  wire [7:0] t_r37_c16_2;
  wire [7:0] t_r37_c16_3;
  wire [7:0] t_r37_c16_4;
  wire [7:0] t_r37_c16_5;
  wire [7:0] t_r37_c16_6;
  wire [7:0] t_r37_c16_7;
  wire [7:0] t_r37_c16_8;
  wire [7:0] t_r37_c16_9;
  wire [7:0] t_r37_c16_10;
  wire [7:0] t_r37_c16_11;
  wire [7:0] t_r37_c16_12;
  wire [7:0] t_r37_c17_0;
  wire [7:0] t_r37_c17_1;
  wire [7:0] t_r37_c17_2;
  wire [7:0] t_r37_c17_3;
  wire [7:0] t_r37_c17_4;
  wire [7:0] t_r37_c17_5;
  wire [7:0] t_r37_c17_6;
  wire [7:0] t_r37_c17_7;
  wire [7:0] t_r37_c17_8;
  wire [7:0] t_r37_c17_9;
  wire [7:0] t_r37_c17_10;
  wire [7:0] t_r37_c17_11;
  wire [7:0] t_r37_c17_12;
  wire [7:0] t_r37_c18_0;
  wire [7:0] t_r37_c18_1;
  wire [7:0] t_r37_c18_2;
  wire [7:0] t_r37_c18_3;
  wire [7:0] t_r37_c18_4;
  wire [7:0] t_r37_c18_5;
  wire [7:0] t_r37_c18_6;
  wire [7:0] t_r37_c18_7;
  wire [7:0] t_r37_c18_8;
  wire [7:0] t_r37_c18_9;
  wire [7:0] t_r37_c18_10;
  wire [7:0] t_r37_c18_11;
  wire [7:0] t_r37_c18_12;
  wire [7:0] t_r37_c19_0;
  wire [7:0] t_r37_c19_1;
  wire [7:0] t_r37_c19_2;
  wire [7:0] t_r37_c19_3;
  wire [7:0] t_r37_c19_4;
  wire [7:0] t_r37_c19_5;
  wire [7:0] t_r37_c19_6;
  wire [7:0] t_r37_c19_7;
  wire [7:0] t_r37_c19_8;
  wire [7:0] t_r37_c19_9;
  wire [7:0] t_r37_c19_10;
  wire [7:0] t_r37_c19_11;
  wire [7:0] t_r37_c19_12;
  wire [7:0] t_r37_c20_0;
  wire [7:0] t_r37_c20_1;
  wire [7:0] t_r37_c20_2;
  wire [7:0] t_r37_c20_3;
  wire [7:0] t_r37_c20_4;
  wire [7:0] t_r37_c20_5;
  wire [7:0] t_r37_c20_6;
  wire [7:0] t_r37_c20_7;
  wire [7:0] t_r37_c20_8;
  wire [7:0] t_r37_c20_9;
  wire [7:0] t_r37_c20_10;
  wire [7:0] t_r37_c20_11;
  wire [7:0] t_r37_c20_12;
  wire [7:0] t_r37_c21_0;
  wire [7:0] t_r37_c21_1;
  wire [7:0] t_r37_c21_2;
  wire [7:0] t_r37_c21_3;
  wire [7:0] t_r37_c21_4;
  wire [7:0] t_r37_c21_5;
  wire [7:0] t_r37_c21_6;
  wire [7:0] t_r37_c21_7;
  wire [7:0] t_r37_c21_8;
  wire [7:0] t_r37_c21_9;
  wire [7:0] t_r37_c21_10;
  wire [7:0] t_r37_c21_11;
  wire [7:0] t_r37_c21_12;
  wire [7:0] t_r37_c22_0;
  wire [7:0] t_r37_c22_1;
  wire [7:0] t_r37_c22_2;
  wire [7:0] t_r37_c22_3;
  wire [7:0] t_r37_c22_4;
  wire [7:0] t_r37_c22_5;
  wire [7:0] t_r37_c22_6;
  wire [7:0] t_r37_c22_7;
  wire [7:0] t_r37_c22_8;
  wire [7:0] t_r37_c22_9;
  wire [7:0] t_r37_c22_10;
  wire [7:0] t_r37_c22_11;
  wire [7:0] t_r37_c22_12;
  wire [7:0] t_r37_c23_0;
  wire [7:0] t_r37_c23_1;
  wire [7:0] t_r37_c23_2;
  wire [7:0] t_r37_c23_3;
  wire [7:0] t_r37_c23_4;
  wire [7:0] t_r37_c23_5;
  wire [7:0] t_r37_c23_6;
  wire [7:0] t_r37_c23_7;
  wire [7:0] t_r37_c23_8;
  wire [7:0] t_r37_c23_9;
  wire [7:0] t_r37_c23_10;
  wire [7:0] t_r37_c23_11;
  wire [7:0] t_r37_c23_12;
  wire [7:0] t_r37_c24_0;
  wire [7:0] t_r37_c24_1;
  wire [7:0] t_r37_c24_2;
  wire [7:0] t_r37_c24_3;
  wire [7:0] t_r37_c24_4;
  wire [7:0] t_r37_c24_5;
  wire [7:0] t_r37_c24_6;
  wire [7:0] t_r37_c24_7;
  wire [7:0] t_r37_c24_8;
  wire [7:0] t_r37_c24_9;
  wire [7:0] t_r37_c24_10;
  wire [7:0] t_r37_c24_11;
  wire [7:0] t_r37_c24_12;
  wire [7:0] t_r37_c25_0;
  wire [7:0] t_r37_c25_1;
  wire [7:0] t_r37_c25_2;
  wire [7:0] t_r37_c25_3;
  wire [7:0] t_r37_c25_4;
  wire [7:0] t_r37_c25_5;
  wire [7:0] t_r37_c25_6;
  wire [7:0] t_r37_c25_7;
  wire [7:0] t_r37_c25_8;
  wire [7:0] t_r37_c25_9;
  wire [7:0] t_r37_c25_10;
  wire [7:0] t_r37_c25_11;
  wire [7:0] t_r37_c25_12;
  wire [7:0] t_r37_c26_0;
  wire [7:0] t_r37_c26_1;
  wire [7:0] t_r37_c26_2;
  wire [7:0] t_r37_c26_3;
  wire [7:0] t_r37_c26_4;
  wire [7:0] t_r37_c26_5;
  wire [7:0] t_r37_c26_6;
  wire [7:0] t_r37_c26_7;
  wire [7:0] t_r37_c26_8;
  wire [7:0] t_r37_c26_9;
  wire [7:0] t_r37_c26_10;
  wire [7:0] t_r37_c26_11;
  wire [7:0] t_r37_c26_12;
  wire [7:0] t_r37_c27_0;
  wire [7:0] t_r37_c27_1;
  wire [7:0] t_r37_c27_2;
  wire [7:0] t_r37_c27_3;
  wire [7:0] t_r37_c27_4;
  wire [7:0] t_r37_c27_5;
  wire [7:0] t_r37_c27_6;
  wire [7:0] t_r37_c27_7;
  wire [7:0] t_r37_c27_8;
  wire [7:0] t_r37_c27_9;
  wire [7:0] t_r37_c27_10;
  wire [7:0] t_r37_c27_11;
  wire [7:0] t_r37_c27_12;
  wire [7:0] t_r37_c28_0;
  wire [7:0] t_r37_c28_1;
  wire [7:0] t_r37_c28_2;
  wire [7:0] t_r37_c28_3;
  wire [7:0] t_r37_c28_4;
  wire [7:0] t_r37_c28_5;
  wire [7:0] t_r37_c28_6;
  wire [7:0] t_r37_c28_7;
  wire [7:0] t_r37_c28_8;
  wire [7:0] t_r37_c28_9;
  wire [7:0] t_r37_c28_10;
  wire [7:0] t_r37_c28_11;
  wire [7:0] t_r37_c28_12;
  wire [7:0] t_r37_c29_0;
  wire [7:0] t_r37_c29_1;
  wire [7:0] t_r37_c29_2;
  wire [7:0] t_r37_c29_3;
  wire [7:0] t_r37_c29_4;
  wire [7:0] t_r37_c29_5;
  wire [7:0] t_r37_c29_6;
  wire [7:0] t_r37_c29_7;
  wire [7:0] t_r37_c29_8;
  wire [7:0] t_r37_c29_9;
  wire [7:0] t_r37_c29_10;
  wire [7:0] t_r37_c29_11;
  wire [7:0] t_r37_c29_12;
  wire [7:0] t_r37_c30_0;
  wire [7:0] t_r37_c30_1;
  wire [7:0] t_r37_c30_2;
  wire [7:0] t_r37_c30_3;
  wire [7:0] t_r37_c30_4;
  wire [7:0] t_r37_c30_5;
  wire [7:0] t_r37_c30_6;
  wire [7:0] t_r37_c30_7;
  wire [7:0] t_r37_c30_8;
  wire [7:0] t_r37_c30_9;
  wire [7:0] t_r37_c30_10;
  wire [7:0] t_r37_c30_11;
  wire [7:0] t_r37_c30_12;
  wire [7:0] t_r37_c31_0;
  wire [7:0] t_r37_c31_1;
  wire [7:0] t_r37_c31_2;
  wire [7:0] t_r37_c31_3;
  wire [7:0] t_r37_c31_4;
  wire [7:0] t_r37_c31_5;
  wire [7:0] t_r37_c31_6;
  wire [7:0] t_r37_c31_7;
  wire [7:0] t_r37_c31_8;
  wire [7:0] t_r37_c31_9;
  wire [7:0] t_r37_c31_10;
  wire [7:0] t_r37_c31_11;
  wire [7:0] t_r37_c31_12;
  wire [7:0] t_r37_c32_0;
  wire [7:0] t_r37_c32_1;
  wire [7:0] t_r37_c32_2;
  wire [7:0] t_r37_c32_3;
  wire [7:0] t_r37_c32_4;
  wire [7:0] t_r37_c32_5;
  wire [7:0] t_r37_c32_6;
  wire [7:0] t_r37_c32_7;
  wire [7:0] t_r37_c32_8;
  wire [7:0] t_r37_c32_9;
  wire [7:0] t_r37_c32_10;
  wire [7:0] t_r37_c32_11;
  wire [7:0] t_r37_c32_12;
  wire [7:0] t_r37_c33_0;
  wire [7:0] t_r37_c33_1;
  wire [7:0] t_r37_c33_2;
  wire [7:0] t_r37_c33_3;
  wire [7:0] t_r37_c33_4;
  wire [7:0] t_r37_c33_5;
  wire [7:0] t_r37_c33_6;
  wire [7:0] t_r37_c33_7;
  wire [7:0] t_r37_c33_8;
  wire [7:0] t_r37_c33_9;
  wire [7:0] t_r37_c33_10;
  wire [7:0] t_r37_c33_11;
  wire [7:0] t_r37_c33_12;
  wire [7:0] t_r37_c34_0;
  wire [7:0] t_r37_c34_1;
  wire [7:0] t_r37_c34_2;
  wire [7:0] t_r37_c34_3;
  wire [7:0] t_r37_c34_4;
  wire [7:0] t_r37_c34_5;
  wire [7:0] t_r37_c34_6;
  wire [7:0] t_r37_c34_7;
  wire [7:0] t_r37_c34_8;
  wire [7:0] t_r37_c34_9;
  wire [7:0] t_r37_c34_10;
  wire [7:0] t_r37_c34_11;
  wire [7:0] t_r37_c34_12;
  wire [7:0] t_r37_c35_0;
  wire [7:0] t_r37_c35_1;
  wire [7:0] t_r37_c35_2;
  wire [7:0] t_r37_c35_3;
  wire [7:0] t_r37_c35_4;
  wire [7:0] t_r37_c35_5;
  wire [7:0] t_r37_c35_6;
  wire [7:0] t_r37_c35_7;
  wire [7:0] t_r37_c35_8;
  wire [7:0] t_r37_c35_9;
  wire [7:0] t_r37_c35_10;
  wire [7:0] t_r37_c35_11;
  wire [7:0] t_r37_c35_12;
  wire [7:0] t_r37_c36_0;
  wire [7:0] t_r37_c36_1;
  wire [7:0] t_r37_c36_2;
  wire [7:0] t_r37_c36_3;
  wire [7:0] t_r37_c36_4;
  wire [7:0] t_r37_c36_5;
  wire [7:0] t_r37_c36_6;
  wire [7:0] t_r37_c36_7;
  wire [7:0] t_r37_c36_8;
  wire [7:0] t_r37_c36_9;
  wire [7:0] t_r37_c36_10;
  wire [7:0] t_r37_c36_11;
  wire [7:0] t_r37_c36_12;
  wire [7:0] t_r37_c37_0;
  wire [7:0] t_r37_c37_1;
  wire [7:0] t_r37_c37_2;
  wire [7:0] t_r37_c37_3;
  wire [7:0] t_r37_c37_4;
  wire [7:0] t_r37_c37_5;
  wire [7:0] t_r37_c37_6;
  wire [7:0] t_r37_c37_7;
  wire [7:0] t_r37_c37_8;
  wire [7:0] t_r37_c37_9;
  wire [7:0] t_r37_c37_10;
  wire [7:0] t_r37_c37_11;
  wire [7:0] t_r37_c37_12;
  wire [7:0] t_r37_c38_0;
  wire [7:0] t_r37_c38_1;
  wire [7:0] t_r37_c38_2;
  wire [7:0] t_r37_c38_3;
  wire [7:0] t_r37_c38_4;
  wire [7:0] t_r37_c38_5;
  wire [7:0] t_r37_c38_6;
  wire [7:0] t_r37_c38_7;
  wire [7:0] t_r37_c38_8;
  wire [7:0] t_r37_c38_9;
  wire [7:0] t_r37_c38_10;
  wire [7:0] t_r37_c38_11;
  wire [7:0] t_r37_c38_12;
  wire [7:0] t_r37_c39_0;
  wire [7:0] t_r37_c39_1;
  wire [7:0] t_r37_c39_2;
  wire [7:0] t_r37_c39_3;
  wire [7:0] t_r37_c39_4;
  wire [7:0] t_r37_c39_5;
  wire [7:0] t_r37_c39_6;
  wire [7:0] t_r37_c39_7;
  wire [7:0] t_r37_c39_8;
  wire [7:0] t_r37_c39_9;
  wire [7:0] t_r37_c39_10;
  wire [7:0] t_r37_c39_11;
  wire [7:0] t_r37_c39_12;
  wire [7:0] t_r37_c40_0;
  wire [7:0] t_r37_c40_1;
  wire [7:0] t_r37_c40_2;
  wire [7:0] t_r37_c40_3;
  wire [7:0] t_r37_c40_4;
  wire [7:0] t_r37_c40_5;
  wire [7:0] t_r37_c40_6;
  wire [7:0] t_r37_c40_7;
  wire [7:0] t_r37_c40_8;
  wire [7:0] t_r37_c40_9;
  wire [7:0] t_r37_c40_10;
  wire [7:0] t_r37_c40_11;
  wire [7:0] t_r37_c40_12;
  wire [7:0] t_r37_c41_0;
  wire [7:0] t_r37_c41_1;
  wire [7:0] t_r37_c41_2;
  wire [7:0] t_r37_c41_3;
  wire [7:0] t_r37_c41_4;
  wire [7:0] t_r37_c41_5;
  wire [7:0] t_r37_c41_6;
  wire [7:0] t_r37_c41_7;
  wire [7:0] t_r37_c41_8;
  wire [7:0] t_r37_c41_9;
  wire [7:0] t_r37_c41_10;
  wire [7:0] t_r37_c41_11;
  wire [7:0] t_r37_c41_12;
  wire [7:0] t_r37_c42_0;
  wire [7:0] t_r37_c42_1;
  wire [7:0] t_r37_c42_2;
  wire [7:0] t_r37_c42_3;
  wire [7:0] t_r37_c42_4;
  wire [7:0] t_r37_c42_5;
  wire [7:0] t_r37_c42_6;
  wire [7:0] t_r37_c42_7;
  wire [7:0] t_r37_c42_8;
  wire [7:0] t_r37_c42_9;
  wire [7:0] t_r37_c42_10;
  wire [7:0] t_r37_c42_11;
  wire [7:0] t_r37_c42_12;
  wire [7:0] t_r37_c43_0;
  wire [7:0] t_r37_c43_1;
  wire [7:0] t_r37_c43_2;
  wire [7:0] t_r37_c43_3;
  wire [7:0] t_r37_c43_4;
  wire [7:0] t_r37_c43_5;
  wire [7:0] t_r37_c43_6;
  wire [7:0] t_r37_c43_7;
  wire [7:0] t_r37_c43_8;
  wire [7:0] t_r37_c43_9;
  wire [7:0] t_r37_c43_10;
  wire [7:0] t_r37_c43_11;
  wire [7:0] t_r37_c43_12;
  wire [7:0] t_r37_c44_0;
  wire [7:0] t_r37_c44_1;
  wire [7:0] t_r37_c44_2;
  wire [7:0] t_r37_c44_3;
  wire [7:0] t_r37_c44_4;
  wire [7:0] t_r37_c44_5;
  wire [7:0] t_r37_c44_6;
  wire [7:0] t_r37_c44_7;
  wire [7:0] t_r37_c44_8;
  wire [7:0] t_r37_c44_9;
  wire [7:0] t_r37_c44_10;
  wire [7:0] t_r37_c44_11;
  wire [7:0] t_r37_c44_12;
  wire [7:0] t_r37_c45_0;
  wire [7:0] t_r37_c45_1;
  wire [7:0] t_r37_c45_2;
  wire [7:0] t_r37_c45_3;
  wire [7:0] t_r37_c45_4;
  wire [7:0] t_r37_c45_5;
  wire [7:0] t_r37_c45_6;
  wire [7:0] t_r37_c45_7;
  wire [7:0] t_r37_c45_8;
  wire [7:0] t_r37_c45_9;
  wire [7:0] t_r37_c45_10;
  wire [7:0] t_r37_c45_11;
  wire [7:0] t_r37_c45_12;
  wire [7:0] t_r37_c46_0;
  wire [7:0] t_r37_c46_1;
  wire [7:0] t_r37_c46_2;
  wire [7:0] t_r37_c46_3;
  wire [7:0] t_r37_c46_4;
  wire [7:0] t_r37_c46_5;
  wire [7:0] t_r37_c46_6;
  wire [7:0] t_r37_c46_7;
  wire [7:0] t_r37_c46_8;
  wire [7:0] t_r37_c46_9;
  wire [7:0] t_r37_c46_10;
  wire [7:0] t_r37_c46_11;
  wire [7:0] t_r37_c46_12;
  wire [7:0] t_r37_c47_0;
  wire [7:0] t_r37_c47_1;
  wire [7:0] t_r37_c47_2;
  wire [7:0] t_r37_c47_3;
  wire [7:0] t_r37_c47_4;
  wire [7:0] t_r37_c47_5;
  wire [7:0] t_r37_c47_6;
  wire [7:0] t_r37_c47_7;
  wire [7:0] t_r37_c47_8;
  wire [7:0] t_r37_c47_9;
  wire [7:0] t_r37_c47_10;
  wire [7:0] t_r37_c47_11;
  wire [7:0] t_r37_c47_12;
  wire [7:0] t_r37_c48_0;
  wire [7:0] t_r37_c48_1;
  wire [7:0] t_r37_c48_2;
  wire [7:0] t_r37_c48_3;
  wire [7:0] t_r37_c48_4;
  wire [7:0] t_r37_c48_5;
  wire [7:0] t_r37_c48_6;
  wire [7:0] t_r37_c48_7;
  wire [7:0] t_r37_c48_8;
  wire [7:0] t_r37_c48_9;
  wire [7:0] t_r37_c48_10;
  wire [7:0] t_r37_c48_11;
  wire [7:0] t_r37_c48_12;
  wire [7:0] t_r37_c49_0;
  wire [7:0] t_r37_c49_1;
  wire [7:0] t_r37_c49_2;
  wire [7:0] t_r37_c49_3;
  wire [7:0] t_r37_c49_4;
  wire [7:0] t_r37_c49_5;
  wire [7:0] t_r37_c49_6;
  wire [7:0] t_r37_c49_7;
  wire [7:0] t_r37_c49_8;
  wire [7:0] t_r37_c49_9;
  wire [7:0] t_r37_c49_10;
  wire [7:0] t_r37_c49_11;
  wire [7:0] t_r37_c49_12;
  wire [7:0] t_r37_c50_0;
  wire [7:0] t_r37_c50_1;
  wire [7:0] t_r37_c50_2;
  wire [7:0] t_r37_c50_3;
  wire [7:0] t_r37_c50_4;
  wire [7:0] t_r37_c50_5;
  wire [7:0] t_r37_c50_6;
  wire [7:0] t_r37_c50_7;
  wire [7:0] t_r37_c50_8;
  wire [7:0] t_r37_c50_9;
  wire [7:0] t_r37_c50_10;
  wire [7:0] t_r37_c50_11;
  wire [7:0] t_r37_c50_12;
  wire [7:0] t_r37_c51_0;
  wire [7:0] t_r37_c51_1;
  wire [7:0] t_r37_c51_2;
  wire [7:0] t_r37_c51_3;
  wire [7:0] t_r37_c51_4;
  wire [7:0] t_r37_c51_5;
  wire [7:0] t_r37_c51_6;
  wire [7:0] t_r37_c51_7;
  wire [7:0] t_r37_c51_8;
  wire [7:0] t_r37_c51_9;
  wire [7:0] t_r37_c51_10;
  wire [7:0] t_r37_c51_11;
  wire [7:0] t_r37_c51_12;
  wire [7:0] t_r37_c52_0;
  wire [7:0] t_r37_c52_1;
  wire [7:0] t_r37_c52_2;
  wire [7:0] t_r37_c52_3;
  wire [7:0] t_r37_c52_4;
  wire [7:0] t_r37_c52_5;
  wire [7:0] t_r37_c52_6;
  wire [7:0] t_r37_c52_7;
  wire [7:0] t_r37_c52_8;
  wire [7:0] t_r37_c52_9;
  wire [7:0] t_r37_c52_10;
  wire [7:0] t_r37_c52_11;
  wire [7:0] t_r37_c52_12;
  wire [7:0] t_r37_c53_0;
  wire [7:0] t_r37_c53_1;
  wire [7:0] t_r37_c53_2;
  wire [7:0] t_r37_c53_3;
  wire [7:0] t_r37_c53_4;
  wire [7:0] t_r37_c53_5;
  wire [7:0] t_r37_c53_6;
  wire [7:0] t_r37_c53_7;
  wire [7:0] t_r37_c53_8;
  wire [7:0] t_r37_c53_9;
  wire [7:0] t_r37_c53_10;
  wire [7:0] t_r37_c53_11;
  wire [7:0] t_r37_c53_12;
  wire [7:0] t_r37_c54_0;
  wire [7:0] t_r37_c54_1;
  wire [7:0] t_r37_c54_2;
  wire [7:0] t_r37_c54_3;
  wire [7:0] t_r37_c54_4;
  wire [7:0] t_r37_c54_5;
  wire [7:0] t_r37_c54_6;
  wire [7:0] t_r37_c54_7;
  wire [7:0] t_r37_c54_8;
  wire [7:0] t_r37_c54_9;
  wire [7:0] t_r37_c54_10;
  wire [7:0] t_r37_c54_11;
  wire [7:0] t_r37_c54_12;
  wire [7:0] t_r37_c55_0;
  wire [7:0] t_r37_c55_1;
  wire [7:0] t_r37_c55_2;
  wire [7:0] t_r37_c55_3;
  wire [7:0] t_r37_c55_4;
  wire [7:0] t_r37_c55_5;
  wire [7:0] t_r37_c55_6;
  wire [7:0] t_r37_c55_7;
  wire [7:0] t_r37_c55_8;
  wire [7:0] t_r37_c55_9;
  wire [7:0] t_r37_c55_10;
  wire [7:0] t_r37_c55_11;
  wire [7:0] t_r37_c55_12;
  wire [7:0] t_r37_c56_0;
  wire [7:0] t_r37_c56_1;
  wire [7:0] t_r37_c56_2;
  wire [7:0] t_r37_c56_3;
  wire [7:0] t_r37_c56_4;
  wire [7:0] t_r37_c56_5;
  wire [7:0] t_r37_c56_6;
  wire [7:0] t_r37_c56_7;
  wire [7:0] t_r37_c56_8;
  wire [7:0] t_r37_c56_9;
  wire [7:0] t_r37_c56_10;
  wire [7:0] t_r37_c56_11;
  wire [7:0] t_r37_c56_12;
  wire [7:0] t_r37_c57_0;
  wire [7:0] t_r37_c57_1;
  wire [7:0] t_r37_c57_2;
  wire [7:0] t_r37_c57_3;
  wire [7:0] t_r37_c57_4;
  wire [7:0] t_r37_c57_5;
  wire [7:0] t_r37_c57_6;
  wire [7:0] t_r37_c57_7;
  wire [7:0] t_r37_c57_8;
  wire [7:0] t_r37_c57_9;
  wire [7:0] t_r37_c57_10;
  wire [7:0] t_r37_c57_11;
  wire [7:0] t_r37_c57_12;
  wire [7:0] t_r37_c58_0;
  wire [7:0] t_r37_c58_1;
  wire [7:0] t_r37_c58_2;
  wire [7:0] t_r37_c58_3;
  wire [7:0] t_r37_c58_4;
  wire [7:0] t_r37_c58_5;
  wire [7:0] t_r37_c58_6;
  wire [7:0] t_r37_c58_7;
  wire [7:0] t_r37_c58_8;
  wire [7:0] t_r37_c58_9;
  wire [7:0] t_r37_c58_10;
  wire [7:0] t_r37_c58_11;
  wire [7:0] t_r37_c58_12;
  wire [7:0] t_r37_c59_0;
  wire [7:0] t_r37_c59_1;
  wire [7:0] t_r37_c59_2;
  wire [7:0] t_r37_c59_3;
  wire [7:0] t_r37_c59_4;
  wire [7:0] t_r37_c59_5;
  wire [7:0] t_r37_c59_6;
  wire [7:0] t_r37_c59_7;
  wire [7:0] t_r37_c59_8;
  wire [7:0] t_r37_c59_9;
  wire [7:0] t_r37_c59_10;
  wire [7:0] t_r37_c59_11;
  wire [7:0] t_r37_c59_12;
  wire [7:0] t_r37_c60_0;
  wire [7:0] t_r37_c60_1;
  wire [7:0] t_r37_c60_2;
  wire [7:0] t_r37_c60_3;
  wire [7:0] t_r37_c60_4;
  wire [7:0] t_r37_c60_5;
  wire [7:0] t_r37_c60_6;
  wire [7:0] t_r37_c60_7;
  wire [7:0] t_r37_c60_8;
  wire [7:0] t_r37_c60_9;
  wire [7:0] t_r37_c60_10;
  wire [7:0] t_r37_c60_11;
  wire [7:0] t_r37_c60_12;
  wire [7:0] t_r37_c61_0;
  wire [7:0] t_r37_c61_1;
  wire [7:0] t_r37_c61_2;
  wire [7:0] t_r37_c61_3;
  wire [7:0] t_r37_c61_4;
  wire [7:0] t_r37_c61_5;
  wire [7:0] t_r37_c61_6;
  wire [7:0] t_r37_c61_7;
  wire [7:0] t_r37_c61_8;
  wire [7:0] t_r37_c61_9;
  wire [7:0] t_r37_c61_10;
  wire [7:0] t_r37_c61_11;
  wire [7:0] t_r37_c61_12;
  wire [7:0] t_r37_c62_0;
  wire [7:0] t_r37_c62_1;
  wire [7:0] t_r37_c62_2;
  wire [7:0] t_r37_c62_3;
  wire [7:0] t_r37_c62_4;
  wire [7:0] t_r37_c62_5;
  wire [7:0] t_r37_c62_6;
  wire [7:0] t_r37_c62_7;
  wire [7:0] t_r37_c62_8;
  wire [7:0] t_r37_c62_9;
  wire [7:0] t_r37_c62_10;
  wire [7:0] t_r37_c62_11;
  wire [7:0] t_r37_c62_12;
  wire [7:0] t_r37_c63_0;
  wire [7:0] t_r37_c63_1;
  wire [7:0] t_r37_c63_2;
  wire [7:0] t_r37_c63_3;
  wire [7:0] t_r37_c63_4;
  wire [7:0] t_r37_c63_5;
  wire [7:0] t_r37_c63_6;
  wire [7:0] t_r37_c63_7;
  wire [7:0] t_r37_c63_8;
  wire [7:0] t_r37_c63_9;
  wire [7:0] t_r37_c63_10;
  wire [7:0] t_r37_c63_11;
  wire [7:0] t_r37_c63_12;
  wire [7:0] t_r37_c64_0;
  wire [7:0] t_r37_c64_1;
  wire [7:0] t_r37_c64_2;
  wire [7:0] t_r37_c64_3;
  wire [7:0] t_r37_c64_4;
  wire [7:0] t_r37_c64_5;
  wire [7:0] t_r37_c64_6;
  wire [7:0] t_r37_c64_7;
  wire [7:0] t_r37_c64_8;
  wire [7:0] t_r37_c64_9;
  wire [7:0] t_r37_c64_10;
  wire [7:0] t_r37_c64_11;
  wire [7:0] t_r37_c64_12;
  wire [7:0] t_r37_c65_0;
  wire [7:0] t_r37_c65_1;
  wire [7:0] t_r37_c65_2;
  wire [7:0] t_r37_c65_3;
  wire [7:0] t_r37_c65_4;
  wire [7:0] t_r37_c65_5;
  wire [7:0] t_r37_c65_6;
  wire [7:0] t_r37_c65_7;
  wire [7:0] t_r37_c65_8;
  wire [7:0] t_r37_c65_9;
  wire [7:0] t_r37_c65_10;
  wire [7:0] t_r37_c65_11;
  wire [7:0] t_r37_c65_12;
  wire [7:0] t_r38_c0_0;
  wire [7:0] t_r38_c0_1;
  wire [7:0] t_r38_c0_2;
  wire [7:0] t_r38_c0_3;
  wire [7:0] t_r38_c0_4;
  wire [7:0] t_r38_c0_5;
  wire [7:0] t_r38_c0_6;
  wire [7:0] t_r38_c0_7;
  wire [7:0] t_r38_c0_8;
  wire [7:0] t_r38_c0_9;
  wire [7:0] t_r38_c0_10;
  wire [7:0] t_r38_c0_11;
  wire [7:0] t_r38_c0_12;
  wire [7:0] t_r38_c1_0;
  wire [7:0] t_r38_c1_1;
  wire [7:0] t_r38_c1_2;
  wire [7:0] t_r38_c1_3;
  wire [7:0] t_r38_c1_4;
  wire [7:0] t_r38_c1_5;
  wire [7:0] t_r38_c1_6;
  wire [7:0] t_r38_c1_7;
  wire [7:0] t_r38_c1_8;
  wire [7:0] t_r38_c1_9;
  wire [7:0] t_r38_c1_10;
  wire [7:0] t_r38_c1_11;
  wire [7:0] t_r38_c1_12;
  wire [7:0] t_r38_c2_0;
  wire [7:0] t_r38_c2_1;
  wire [7:0] t_r38_c2_2;
  wire [7:0] t_r38_c2_3;
  wire [7:0] t_r38_c2_4;
  wire [7:0] t_r38_c2_5;
  wire [7:0] t_r38_c2_6;
  wire [7:0] t_r38_c2_7;
  wire [7:0] t_r38_c2_8;
  wire [7:0] t_r38_c2_9;
  wire [7:0] t_r38_c2_10;
  wire [7:0] t_r38_c2_11;
  wire [7:0] t_r38_c2_12;
  wire [7:0] t_r38_c3_0;
  wire [7:0] t_r38_c3_1;
  wire [7:0] t_r38_c3_2;
  wire [7:0] t_r38_c3_3;
  wire [7:0] t_r38_c3_4;
  wire [7:0] t_r38_c3_5;
  wire [7:0] t_r38_c3_6;
  wire [7:0] t_r38_c3_7;
  wire [7:0] t_r38_c3_8;
  wire [7:0] t_r38_c3_9;
  wire [7:0] t_r38_c3_10;
  wire [7:0] t_r38_c3_11;
  wire [7:0] t_r38_c3_12;
  wire [7:0] t_r38_c4_0;
  wire [7:0] t_r38_c4_1;
  wire [7:0] t_r38_c4_2;
  wire [7:0] t_r38_c4_3;
  wire [7:0] t_r38_c4_4;
  wire [7:0] t_r38_c4_5;
  wire [7:0] t_r38_c4_6;
  wire [7:0] t_r38_c4_7;
  wire [7:0] t_r38_c4_8;
  wire [7:0] t_r38_c4_9;
  wire [7:0] t_r38_c4_10;
  wire [7:0] t_r38_c4_11;
  wire [7:0] t_r38_c4_12;
  wire [7:0] t_r38_c5_0;
  wire [7:0] t_r38_c5_1;
  wire [7:0] t_r38_c5_2;
  wire [7:0] t_r38_c5_3;
  wire [7:0] t_r38_c5_4;
  wire [7:0] t_r38_c5_5;
  wire [7:0] t_r38_c5_6;
  wire [7:0] t_r38_c5_7;
  wire [7:0] t_r38_c5_8;
  wire [7:0] t_r38_c5_9;
  wire [7:0] t_r38_c5_10;
  wire [7:0] t_r38_c5_11;
  wire [7:0] t_r38_c5_12;
  wire [7:0] t_r38_c6_0;
  wire [7:0] t_r38_c6_1;
  wire [7:0] t_r38_c6_2;
  wire [7:0] t_r38_c6_3;
  wire [7:0] t_r38_c6_4;
  wire [7:0] t_r38_c6_5;
  wire [7:0] t_r38_c6_6;
  wire [7:0] t_r38_c6_7;
  wire [7:0] t_r38_c6_8;
  wire [7:0] t_r38_c6_9;
  wire [7:0] t_r38_c6_10;
  wire [7:0] t_r38_c6_11;
  wire [7:0] t_r38_c6_12;
  wire [7:0] t_r38_c7_0;
  wire [7:0] t_r38_c7_1;
  wire [7:0] t_r38_c7_2;
  wire [7:0] t_r38_c7_3;
  wire [7:0] t_r38_c7_4;
  wire [7:0] t_r38_c7_5;
  wire [7:0] t_r38_c7_6;
  wire [7:0] t_r38_c7_7;
  wire [7:0] t_r38_c7_8;
  wire [7:0] t_r38_c7_9;
  wire [7:0] t_r38_c7_10;
  wire [7:0] t_r38_c7_11;
  wire [7:0] t_r38_c7_12;
  wire [7:0] t_r38_c8_0;
  wire [7:0] t_r38_c8_1;
  wire [7:0] t_r38_c8_2;
  wire [7:0] t_r38_c8_3;
  wire [7:0] t_r38_c8_4;
  wire [7:0] t_r38_c8_5;
  wire [7:0] t_r38_c8_6;
  wire [7:0] t_r38_c8_7;
  wire [7:0] t_r38_c8_8;
  wire [7:0] t_r38_c8_9;
  wire [7:0] t_r38_c8_10;
  wire [7:0] t_r38_c8_11;
  wire [7:0] t_r38_c8_12;
  wire [7:0] t_r38_c9_0;
  wire [7:0] t_r38_c9_1;
  wire [7:0] t_r38_c9_2;
  wire [7:0] t_r38_c9_3;
  wire [7:0] t_r38_c9_4;
  wire [7:0] t_r38_c9_5;
  wire [7:0] t_r38_c9_6;
  wire [7:0] t_r38_c9_7;
  wire [7:0] t_r38_c9_8;
  wire [7:0] t_r38_c9_9;
  wire [7:0] t_r38_c9_10;
  wire [7:0] t_r38_c9_11;
  wire [7:0] t_r38_c9_12;
  wire [7:0] t_r38_c10_0;
  wire [7:0] t_r38_c10_1;
  wire [7:0] t_r38_c10_2;
  wire [7:0] t_r38_c10_3;
  wire [7:0] t_r38_c10_4;
  wire [7:0] t_r38_c10_5;
  wire [7:0] t_r38_c10_6;
  wire [7:0] t_r38_c10_7;
  wire [7:0] t_r38_c10_8;
  wire [7:0] t_r38_c10_9;
  wire [7:0] t_r38_c10_10;
  wire [7:0] t_r38_c10_11;
  wire [7:0] t_r38_c10_12;
  wire [7:0] t_r38_c11_0;
  wire [7:0] t_r38_c11_1;
  wire [7:0] t_r38_c11_2;
  wire [7:0] t_r38_c11_3;
  wire [7:0] t_r38_c11_4;
  wire [7:0] t_r38_c11_5;
  wire [7:0] t_r38_c11_6;
  wire [7:0] t_r38_c11_7;
  wire [7:0] t_r38_c11_8;
  wire [7:0] t_r38_c11_9;
  wire [7:0] t_r38_c11_10;
  wire [7:0] t_r38_c11_11;
  wire [7:0] t_r38_c11_12;
  wire [7:0] t_r38_c12_0;
  wire [7:0] t_r38_c12_1;
  wire [7:0] t_r38_c12_2;
  wire [7:0] t_r38_c12_3;
  wire [7:0] t_r38_c12_4;
  wire [7:0] t_r38_c12_5;
  wire [7:0] t_r38_c12_6;
  wire [7:0] t_r38_c12_7;
  wire [7:0] t_r38_c12_8;
  wire [7:0] t_r38_c12_9;
  wire [7:0] t_r38_c12_10;
  wire [7:0] t_r38_c12_11;
  wire [7:0] t_r38_c12_12;
  wire [7:0] t_r38_c13_0;
  wire [7:0] t_r38_c13_1;
  wire [7:0] t_r38_c13_2;
  wire [7:0] t_r38_c13_3;
  wire [7:0] t_r38_c13_4;
  wire [7:0] t_r38_c13_5;
  wire [7:0] t_r38_c13_6;
  wire [7:0] t_r38_c13_7;
  wire [7:0] t_r38_c13_8;
  wire [7:0] t_r38_c13_9;
  wire [7:0] t_r38_c13_10;
  wire [7:0] t_r38_c13_11;
  wire [7:0] t_r38_c13_12;
  wire [7:0] t_r38_c14_0;
  wire [7:0] t_r38_c14_1;
  wire [7:0] t_r38_c14_2;
  wire [7:0] t_r38_c14_3;
  wire [7:0] t_r38_c14_4;
  wire [7:0] t_r38_c14_5;
  wire [7:0] t_r38_c14_6;
  wire [7:0] t_r38_c14_7;
  wire [7:0] t_r38_c14_8;
  wire [7:0] t_r38_c14_9;
  wire [7:0] t_r38_c14_10;
  wire [7:0] t_r38_c14_11;
  wire [7:0] t_r38_c14_12;
  wire [7:0] t_r38_c15_0;
  wire [7:0] t_r38_c15_1;
  wire [7:0] t_r38_c15_2;
  wire [7:0] t_r38_c15_3;
  wire [7:0] t_r38_c15_4;
  wire [7:0] t_r38_c15_5;
  wire [7:0] t_r38_c15_6;
  wire [7:0] t_r38_c15_7;
  wire [7:0] t_r38_c15_8;
  wire [7:0] t_r38_c15_9;
  wire [7:0] t_r38_c15_10;
  wire [7:0] t_r38_c15_11;
  wire [7:0] t_r38_c15_12;
  wire [7:0] t_r38_c16_0;
  wire [7:0] t_r38_c16_1;
  wire [7:0] t_r38_c16_2;
  wire [7:0] t_r38_c16_3;
  wire [7:0] t_r38_c16_4;
  wire [7:0] t_r38_c16_5;
  wire [7:0] t_r38_c16_6;
  wire [7:0] t_r38_c16_7;
  wire [7:0] t_r38_c16_8;
  wire [7:0] t_r38_c16_9;
  wire [7:0] t_r38_c16_10;
  wire [7:0] t_r38_c16_11;
  wire [7:0] t_r38_c16_12;
  wire [7:0] t_r38_c17_0;
  wire [7:0] t_r38_c17_1;
  wire [7:0] t_r38_c17_2;
  wire [7:0] t_r38_c17_3;
  wire [7:0] t_r38_c17_4;
  wire [7:0] t_r38_c17_5;
  wire [7:0] t_r38_c17_6;
  wire [7:0] t_r38_c17_7;
  wire [7:0] t_r38_c17_8;
  wire [7:0] t_r38_c17_9;
  wire [7:0] t_r38_c17_10;
  wire [7:0] t_r38_c17_11;
  wire [7:0] t_r38_c17_12;
  wire [7:0] t_r38_c18_0;
  wire [7:0] t_r38_c18_1;
  wire [7:0] t_r38_c18_2;
  wire [7:0] t_r38_c18_3;
  wire [7:0] t_r38_c18_4;
  wire [7:0] t_r38_c18_5;
  wire [7:0] t_r38_c18_6;
  wire [7:0] t_r38_c18_7;
  wire [7:0] t_r38_c18_8;
  wire [7:0] t_r38_c18_9;
  wire [7:0] t_r38_c18_10;
  wire [7:0] t_r38_c18_11;
  wire [7:0] t_r38_c18_12;
  wire [7:0] t_r38_c19_0;
  wire [7:0] t_r38_c19_1;
  wire [7:0] t_r38_c19_2;
  wire [7:0] t_r38_c19_3;
  wire [7:0] t_r38_c19_4;
  wire [7:0] t_r38_c19_5;
  wire [7:0] t_r38_c19_6;
  wire [7:0] t_r38_c19_7;
  wire [7:0] t_r38_c19_8;
  wire [7:0] t_r38_c19_9;
  wire [7:0] t_r38_c19_10;
  wire [7:0] t_r38_c19_11;
  wire [7:0] t_r38_c19_12;
  wire [7:0] t_r38_c20_0;
  wire [7:0] t_r38_c20_1;
  wire [7:0] t_r38_c20_2;
  wire [7:0] t_r38_c20_3;
  wire [7:0] t_r38_c20_4;
  wire [7:0] t_r38_c20_5;
  wire [7:0] t_r38_c20_6;
  wire [7:0] t_r38_c20_7;
  wire [7:0] t_r38_c20_8;
  wire [7:0] t_r38_c20_9;
  wire [7:0] t_r38_c20_10;
  wire [7:0] t_r38_c20_11;
  wire [7:0] t_r38_c20_12;
  wire [7:0] t_r38_c21_0;
  wire [7:0] t_r38_c21_1;
  wire [7:0] t_r38_c21_2;
  wire [7:0] t_r38_c21_3;
  wire [7:0] t_r38_c21_4;
  wire [7:0] t_r38_c21_5;
  wire [7:0] t_r38_c21_6;
  wire [7:0] t_r38_c21_7;
  wire [7:0] t_r38_c21_8;
  wire [7:0] t_r38_c21_9;
  wire [7:0] t_r38_c21_10;
  wire [7:0] t_r38_c21_11;
  wire [7:0] t_r38_c21_12;
  wire [7:0] t_r38_c22_0;
  wire [7:0] t_r38_c22_1;
  wire [7:0] t_r38_c22_2;
  wire [7:0] t_r38_c22_3;
  wire [7:0] t_r38_c22_4;
  wire [7:0] t_r38_c22_5;
  wire [7:0] t_r38_c22_6;
  wire [7:0] t_r38_c22_7;
  wire [7:0] t_r38_c22_8;
  wire [7:0] t_r38_c22_9;
  wire [7:0] t_r38_c22_10;
  wire [7:0] t_r38_c22_11;
  wire [7:0] t_r38_c22_12;
  wire [7:0] t_r38_c23_0;
  wire [7:0] t_r38_c23_1;
  wire [7:0] t_r38_c23_2;
  wire [7:0] t_r38_c23_3;
  wire [7:0] t_r38_c23_4;
  wire [7:0] t_r38_c23_5;
  wire [7:0] t_r38_c23_6;
  wire [7:0] t_r38_c23_7;
  wire [7:0] t_r38_c23_8;
  wire [7:0] t_r38_c23_9;
  wire [7:0] t_r38_c23_10;
  wire [7:0] t_r38_c23_11;
  wire [7:0] t_r38_c23_12;
  wire [7:0] t_r38_c24_0;
  wire [7:0] t_r38_c24_1;
  wire [7:0] t_r38_c24_2;
  wire [7:0] t_r38_c24_3;
  wire [7:0] t_r38_c24_4;
  wire [7:0] t_r38_c24_5;
  wire [7:0] t_r38_c24_6;
  wire [7:0] t_r38_c24_7;
  wire [7:0] t_r38_c24_8;
  wire [7:0] t_r38_c24_9;
  wire [7:0] t_r38_c24_10;
  wire [7:0] t_r38_c24_11;
  wire [7:0] t_r38_c24_12;
  wire [7:0] t_r38_c25_0;
  wire [7:0] t_r38_c25_1;
  wire [7:0] t_r38_c25_2;
  wire [7:0] t_r38_c25_3;
  wire [7:0] t_r38_c25_4;
  wire [7:0] t_r38_c25_5;
  wire [7:0] t_r38_c25_6;
  wire [7:0] t_r38_c25_7;
  wire [7:0] t_r38_c25_8;
  wire [7:0] t_r38_c25_9;
  wire [7:0] t_r38_c25_10;
  wire [7:0] t_r38_c25_11;
  wire [7:0] t_r38_c25_12;
  wire [7:0] t_r38_c26_0;
  wire [7:0] t_r38_c26_1;
  wire [7:0] t_r38_c26_2;
  wire [7:0] t_r38_c26_3;
  wire [7:0] t_r38_c26_4;
  wire [7:0] t_r38_c26_5;
  wire [7:0] t_r38_c26_6;
  wire [7:0] t_r38_c26_7;
  wire [7:0] t_r38_c26_8;
  wire [7:0] t_r38_c26_9;
  wire [7:0] t_r38_c26_10;
  wire [7:0] t_r38_c26_11;
  wire [7:0] t_r38_c26_12;
  wire [7:0] t_r38_c27_0;
  wire [7:0] t_r38_c27_1;
  wire [7:0] t_r38_c27_2;
  wire [7:0] t_r38_c27_3;
  wire [7:0] t_r38_c27_4;
  wire [7:0] t_r38_c27_5;
  wire [7:0] t_r38_c27_6;
  wire [7:0] t_r38_c27_7;
  wire [7:0] t_r38_c27_8;
  wire [7:0] t_r38_c27_9;
  wire [7:0] t_r38_c27_10;
  wire [7:0] t_r38_c27_11;
  wire [7:0] t_r38_c27_12;
  wire [7:0] t_r38_c28_0;
  wire [7:0] t_r38_c28_1;
  wire [7:0] t_r38_c28_2;
  wire [7:0] t_r38_c28_3;
  wire [7:0] t_r38_c28_4;
  wire [7:0] t_r38_c28_5;
  wire [7:0] t_r38_c28_6;
  wire [7:0] t_r38_c28_7;
  wire [7:0] t_r38_c28_8;
  wire [7:0] t_r38_c28_9;
  wire [7:0] t_r38_c28_10;
  wire [7:0] t_r38_c28_11;
  wire [7:0] t_r38_c28_12;
  wire [7:0] t_r38_c29_0;
  wire [7:0] t_r38_c29_1;
  wire [7:0] t_r38_c29_2;
  wire [7:0] t_r38_c29_3;
  wire [7:0] t_r38_c29_4;
  wire [7:0] t_r38_c29_5;
  wire [7:0] t_r38_c29_6;
  wire [7:0] t_r38_c29_7;
  wire [7:0] t_r38_c29_8;
  wire [7:0] t_r38_c29_9;
  wire [7:0] t_r38_c29_10;
  wire [7:0] t_r38_c29_11;
  wire [7:0] t_r38_c29_12;
  wire [7:0] t_r38_c30_0;
  wire [7:0] t_r38_c30_1;
  wire [7:0] t_r38_c30_2;
  wire [7:0] t_r38_c30_3;
  wire [7:0] t_r38_c30_4;
  wire [7:0] t_r38_c30_5;
  wire [7:0] t_r38_c30_6;
  wire [7:0] t_r38_c30_7;
  wire [7:0] t_r38_c30_8;
  wire [7:0] t_r38_c30_9;
  wire [7:0] t_r38_c30_10;
  wire [7:0] t_r38_c30_11;
  wire [7:0] t_r38_c30_12;
  wire [7:0] t_r38_c31_0;
  wire [7:0] t_r38_c31_1;
  wire [7:0] t_r38_c31_2;
  wire [7:0] t_r38_c31_3;
  wire [7:0] t_r38_c31_4;
  wire [7:0] t_r38_c31_5;
  wire [7:0] t_r38_c31_6;
  wire [7:0] t_r38_c31_7;
  wire [7:0] t_r38_c31_8;
  wire [7:0] t_r38_c31_9;
  wire [7:0] t_r38_c31_10;
  wire [7:0] t_r38_c31_11;
  wire [7:0] t_r38_c31_12;
  wire [7:0] t_r38_c32_0;
  wire [7:0] t_r38_c32_1;
  wire [7:0] t_r38_c32_2;
  wire [7:0] t_r38_c32_3;
  wire [7:0] t_r38_c32_4;
  wire [7:0] t_r38_c32_5;
  wire [7:0] t_r38_c32_6;
  wire [7:0] t_r38_c32_7;
  wire [7:0] t_r38_c32_8;
  wire [7:0] t_r38_c32_9;
  wire [7:0] t_r38_c32_10;
  wire [7:0] t_r38_c32_11;
  wire [7:0] t_r38_c32_12;
  wire [7:0] t_r38_c33_0;
  wire [7:0] t_r38_c33_1;
  wire [7:0] t_r38_c33_2;
  wire [7:0] t_r38_c33_3;
  wire [7:0] t_r38_c33_4;
  wire [7:0] t_r38_c33_5;
  wire [7:0] t_r38_c33_6;
  wire [7:0] t_r38_c33_7;
  wire [7:0] t_r38_c33_8;
  wire [7:0] t_r38_c33_9;
  wire [7:0] t_r38_c33_10;
  wire [7:0] t_r38_c33_11;
  wire [7:0] t_r38_c33_12;
  wire [7:0] t_r38_c34_0;
  wire [7:0] t_r38_c34_1;
  wire [7:0] t_r38_c34_2;
  wire [7:0] t_r38_c34_3;
  wire [7:0] t_r38_c34_4;
  wire [7:0] t_r38_c34_5;
  wire [7:0] t_r38_c34_6;
  wire [7:0] t_r38_c34_7;
  wire [7:0] t_r38_c34_8;
  wire [7:0] t_r38_c34_9;
  wire [7:0] t_r38_c34_10;
  wire [7:0] t_r38_c34_11;
  wire [7:0] t_r38_c34_12;
  wire [7:0] t_r38_c35_0;
  wire [7:0] t_r38_c35_1;
  wire [7:0] t_r38_c35_2;
  wire [7:0] t_r38_c35_3;
  wire [7:0] t_r38_c35_4;
  wire [7:0] t_r38_c35_5;
  wire [7:0] t_r38_c35_6;
  wire [7:0] t_r38_c35_7;
  wire [7:0] t_r38_c35_8;
  wire [7:0] t_r38_c35_9;
  wire [7:0] t_r38_c35_10;
  wire [7:0] t_r38_c35_11;
  wire [7:0] t_r38_c35_12;
  wire [7:0] t_r38_c36_0;
  wire [7:0] t_r38_c36_1;
  wire [7:0] t_r38_c36_2;
  wire [7:0] t_r38_c36_3;
  wire [7:0] t_r38_c36_4;
  wire [7:0] t_r38_c36_5;
  wire [7:0] t_r38_c36_6;
  wire [7:0] t_r38_c36_7;
  wire [7:0] t_r38_c36_8;
  wire [7:0] t_r38_c36_9;
  wire [7:0] t_r38_c36_10;
  wire [7:0] t_r38_c36_11;
  wire [7:0] t_r38_c36_12;
  wire [7:0] t_r38_c37_0;
  wire [7:0] t_r38_c37_1;
  wire [7:0] t_r38_c37_2;
  wire [7:0] t_r38_c37_3;
  wire [7:0] t_r38_c37_4;
  wire [7:0] t_r38_c37_5;
  wire [7:0] t_r38_c37_6;
  wire [7:0] t_r38_c37_7;
  wire [7:0] t_r38_c37_8;
  wire [7:0] t_r38_c37_9;
  wire [7:0] t_r38_c37_10;
  wire [7:0] t_r38_c37_11;
  wire [7:0] t_r38_c37_12;
  wire [7:0] t_r38_c38_0;
  wire [7:0] t_r38_c38_1;
  wire [7:0] t_r38_c38_2;
  wire [7:0] t_r38_c38_3;
  wire [7:0] t_r38_c38_4;
  wire [7:0] t_r38_c38_5;
  wire [7:0] t_r38_c38_6;
  wire [7:0] t_r38_c38_7;
  wire [7:0] t_r38_c38_8;
  wire [7:0] t_r38_c38_9;
  wire [7:0] t_r38_c38_10;
  wire [7:0] t_r38_c38_11;
  wire [7:0] t_r38_c38_12;
  wire [7:0] t_r38_c39_0;
  wire [7:0] t_r38_c39_1;
  wire [7:0] t_r38_c39_2;
  wire [7:0] t_r38_c39_3;
  wire [7:0] t_r38_c39_4;
  wire [7:0] t_r38_c39_5;
  wire [7:0] t_r38_c39_6;
  wire [7:0] t_r38_c39_7;
  wire [7:0] t_r38_c39_8;
  wire [7:0] t_r38_c39_9;
  wire [7:0] t_r38_c39_10;
  wire [7:0] t_r38_c39_11;
  wire [7:0] t_r38_c39_12;
  wire [7:0] t_r38_c40_0;
  wire [7:0] t_r38_c40_1;
  wire [7:0] t_r38_c40_2;
  wire [7:0] t_r38_c40_3;
  wire [7:0] t_r38_c40_4;
  wire [7:0] t_r38_c40_5;
  wire [7:0] t_r38_c40_6;
  wire [7:0] t_r38_c40_7;
  wire [7:0] t_r38_c40_8;
  wire [7:0] t_r38_c40_9;
  wire [7:0] t_r38_c40_10;
  wire [7:0] t_r38_c40_11;
  wire [7:0] t_r38_c40_12;
  wire [7:0] t_r38_c41_0;
  wire [7:0] t_r38_c41_1;
  wire [7:0] t_r38_c41_2;
  wire [7:0] t_r38_c41_3;
  wire [7:0] t_r38_c41_4;
  wire [7:0] t_r38_c41_5;
  wire [7:0] t_r38_c41_6;
  wire [7:0] t_r38_c41_7;
  wire [7:0] t_r38_c41_8;
  wire [7:0] t_r38_c41_9;
  wire [7:0] t_r38_c41_10;
  wire [7:0] t_r38_c41_11;
  wire [7:0] t_r38_c41_12;
  wire [7:0] t_r38_c42_0;
  wire [7:0] t_r38_c42_1;
  wire [7:0] t_r38_c42_2;
  wire [7:0] t_r38_c42_3;
  wire [7:0] t_r38_c42_4;
  wire [7:0] t_r38_c42_5;
  wire [7:0] t_r38_c42_6;
  wire [7:0] t_r38_c42_7;
  wire [7:0] t_r38_c42_8;
  wire [7:0] t_r38_c42_9;
  wire [7:0] t_r38_c42_10;
  wire [7:0] t_r38_c42_11;
  wire [7:0] t_r38_c42_12;
  wire [7:0] t_r38_c43_0;
  wire [7:0] t_r38_c43_1;
  wire [7:0] t_r38_c43_2;
  wire [7:0] t_r38_c43_3;
  wire [7:0] t_r38_c43_4;
  wire [7:0] t_r38_c43_5;
  wire [7:0] t_r38_c43_6;
  wire [7:0] t_r38_c43_7;
  wire [7:0] t_r38_c43_8;
  wire [7:0] t_r38_c43_9;
  wire [7:0] t_r38_c43_10;
  wire [7:0] t_r38_c43_11;
  wire [7:0] t_r38_c43_12;
  wire [7:0] t_r38_c44_0;
  wire [7:0] t_r38_c44_1;
  wire [7:0] t_r38_c44_2;
  wire [7:0] t_r38_c44_3;
  wire [7:0] t_r38_c44_4;
  wire [7:0] t_r38_c44_5;
  wire [7:0] t_r38_c44_6;
  wire [7:0] t_r38_c44_7;
  wire [7:0] t_r38_c44_8;
  wire [7:0] t_r38_c44_9;
  wire [7:0] t_r38_c44_10;
  wire [7:0] t_r38_c44_11;
  wire [7:0] t_r38_c44_12;
  wire [7:0] t_r38_c45_0;
  wire [7:0] t_r38_c45_1;
  wire [7:0] t_r38_c45_2;
  wire [7:0] t_r38_c45_3;
  wire [7:0] t_r38_c45_4;
  wire [7:0] t_r38_c45_5;
  wire [7:0] t_r38_c45_6;
  wire [7:0] t_r38_c45_7;
  wire [7:0] t_r38_c45_8;
  wire [7:0] t_r38_c45_9;
  wire [7:0] t_r38_c45_10;
  wire [7:0] t_r38_c45_11;
  wire [7:0] t_r38_c45_12;
  wire [7:0] t_r38_c46_0;
  wire [7:0] t_r38_c46_1;
  wire [7:0] t_r38_c46_2;
  wire [7:0] t_r38_c46_3;
  wire [7:0] t_r38_c46_4;
  wire [7:0] t_r38_c46_5;
  wire [7:0] t_r38_c46_6;
  wire [7:0] t_r38_c46_7;
  wire [7:0] t_r38_c46_8;
  wire [7:0] t_r38_c46_9;
  wire [7:0] t_r38_c46_10;
  wire [7:0] t_r38_c46_11;
  wire [7:0] t_r38_c46_12;
  wire [7:0] t_r38_c47_0;
  wire [7:0] t_r38_c47_1;
  wire [7:0] t_r38_c47_2;
  wire [7:0] t_r38_c47_3;
  wire [7:0] t_r38_c47_4;
  wire [7:0] t_r38_c47_5;
  wire [7:0] t_r38_c47_6;
  wire [7:0] t_r38_c47_7;
  wire [7:0] t_r38_c47_8;
  wire [7:0] t_r38_c47_9;
  wire [7:0] t_r38_c47_10;
  wire [7:0] t_r38_c47_11;
  wire [7:0] t_r38_c47_12;
  wire [7:0] t_r38_c48_0;
  wire [7:0] t_r38_c48_1;
  wire [7:0] t_r38_c48_2;
  wire [7:0] t_r38_c48_3;
  wire [7:0] t_r38_c48_4;
  wire [7:0] t_r38_c48_5;
  wire [7:0] t_r38_c48_6;
  wire [7:0] t_r38_c48_7;
  wire [7:0] t_r38_c48_8;
  wire [7:0] t_r38_c48_9;
  wire [7:0] t_r38_c48_10;
  wire [7:0] t_r38_c48_11;
  wire [7:0] t_r38_c48_12;
  wire [7:0] t_r38_c49_0;
  wire [7:0] t_r38_c49_1;
  wire [7:0] t_r38_c49_2;
  wire [7:0] t_r38_c49_3;
  wire [7:0] t_r38_c49_4;
  wire [7:0] t_r38_c49_5;
  wire [7:0] t_r38_c49_6;
  wire [7:0] t_r38_c49_7;
  wire [7:0] t_r38_c49_8;
  wire [7:0] t_r38_c49_9;
  wire [7:0] t_r38_c49_10;
  wire [7:0] t_r38_c49_11;
  wire [7:0] t_r38_c49_12;
  wire [7:0] t_r38_c50_0;
  wire [7:0] t_r38_c50_1;
  wire [7:0] t_r38_c50_2;
  wire [7:0] t_r38_c50_3;
  wire [7:0] t_r38_c50_4;
  wire [7:0] t_r38_c50_5;
  wire [7:0] t_r38_c50_6;
  wire [7:0] t_r38_c50_7;
  wire [7:0] t_r38_c50_8;
  wire [7:0] t_r38_c50_9;
  wire [7:0] t_r38_c50_10;
  wire [7:0] t_r38_c50_11;
  wire [7:0] t_r38_c50_12;
  wire [7:0] t_r38_c51_0;
  wire [7:0] t_r38_c51_1;
  wire [7:0] t_r38_c51_2;
  wire [7:0] t_r38_c51_3;
  wire [7:0] t_r38_c51_4;
  wire [7:0] t_r38_c51_5;
  wire [7:0] t_r38_c51_6;
  wire [7:0] t_r38_c51_7;
  wire [7:0] t_r38_c51_8;
  wire [7:0] t_r38_c51_9;
  wire [7:0] t_r38_c51_10;
  wire [7:0] t_r38_c51_11;
  wire [7:0] t_r38_c51_12;
  wire [7:0] t_r38_c52_0;
  wire [7:0] t_r38_c52_1;
  wire [7:0] t_r38_c52_2;
  wire [7:0] t_r38_c52_3;
  wire [7:0] t_r38_c52_4;
  wire [7:0] t_r38_c52_5;
  wire [7:0] t_r38_c52_6;
  wire [7:0] t_r38_c52_7;
  wire [7:0] t_r38_c52_8;
  wire [7:0] t_r38_c52_9;
  wire [7:0] t_r38_c52_10;
  wire [7:0] t_r38_c52_11;
  wire [7:0] t_r38_c52_12;
  wire [7:0] t_r38_c53_0;
  wire [7:0] t_r38_c53_1;
  wire [7:0] t_r38_c53_2;
  wire [7:0] t_r38_c53_3;
  wire [7:0] t_r38_c53_4;
  wire [7:0] t_r38_c53_5;
  wire [7:0] t_r38_c53_6;
  wire [7:0] t_r38_c53_7;
  wire [7:0] t_r38_c53_8;
  wire [7:0] t_r38_c53_9;
  wire [7:0] t_r38_c53_10;
  wire [7:0] t_r38_c53_11;
  wire [7:0] t_r38_c53_12;
  wire [7:0] t_r38_c54_0;
  wire [7:0] t_r38_c54_1;
  wire [7:0] t_r38_c54_2;
  wire [7:0] t_r38_c54_3;
  wire [7:0] t_r38_c54_4;
  wire [7:0] t_r38_c54_5;
  wire [7:0] t_r38_c54_6;
  wire [7:0] t_r38_c54_7;
  wire [7:0] t_r38_c54_8;
  wire [7:0] t_r38_c54_9;
  wire [7:0] t_r38_c54_10;
  wire [7:0] t_r38_c54_11;
  wire [7:0] t_r38_c54_12;
  wire [7:0] t_r38_c55_0;
  wire [7:0] t_r38_c55_1;
  wire [7:0] t_r38_c55_2;
  wire [7:0] t_r38_c55_3;
  wire [7:0] t_r38_c55_4;
  wire [7:0] t_r38_c55_5;
  wire [7:0] t_r38_c55_6;
  wire [7:0] t_r38_c55_7;
  wire [7:0] t_r38_c55_8;
  wire [7:0] t_r38_c55_9;
  wire [7:0] t_r38_c55_10;
  wire [7:0] t_r38_c55_11;
  wire [7:0] t_r38_c55_12;
  wire [7:0] t_r38_c56_0;
  wire [7:0] t_r38_c56_1;
  wire [7:0] t_r38_c56_2;
  wire [7:0] t_r38_c56_3;
  wire [7:0] t_r38_c56_4;
  wire [7:0] t_r38_c56_5;
  wire [7:0] t_r38_c56_6;
  wire [7:0] t_r38_c56_7;
  wire [7:0] t_r38_c56_8;
  wire [7:0] t_r38_c56_9;
  wire [7:0] t_r38_c56_10;
  wire [7:0] t_r38_c56_11;
  wire [7:0] t_r38_c56_12;
  wire [7:0] t_r38_c57_0;
  wire [7:0] t_r38_c57_1;
  wire [7:0] t_r38_c57_2;
  wire [7:0] t_r38_c57_3;
  wire [7:0] t_r38_c57_4;
  wire [7:0] t_r38_c57_5;
  wire [7:0] t_r38_c57_6;
  wire [7:0] t_r38_c57_7;
  wire [7:0] t_r38_c57_8;
  wire [7:0] t_r38_c57_9;
  wire [7:0] t_r38_c57_10;
  wire [7:0] t_r38_c57_11;
  wire [7:0] t_r38_c57_12;
  wire [7:0] t_r38_c58_0;
  wire [7:0] t_r38_c58_1;
  wire [7:0] t_r38_c58_2;
  wire [7:0] t_r38_c58_3;
  wire [7:0] t_r38_c58_4;
  wire [7:0] t_r38_c58_5;
  wire [7:0] t_r38_c58_6;
  wire [7:0] t_r38_c58_7;
  wire [7:0] t_r38_c58_8;
  wire [7:0] t_r38_c58_9;
  wire [7:0] t_r38_c58_10;
  wire [7:0] t_r38_c58_11;
  wire [7:0] t_r38_c58_12;
  wire [7:0] t_r38_c59_0;
  wire [7:0] t_r38_c59_1;
  wire [7:0] t_r38_c59_2;
  wire [7:0] t_r38_c59_3;
  wire [7:0] t_r38_c59_4;
  wire [7:0] t_r38_c59_5;
  wire [7:0] t_r38_c59_6;
  wire [7:0] t_r38_c59_7;
  wire [7:0] t_r38_c59_8;
  wire [7:0] t_r38_c59_9;
  wire [7:0] t_r38_c59_10;
  wire [7:0] t_r38_c59_11;
  wire [7:0] t_r38_c59_12;
  wire [7:0] t_r38_c60_0;
  wire [7:0] t_r38_c60_1;
  wire [7:0] t_r38_c60_2;
  wire [7:0] t_r38_c60_3;
  wire [7:0] t_r38_c60_4;
  wire [7:0] t_r38_c60_5;
  wire [7:0] t_r38_c60_6;
  wire [7:0] t_r38_c60_7;
  wire [7:0] t_r38_c60_8;
  wire [7:0] t_r38_c60_9;
  wire [7:0] t_r38_c60_10;
  wire [7:0] t_r38_c60_11;
  wire [7:0] t_r38_c60_12;
  wire [7:0] t_r38_c61_0;
  wire [7:0] t_r38_c61_1;
  wire [7:0] t_r38_c61_2;
  wire [7:0] t_r38_c61_3;
  wire [7:0] t_r38_c61_4;
  wire [7:0] t_r38_c61_5;
  wire [7:0] t_r38_c61_6;
  wire [7:0] t_r38_c61_7;
  wire [7:0] t_r38_c61_8;
  wire [7:0] t_r38_c61_9;
  wire [7:0] t_r38_c61_10;
  wire [7:0] t_r38_c61_11;
  wire [7:0] t_r38_c61_12;
  wire [7:0] t_r38_c62_0;
  wire [7:0] t_r38_c62_1;
  wire [7:0] t_r38_c62_2;
  wire [7:0] t_r38_c62_3;
  wire [7:0] t_r38_c62_4;
  wire [7:0] t_r38_c62_5;
  wire [7:0] t_r38_c62_6;
  wire [7:0] t_r38_c62_7;
  wire [7:0] t_r38_c62_8;
  wire [7:0] t_r38_c62_9;
  wire [7:0] t_r38_c62_10;
  wire [7:0] t_r38_c62_11;
  wire [7:0] t_r38_c62_12;
  wire [7:0] t_r38_c63_0;
  wire [7:0] t_r38_c63_1;
  wire [7:0] t_r38_c63_2;
  wire [7:0] t_r38_c63_3;
  wire [7:0] t_r38_c63_4;
  wire [7:0] t_r38_c63_5;
  wire [7:0] t_r38_c63_6;
  wire [7:0] t_r38_c63_7;
  wire [7:0] t_r38_c63_8;
  wire [7:0] t_r38_c63_9;
  wire [7:0] t_r38_c63_10;
  wire [7:0] t_r38_c63_11;
  wire [7:0] t_r38_c63_12;
  wire [7:0] t_r38_c64_0;
  wire [7:0] t_r38_c64_1;
  wire [7:0] t_r38_c64_2;
  wire [7:0] t_r38_c64_3;
  wire [7:0] t_r38_c64_4;
  wire [7:0] t_r38_c64_5;
  wire [7:0] t_r38_c64_6;
  wire [7:0] t_r38_c64_7;
  wire [7:0] t_r38_c64_8;
  wire [7:0] t_r38_c64_9;
  wire [7:0] t_r38_c64_10;
  wire [7:0] t_r38_c64_11;
  wire [7:0] t_r38_c64_12;
  wire [7:0] t_r38_c65_0;
  wire [7:0] t_r38_c65_1;
  wire [7:0] t_r38_c65_2;
  wire [7:0] t_r38_c65_3;
  wire [7:0] t_r38_c65_4;
  wire [7:0] t_r38_c65_5;
  wire [7:0] t_r38_c65_6;
  wire [7:0] t_r38_c65_7;
  wire [7:0] t_r38_c65_8;
  wire [7:0] t_r38_c65_9;
  wire [7:0] t_r38_c65_10;
  wire [7:0] t_r38_c65_11;
  wire [7:0] t_r38_c65_12;
  wire [7:0] t_r39_c0_0;
  wire [7:0] t_r39_c0_1;
  wire [7:0] t_r39_c0_2;
  wire [7:0] t_r39_c0_3;
  wire [7:0] t_r39_c0_4;
  wire [7:0] t_r39_c0_5;
  wire [7:0] t_r39_c0_6;
  wire [7:0] t_r39_c0_7;
  wire [7:0] t_r39_c0_8;
  wire [7:0] t_r39_c0_9;
  wire [7:0] t_r39_c0_10;
  wire [7:0] t_r39_c0_11;
  wire [7:0] t_r39_c0_12;
  wire [7:0] t_r39_c1_0;
  wire [7:0] t_r39_c1_1;
  wire [7:0] t_r39_c1_2;
  wire [7:0] t_r39_c1_3;
  wire [7:0] t_r39_c1_4;
  wire [7:0] t_r39_c1_5;
  wire [7:0] t_r39_c1_6;
  wire [7:0] t_r39_c1_7;
  wire [7:0] t_r39_c1_8;
  wire [7:0] t_r39_c1_9;
  wire [7:0] t_r39_c1_10;
  wire [7:0] t_r39_c1_11;
  wire [7:0] t_r39_c1_12;
  wire [7:0] t_r39_c2_0;
  wire [7:0] t_r39_c2_1;
  wire [7:0] t_r39_c2_2;
  wire [7:0] t_r39_c2_3;
  wire [7:0] t_r39_c2_4;
  wire [7:0] t_r39_c2_5;
  wire [7:0] t_r39_c2_6;
  wire [7:0] t_r39_c2_7;
  wire [7:0] t_r39_c2_8;
  wire [7:0] t_r39_c2_9;
  wire [7:0] t_r39_c2_10;
  wire [7:0] t_r39_c2_11;
  wire [7:0] t_r39_c2_12;
  wire [7:0] t_r39_c3_0;
  wire [7:0] t_r39_c3_1;
  wire [7:0] t_r39_c3_2;
  wire [7:0] t_r39_c3_3;
  wire [7:0] t_r39_c3_4;
  wire [7:0] t_r39_c3_5;
  wire [7:0] t_r39_c3_6;
  wire [7:0] t_r39_c3_7;
  wire [7:0] t_r39_c3_8;
  wire [7:0] t_r39_c3_9;
  wire [7:0] t_r39_c3_10;
  wire [7:0] t_r39_c3_11;
  wire [7:0] t_r39_c3_12;
  wire [7:0] t_r39_c4_0;
  wire [7:0] t_r39_c4_1;
  wire [7:0] t_r39_c4_2;
  wire [7:0] t_r39_c4_3;
  wire [7:0] t_r39_c4_4;
  wire [7:0] t_r39_c4_5;
  wire [7:0] t_r39_c4_6;
  wire [7:0] t_r39_c4_7;
  wire [7:0] t_r39_c4_8;
  wire [7:0] t_r39_c4_9;
  wire [7:0] t_r39_c4_10;
  wire [7:0] t_r39_c4_11;
  wire [7:0] t_r39_c4_12;
  wire [7:0] t_r39_c5_0;
  wire [7:0] t_r39_c5_1;
  wire [7:0] t_r39_c5_2;
  wire [7:0] t_r39_c5_3;
  wire [7:0] t_r39_c5_4;
  wire [7:0] t_r39_c5_5;
  wire [7:0] t_r39_c5_6;
  wire [7:0] t_r39_c5_7;
  wire [7:0] t_r39_c5_8;
  wire [7:0] t_r39_c5_9;
  wire [7:0] t_r39_c5_10;
  wire [7:0] t_r39_c5_11;
  wire [7:0] t_r39_c5_12;
  wire [7:0] t_r39_c6_0;
  wire [7:0] t_r39_c6_1;
  wire [7:0] t_r39_c6_2;
  wire [7:0] t_r39_c6_3;
  wire [7:0] t_r39_c6_4;
  wire [7:0] t_r39_c6_5;
  wire [7:0] t_r39_c6_6;
  wire [7:0] t_r39_c6_7;
  wire [7:0] t_r39_c6_8;
  wire [7:0] t_r39_c6_9;
  wire [7:0] t_r39_c6_10;
  wire [7:0] t_r39_c6_11;
  wire [7:0] t_r39_c6_12;
  wire [7:0] t_r39_c7_0;
  wire [7:0] t_r39_c7_1;
  wire [7:0] t_r39_c7_2;
  wire [7:0] t_r39_c7_3;
  wire [7:0] t_r39_c7_4;
  wire [7:0] t_r39_c7_5;
  wire [7:0] t_r39_c7_6;
  wire [7:0] t_r39_c7_7;
  wire [7:0] t_r39_c7_8;
  wire [7:0] t_r39_c7_9;
  wire [7:0] t_r39_c7_10;
  wire [7:0] t_r39_c7_11;
  wire [7:0] t_r39_c7_12;
  wire [7:0] t_r39_c8_0;
  wire [7:0] t_r39_c8_1;
  wire [7:0] t_r39_c8_2;
  wire [7:0] t_r39_c8_3;
  wire [7:0] t_r39_c8_4;
  wire [7:0] t_r39_c8_5;
  wire [7:0] t_r39_c8_6;
  wire [7:0] t_r39_c8_7;
  wire [7:0] t_r39_c8_8;
  wire [7:0] t_r39_c8_9;
  wire [7:0] t_r39_c8_10;
  wire [7:0] t_r39_c8_11;
  wire [7:0] t_r39_c8_12;
  wire [7:0] t_r39_c9_0;
  wire [7:0] t_r39_c9_1;
  wire [7:0] t_r39_c9_2;
  wire [7:0] t_r39_c9_3;
  wire [7:0] t_r39_c9_4;
  wire [7:0] t_r39_c9_5;
  wire [7:0] t_r39_c9_6;
  wire [7:0] t_r39_c9_7;
  wire [7:0] t_r39_c9_8;
  wire [7:0] t_r39_c9_9;
  wire [7:0] t_r39_c9_10;
  wire [7:0] t_r39_c9_11;
  wire [7:0] t_r39_c9_12;
  wire [7:0] t_r39_c10_0;
  wire [7:0] t_r39_c10_1;
  wire [7:0] t_r39_c10_2;
  wire [7:0] t_r39_c10_3;
  wire [7:0] t_r39_c10_4;
  wire [7:0] t_r39_c10_5;
  wire [7:0] t_r39_c10_6;
  wire [7:0] t_r39_c10_7;
  wire [7:0] t_r39_c10_8;
  wire [7:0] t_r39_c10_9;
  wire [7:0] t_r39_c10_10;
  wire [7:0] t_r39_c10_11;
  wire [7:0] t_r39_c10_12;
  wire [7:0] t_r39_c11_0;
  wire [7:0] t_r39_c11_1;
  wire [7:0] t_r39_c11_2;
  wire [7:0] t_r39_c11_3;
  wire [7:0] t_r39_c11_4;
  wire [7:0] t_r39_c11_5;
  wire [7:0] t_r39_c11_6;
  wire [7:0] t_r39_c11_7;
  wire [7:0] t_r39_c11_8;
  wire [7:0] t_r39_c11_9;
  wire [7:0] t_r39_c11_10;
  wire [7:0] t_r39_c11_11;
  wire [7:0] t_r39_c11_12;
  wire [7:0] t_r39_c12_0;
  wire [7:0] t_r39_c12_1;
  wire [7:0] t_r39_c12_2;
  wire [7:0] t_r39_c12_3;
  wire [7:0] t_r39_c12_4;
  wire [7:0] t_r39_c12_5;
  wire [7:0] t_r39_c12_6;
  wire [7:0] t_r39_c12_7;
  wire [7:0] t_r39_c12_8;
  wire [7:0] t_r39_c12_9;
  wire [7:0] t_r39_c12_10;
  wire [7:0] t_r39_c12_11;
  wire [7:0] t_r39_c12_12;
  wire [7:0] t_r39_c13_0;
  wire [7:0] t_r39_c13_1;
  wire [7:0] t_r39_c13_2;
  wire [7:0] t_r39_c13_3;
  wire [7:0] t_r39_c13_4;
  wire [7:0] t_r39_c13_5;
  wire [7:0] t_r39_c13_6;
  wire [7:0] t_r39_c13_7;
  wire [7:0] t_r39_c13_8;
  wire [7:0] t_r39_c13_9;
  wire [7:0] t_r39_c13_10;
  wire [7:0] t_r39_c13_11;
  wire [7:0] t_r39_c13_12;
  wire [7:0] t_r39_c14_0;
  wire [7:0] t_r39_c14_1;
  wire [7:0] t_r39_c14_2;
  wire [7:0] t_r39_c14_3;
  wire [7:0] t_r39_c14_4;
  wire [7:0] t_r39_c14_5;
  wire [7:0] t_r39_c14_6;
  wire [7:0] t_r39_c14_7;
  wire [7:0] t_r39_c14_8;
  wire [7:0] t_r39_c14_9;
  wire [7:0] t_r39_c14_10;
  wire [7:0] t_r39_c14_11;
  wire [7:0] t_r39_c14_12;
  wire [7:0] t_r39_c15_0;
  wire [7:0] t_r39_c15_1;
  wire [7:0] t_r39_c15_2;
  wire [7:0] t_r39_c15_3;
  wire [7:0] t_r39_c15_4;
  wire [7:0] t_r39_c15_5;
  wire [7:0] t_r39_c15_6;
  wire [7:0] t_r39_c15_7;
  wire [7:0] t_r39_c15_8;
  wire [7:0] t_r39_c15_9;
  wire [7:0] t_r39_c15_10;
  wire [7:0] t_r39_c15_11;
  wire [7:0] t_r39_c15_12;
  wire [7:0] t_r39_c16_0;
  wire [7:0] t_r39_c16_1;
  wire [7:0] t_r39_c16_2;
  wire [7:0] t_r39_c16_3;
  wire [7:0] t_r39_c16_4;
  wire [7:0] t_r39_c16_5;
  wire [7:0] t_r39_c16_6;
  wire [7:0] t_r39_c16_7;
  wire [7:0] t_r39_c16_8;
  wire [7:0] t_r39_c16_9;
  wire [7:0] t_r39_c16_10;
  wire [7:0] t_r39_c16_11;
  wire [7:0] t_r39_c16_12;
  wire [7:0] t_r39_c17_0;
  wire [7:0] t_r39_c17_1;
  wire [7:0] t_r39_c17_2;
  wire [7:0] t_r39_c17_3;
  wire [7:0] t_r39_c17_4;
  wire [7:0] t_r39_c17_5;
  wire [7:0] t_r39_c17_6;
  wire [7:0] t_r39_c17_7;
  wire [7:0] t_r39_c17_8;
  wire [7:0] t_r39_c17_9;
  wire [7:0] t_r39_c17_10;
  wire [7:0] t_r39_c17_11;
  wire [7:0] t_r39_c17_12;
  wire [7:0] t_r39_c18_0;
  wire [7:0] t_r39_c18_1;
  wire [7:0] t_r39_c18_2;
  wire [7:0] t_r39_c18_3;
  wire [7:0] t_r39_c18_4;
  wire [7:0] t_r39_c18_5;
  wire [7:0] t_r39_c18_6;
  wire [7:0] t_r39_c18_7;
  wire [7:0] t_r39_c18_8;
  wire [7:0] t_r39_c18_9;
  wire [7:0] t_r39_c18_10;
  wire [7:0] t_r39_c18_11;
  wire [7:0] t_r39_c18_12;
  wire [7:0] t_r39_c19_0;
  wire [7:0] t_r39_c19_1;
  wire [7:0] t_r39_c19_2;
  wire [7:0] t_r39_c19_3;
  wire [7:0] t_r39_c19_4;
  wire [7:0] t_r39_c19_5;
  wire [7:0] t_r39_c19_6;
  wire [7:0] t_r39_c19_7;
  wire [7:0] t_r39_c19_8;
  wire [7:0] t_r39_c19_9;
  wire [7:0] t_r39_c19_10;
  wire [7:0] t_r39_c19_11;
  wire [7:0] t_r39_c19_12;
  wire [7:0] t_r39_c20_0;
  wire [7:0] t_r39_c20_1;
  wire [7:0] t_r39_c20_2;
  wire [7:0] t_r39_c20_3;
  wire [7:0] t_r39_c20_4;
  wire [7:0] t_r39_c20_5;
  wire [7:0] t_r39_c20_6;
  wire [7:0] t_r39_c20_7;
  wire [7:0] t_r39_c20_8;
  wire [7:0] t_r39_c20_9;
  wire [7:0] t_r39_c20_10;
  wire [7:0] t_r39_c20_11;
  wire [7:0] t_r39_c20_12;
  wire [7:0] t_r39_c21_0;
  wire [7:0] t_r39_c21_1;
  wire [7:0] t_r39_c21_2;
  wire [7:0] t_r39_c21_3;
  wire [7:0] t_r39_c21_4;
  wire [7:0] t_r39_c21_5;
  wire [7:0] t_r39_c21_6;
  wire [7:0] t_r39_c21_7;
  wire [7:0] t_r39_c21_8;
  wire [7:0] t_r39_c21_9;
  wire [7:0] t_r39_c21_10;
  wire [7:0] t_r39_c21_11;
  wire [7:0] t_r39_c21_12;
  wire [7:0] t_r39_c22_0;
  wire [7:0] t_r39_c22_1;
  wire [7:0] t_r39_c22_2;
  wire [7:0] t_r39_c22_3;
  wire [7:0] t_r39_c22_4;
  wire [7:0] t_r39_c22_5;
  wire [7:0] t_r39_c22_6;
  wire [7:0] t_r39_c22_7;
  wire [7:0] t_r39_c22_8;
  wire [7:0] t_r39_c22_9;
  wire [7:0] t_r39_c22_10;
  wire [7:0] t_r39_c22_11;
  wire [7:0] t_r39_c22_12;
  wire [7:0] t_r39_c23_0;
  wire [7:0] t_r39_c23_1;
  wire [7:0] t_r39_c23_2;
  wire [7:0] t_r39_c23_3;
  wire [7:0] t_r39_c23_4;
  wire [7:0] t_r39_c23_5;
  wire [7:0] t_r39_c23_6;
  wire [7:0] t_r39_c23_7;
  wire [7:0] t_r39_c23_8;
  wire [7:0] t_r39_c23_9;
  wire [7:0] t_r39_c23_10;
  wire [7:0] t_r39_c23_11;
  wire [7:0] t_r39_c23_12;
  wire [7:0] t_r39_c24_0;
  wire [7:0] t_r39_c24_1;
  wire [7:0] t_r39_c24_2;
  wire [7:0] t_r39_c24_3;
  wire [7:0] t_r39_c24_4;
  wire [7:0] t_r39_c24_5;
  wire [7:0] t_r39_c24_6;
  wire [7:0] t_r39_c24_7;
  wire [7:0] t_r39_c24_8;
  wire [7:0] t_r39_c24_9;
  wire [7:0] t_r39_c24_10;
  wire [7:0] t_r39_c24_11;
  wire [7:0] t_r39_c24_12;
  wire [7:0] t_r39_c25_0;
  wire [7:0] t_r39_c25_1;
  wire [7:0] t_r39_c25_2;
  wire [7:0] t_r39_c25_3;
  wire [7:0] t_r39_c25_4;
  wire [7:0] t_r39_c25_5;
  wire [7:0] t_r39_c25_6;
  wire [7:0] t_r39_c25_7;
  wire [7:0] t_r39_c25_8;
  wire [7:0] t_r39_c25_9;
  wire [7:0] t_r39_c25_10;
  wire [7:0] t_r39_c25_11;
  wire [7:0] t_r39_c25_12;
  wire [7:0] t_r39_c26_0;
  wire [7:0] t_r39_c26_1;
  wire [7:0] t_r39_c26_2;
  wire [7:0] t_r39_c26_3;
  wire [7:0] t_r39_c26_4;
  wire [7:0] t_r39_c26_5;
  wire [7:0] t_r39_c26_6;
  wire [7:0] t_r39_c26_7;
  wire [7:0] t_r39_c26_8;
  wire [7:0] t_r39_c26_9;
  wire [7:0] t_r39_c26_10;
  wire [7:0] t_r39_c26_11;
  wire [7:0] t_r39_c26_12;
  wire [7:0] t_r39_c27_0;
  wire [7:0] t_r39_c27_1;
  wire [7:0] t_r39_c27_2;
  wire [7:0] t_r39_c27_3;
  wire [7:0] t_r39_c27_4;
  wire [7:0] t_r39_c27_5;
  wire [7:0] t_r39_c27_6;
  wire [7:0] t_r39_c27_7;
  wire [7:0] t_r39_c27_8;
  wire [7:0] t_r39_c27_9;
  wire [7:0] t_r39_c27_10;
  wire [7:0] t_r39_c27_11;
  wire [7:0] t_r39_c27_12;
  wire [7:0] t_r39_c28_0;
  wire [7:0] t_r39_c28_1;
  wire [7:0] t_r39_c28_2;
  wire [7:0] t_r39_c28_3;
  wire [7:0] t_r39_c28_4;
  wire [7:0] t_r39_c28_5;
  wire [7:0] t_r39_c28_6;
  wire [7:0] t_r39_c28_7;
  wire [7:0] t_r39_c28_8;
  wire [7:0] t_r39_c28_9;
  wire [7:0] t_r39_c28_10;
  wire [7:0] t_r39_c28_11;
  wire [7:0] t_r39_c28_12;
  wire [7:0] t_r39_c29_0;
  wire [7:0] t_r39_c29_1;
  wire [7:0] t_r39_c29_2;
  wire [7:0] t_r39_c29_3;
  wire [7:0] t_r39_c29_4;
  wire [7:0] t_r39_c29_5;
  wire [7:0] t_r39_c29_6;
  wire [7:0] t_r39_c29_7;
  wire [7:0] t_r39_c29_8;
  wire [7:0] t_r39_c29_9;
  wire [7:0] t_r39_c29_10;
  wire [7:0] t_r39_c29_11;
  wire [7:0] t_r39_c29_12;
  wire [7:0] t_r39_c30_0;
  wire [7:0] t_r39_c30_1;
  wire [7:0] t_r39_c30_2;
  wire [7:0] t_r39_c30_3;
  wire [7:0] t_r39_c30_4;
  wire [7:0] t_r39_c30_5;
  wire [7:0] t_r39_c30_6;
  wire [7:0] t_r39_c30_7;
  wire [7:0] t_r39_c30_8;
  wire [7:0] t_r39_c30_9;
  wire [7:0] t_r39_c30_10;
  wire [7:0] t_r39_c30_11;
  wire [7:0] t_r39_c30_12;
  wire [7:0] t_r39_c31_0;
  wire [7:0] t_r39_c31_1;
  wire [7:0] t_r39_c31_2;
  wire [7:0] t_r39_c31_3;
  wire [7:0] t_r39_c31_4;
  wire [7:0] t_r39_c31_5;
  wire [7:0] t_r39_c31_6;
  wire [7:0] t_r39_c31_7;
  wire [7:0] t_r39_c31_8;
  wire [7:0] t_r39_c31_9;
  wire [7:0] t_r39_c31_10;
  wire [7:0] t_r39_c31_11;
  wire [7:0] t_r39_c31_12;
  wire [7:0] t_r39_c32_0;
  wire [7:0] t_r39_c32_1;
  wire [7:0] t_r39_c32_2;
  wire [7:0] t_r39_c32_3;
  wire [7:0] t_r39_c32_4;
  wire [7:0] t_r39_c32_5;
  wire [7:0] t_r39_c32_6;
  wire [7:0] t_r39_c32_7;
  wire [7:0] t_r39_c32_8;
  wire [7:0] t_r39_c32_9;
  wire [7:0] t_r39_c32_10;
  wire [7:0] t_r39_c32_11;
  wire [7:0] t_r39_c32_12;
  wire [7:0] t_r39_c33_0;
  wire [7:0] t_r39_c33_1;
  wire [7:0] t_r39_c33_2;
  wire [7:0] t_r39_c33_3;
  wire [7:0] t_r39_c33_4;
  wire [7:0] t_r39_c33_5;
  wire [7:0] t_r39_c33_6;
  wire [7:0] t_r39_c33_7;
  wire [7:0] t_r39_c33_8;
  wire [7:0] t_r39_c33_9;
  wire [7:0] t_r39_c33_10;
  wire [7:0] t_r39_c33_11;
  wire [7:0] t_r39_c33_12;
  wire [7:0] t_r39_c34_0;
  wire [7:0] t_r39_c34_1;
  wire [7:0] t_r39_c34_2;
  wire [7:0] t_r39_c34_3;
  wire [7:0] t_r39_c34_4;
  wire [7:0] t_r39_c34_5;
  wire [7:0] t_r39_c34_6;
  wire [7:0] t_r39_c34_7;
  wire [7:0] t_r39_c34_8;
  wire [7:0] t_r39_c34_9;
  wire [7:0] t_r39_c34_10;
  wire [7:0] t_r39_c34_11;
  wire [7:0] t_r39_c34_12;
  wire [7:0] t_r39_c35_0;
  wire [7:0] t_r39_c35_1;
  wire [7:0] t_r39_c35_2;
  wire [7:0] t_r39_c35_3;
  wire [7:0] t_r39_c35_4;
  wire [7:0] t_r39_c35_5;
  wire [7:0] t_r39_c35_6;
  wire [7:0] t_r39_c35_7;
  wire [7:0] t_r39_c35_8;
  wire [7:0] t_r39_c35_9;
  wire [7:0] t_r39_c35_10;
  wire [7:0] t_r39_c35_11;
  wire [7:0] t_r39_c35_12;
  wire [7:0] t_r39_c36_0;
  wire [7:0] t_r39_c36_1;
  wire [7:0] t_r39_c36_2;
  wire [7:0] t_r39_c36_3;
  wire [7:0] t_r39_c36_4;
  wire [7:0] t_r39_c36_5;
  wire [7:0] t_r39_c36_6;
  wire [7:0] t_r39_c36_7;
  wire [7:0] t_r39_c36_8;
  wire [7:0] t_r39_c36_9;
  wire [7:0] t_r39_c36_10;
  wire [7:0] t_r39_c36_11;
  wire [7:0] t_r39_c36_12;
  wire [7:0] t_r39_c37_0;
  wire [7:0] t_r39_c37_1;
  wire [7:0] t_r39_c37_2;
  wire [7:0] t_r39_c37_3;
  wire [7:0] t_r39_c37_4;
  wire [7:0] t_r39_c37_5;
  wire [7:0] t_r39_c37_6;
  wire [7:0] t_r39_c37_7;
  wire [7:0] t_r39_c37_8;
  wire [7:0] t_r39_c37_9;
  wire [7:0] t_r39_c37_10;
  wire [7:0] t_r39_c37_11;
  wire [7:0] t_r39_c37_12;
  wire [7:0] t_r39_c38_0;
  wire [7:0] t_r39_c38_1;
  wire [7:0] t_r39_c38_2;
  wire [7:0] t_r39_c38_3;
  wire [7:0] t_r39_c38_4;
  wire [7:0] t_r39_c38_5;
  wire [7:0] t_r39_c38_6;
  wire [7:0] t_r39_c38_7;
  wire [7:0] t_r39_c38_8;
  wire [7:0] t_r39_c38_9;
  wire [7:0] t_r39_c38_10;
  wire [7:0] t_r39_c38_11;
  wire [7:0] t_r39_c38_12;
  wire [7:0] t_r39_c39_0;
  wire [7:0] t_r39_c39_1;
  wire [7:0] t_r39_c39_2;
  wire [7:0] t_r39_c39_3;
  wire [7:0] t_r39_c39_4;
  wire [7:0] t_r39_c39_5;
  wire [7:0] t_r39_c39_6;
  wire [7:0] t_r39_c39_7;
  wire [7:0] t_r39_c39_8;
  wire [7:0] t_r39_c39_9;
  wire [7:0] t_r39_c39_10;
  wire [7:0] t_r39_c39_11;
  wire [7:0] t_r39_c39_12;
  wire [7:0] t_r39_c40_0;
  wire [7:0] t_r39_c40_1;
  wire [7:0] t_r39_c40_2;
  wire [7:0] t_r39_c40_3;
  wire [7:0] t_r39_c40_4;
  wire [7:0] t_r39_c40_5;
  wire [7:0] t_r39_c40_6;
  wire [7:0] t_r39_c40_7;
  wire [7:0] t_r39_c40_8;
  wire [7:0] t_r39_c40_9;
  wire [7:0] t_r39_c40_10;
  wire [7:0] t_r39_c40_11;
  wire [7:0] t_r39_c40_12;
  wire [7:0] t_r39_c41_0;
  wire [7:0] t_r39_c41_1;
  wire [7:0] t_r39_c41_2;
  wire [7:0] t_r39_c41_3;
  wire [7:0] t_r39_c41_4;
  wire [7:0] t_r39_c41_5;
  wire [7:0] t_r39_c41_6;
  wire [7:0] t_r39_c41_7;
  wire [7:0] t_r39_c41_8;
  wire [7:0] t_r39_c41_9;
  wire [7:0] t_r39_c41_10;
  wire [7:0] t_r39_c41_11;
  wire [7:0] t_r39_c41_12;
  wire [7:0] t_r39_c42_0;
  wire [7:0] t_r39_c42_1;
  wire [7:0] t_r39_c42_2;
  wire [7:0] t_r39_c42_3;
  wire [7:0] t_r39_c42_4;
  wire [7:0] t_r39_c42_5;
  wire [7:0] t_r39_c42_6;
  wire [7:0] t_r39_c42_7;
  wire [7:0] t_r39_c42_8;
  wire [7:0] t_r39_c42_9;
  wire [7:0] t_r39_c42_10;
  wire [7:0] t_r39_c42_11;
  wire [7:0] t_r39_c42_12;
  wire [7:0] t_r39_c43_0;
  wire [7:0] t_r39_c43_1;
  wire [7:0] t_r39_c43_2;
  wire [7:0] t_r39_c43_3;
  wire [7:0] t_r39_c43_4;
  wire [7:0] t_r39_c43_5;
  wire [7:0] t_r39_c43_6;
  wire [7:0] t_r39_c43_7;
  wire [7:0] t_r39_c43_8;
  wire [7:0] t_r39_c43_9;
  wire [7:0] t_r39_c43_10;
  wire [7:0] t_r39_c43_11;
  wire [7:0] t_r39_c43_12;
  wire [7:0] t_r39_c44_0;
  wire [7:0] t_r39_c44_1;
  wire [7:0] t_r39_c44_2;
  wire [7:0] t_r39_c44_3;
  wire [7:0] t_r39_c44_4;
  wire [7:0] t_r39_c44_5;
  wire [7:0] t_r39_c44_6;
  wire [7:0] t_r39_c44_7;
  wire [7:0] t_r39_c44_8;
  wire [7:0] t_r39_c44_9;
  wire [7:0] t_r39_c44_10;
  wire [7:0] t_r39_c44_11;
  wire [7:0] t_r39_c44_12;
  wire [7:0] t_r39_c45_0;
  wire [7:0] t_r39_c45_1;
  wire [7:0] t_r39_c45_2;
  wire [7:0] t_r39_c45_3;
  wire [7:0] t_r39_c45_4;
  wire [7:0] t_r39_c45_5;
  wire [7:0] t_r39_c45_6;
  wire [7:0] t_r39_c45_7;
  wire [7:0] t_r39_c45_8;
  wire [7:0] t_r39_c45_9;
  wire [7:0] t_r39_c45_10;
  wire [7:0] t_r39_c45_11;
  wire [7:0] t_r39_c45_12;
  wire [7:0] t_r39_c46_0;
  wire [7:0] t_r39_c46_1;
  wire [7:0] t_r39_c46_2;
  wire [7:0] t_r39_c46_3;
  wire [7:0] t_r39_c46_4;
  wire [7:0] t_r39_c46_5;
  wire [7:0] t_r39_c46_6;
  wire [7:0] t_r39_c46_7;
  wire [7:0] t_r39_c46_8;
  wire [7:0] t_r39_c46_9;
  wire [7:0] t_r39_c46_10;
  wire [7:0] t_r39_c46_11;
  wire [7:0] t_r39_c46_12;
  wire [7:0] t_r39_c47_0;
  wire [7:0] t_r39_c47_1;
  wire [7:0] t_r39_c47_2;
  wire [7:0] t_r39_c47_3;
  wire [7:0] t_r39_c47_4;
  wire [7:0] t_r39_c47_5;
  wire [7:0] t_r39_c47_6;
  wire [7:0] t_r39_c47_7;
  wire [7:0] t_r39_c47_8;
  wire [7:0] t_r39_c47_9;
  wire [7:0] t_r39_c47_10;
  wire [7:0] t_r39_c47_11;
  wire [7:0] t_r39_c47_12;
  wire [7:0] t_r39_c48_0;
  wire [7:0] t_r39_c48_1;
  wire [7:0] t_r39_c48_2;
  wire [7:0] t_r39_c48_3;
  wire [7:0] t_r39_c48_4;
  wire [7:0] t_r39_c48_5;
  wire [7:0] t_r39_c48_6;
  wire [7:0] t_r39_c48_7;
  wire [7:0] t_r39_c48_8;
  wire [7:0] t_r39_c48_9;
  wire [7:0] t_r39_c48_10;
  wire [7:0] t_r39_c48_11;
  wire [7:0] t_r39_c48_12;
  wire [7:0] t_r39_c49_0;
  wire [7:0] t_r39_c49_1;
  wire [7:0] t_r39_c49_2;
  wire [7:0] t_r39_c49_3;
  wire [7:0] t_r39_c49_4;
  wire [7:0] t_r39_c49_5;
  wire [7:0] t_r39_c49_6;
  wire [7:0] t_r39_c49_7;
  wire [7:0] t_r39_c49_8;
  wire [7:0] t_r39_c49_9;
  wire [7:0] t_r39_c49_10;
  wire [7:0] t_r39_c49_11;
  wire [7:0] t_r39_c49_12;
  wire [7:0] t_r39_c50_0;
  wire [7:0] t_r39_c50_1;
  wire [7:0] t_r39_c50_2;
  wire [7:0] t_r39_c50_3;
  wire [7:0] t_r39_c50_4;
  wire [7:0] t_r39_c50_5;
  wire [7:0] t_r39_c50_6;
  wire [7:0] t_r39_c50_7;
  wire [7:0] t_r39_c50_8;
  wire [7:0] t_r39_c50_9;
  wire [7:0] t_r39_c50_10;
  wire [7:0] t_r39_c50_11;
  wire [7:0] t_r39_c50_12;
  wire [7:0] t_r39_c51_0;
  wire [7:0] t_r39_c51_1;
  wire [7:0] t_r39_c51_2;
  wire [7:0] t_r39_c51_3;
  wire [7:0] t_r39_c51_4;
  wire [7:0] t_r39_c51_5;
  wire [7:0] t_r39_c51_6;
  wire [7:0] t_r39_c51_7;
  wire [7:0] t_r39_c51_8;
  wire [7:0] t_r39_c51_9;
  wire [7:0] t_r39_c51_10;
  wire [7:0] t_r39_c51_11;
  wire [7:0] t_r39_c51_12;
  wire [7:0] t_r39_c52_0;
  wire [7:0] t_r39_c52_1;
  wire [7:0] t_r39_c52_2;
  wire [7:0] t_r39_c52_3;
  wire [7:0] t_r39_c52_4;
  wire [7:0] t_r39_c52_5;
  wire [7:0] t_r39_c52_6;
  wire [7:0] t_r39_c52_7;
  wire [7:0] t_r39_c52_8;
  wire [7:0] t_r39_c52_9;
  wire [7:0] t_r39_c52_10;
  wire [7:0] t_r39_c52_11;
  wire [7:0] t_r39_c52_12;
  wire [7:0] t_r39_c53_0;
  wire [7:0] t_r39_c53_1;
  wire [7:0] t_r39_c53_2;
  wire [7:0] t_r39_c53_3;
  wire [7:0] t_r39_c53_4;
  wire [7:0] t_r39_c53_5;
  wire [7:0] t_r39_c53_6;
  wire [7:0] t_r39_c53_7;
  wire [7:0] t_r39_c53_8;
  wire [7:0] t_r39_c53_9;
  wire [7:0] t_r39_c53_10;
  wire [7:0] t_r39_c53_11;
  wire [7:0] t_r39_c53_12;
  wire [7:0] t_r39_c54_0;
  wire [7:0] t_r39_c54_1;
  wire [7:0] t_r39_c54_2;
  wire [7:0] t_r39_c54_3;
  wire [7:0] t_r39_c54_4;
  wire [7:0] t_r39_c54_5;
  wire [7:0] t_r39_c54_6;
  wire [7:0] t_r39_c54_7;
  wire [7:0] t_r39_c54_8;
  wire [7:0] t_r39_c54_9;
  wire [7:0] t_r39_c54_10;
  wire [7:0] t_r39_c54_11;
  wire [7:0] t_r39_c54_12;
  wire [7:0] t_r39_c55_0;
  wire [7:0] t_r39_c55_1;
  wire [7:0] t_r39_c55_2;
  wire [7:0] t_r39_c55_3;
  wire [7:0] t_r39_c55_4;
  wire [7:0] t_r39_c55_5;
  wire [7:0] t_r39_c55_6;
  wire [7:0] t_r39_c55_7;
  wire [7:0] t_r39_c55_8;
  wire [7:0] t_r39_c55_9;
  wire [7:0] t_r39_c55_10;
  wire [7:0] t_r39_c55_11;
  wire [7:0] t_r39_c55_12;
  wire [7:0] t_r39_c56_0;
  wire [7:0] t_r39_c56_1;
  wire [7:0] t_r39_c56_2;
  wire [7:0] t_r39_c56_3;
  wire [7:0] t_r39_c56_4;
  wire [7:0] t_r39_c56_5;
  wire [7:0] t_r39_c56_6;
  wire [7:0] t_r39_c56_7;
  wire [7:0] t_r39_c56_8;
  wire [7:0] t_r39_c56_9;
  wire [7:0] t_r39_c56_10;
  wire [7:0] t_r39_c56_11;
  wire [7:0] t_r39_c56_12;
  wire [7:0] t_r39_c57_0;
  wire [7:0] t_r39_c57_1;
  wire [7:0] t_r39_c57_2;
  wire [7:0] t_r39_c57_3;
  wire [7:0] t_r39_c57_4;
  wire [7:0] t_r39_c57_5;
  wire [7:0] t_r39_c57_6;
  wire [7:0] t_r39_c57_7;
  wire [7:0] t_r39_c57_8;
  wire [7:0] t_r39_c57_9;
  wire [7:0] t_r39_c57_10;
  wire [7:0] t_r39_c57_11;
  wire [7:0] t_r39_c57_12;
  wire [7:0] t_r39_c58_0;
  wire [7:0] t_r39_c58_1;
  wire [7:0] t_r39_c58_2;
  wire [7:0] t_r39_c58_3;
  wire [7:0] t_r39_c58_4;
  wire [7:0] t_r39_c58_5;
  wire [7:0] t_r39_c58_6;
  wire [7:0] t_r39_c58_7;
  wire [7:0] t_r39_c58_8;
  wire [7:0] t_r39_c58_9;
  wire [7:0] t_r39_c58_10;
  wire [7:0] t_r39_c58_11;
  wire [7:0] t_r39_c58_12;
  wire [7:0] t_r39_c59_0;
  wire [7:0] t_r39_c59_1;
  wire [7:0] t_r39_c59_2;
  wire [7:0] t_r39_c59_3;
  wire [7:0] t_r39_c59_4;
  wire [7:0] t_r39_c59_5;
  wire [7:0] t_r39_c59_6;
  wire [7:0] t_r39_c59_7;
  wire [7:0] t_r39_c59_8;
  wire [7:0] t_r39_c59_9;
  wire [7:0] t_r39_c59_10;
  wire [7:0] t_r39_c59_11;
  wire [7:0] t_r39_c59_12;
  wire [7:0] t_r39_c60_0;
  wire [7:0] t_r39_c60_1;
  wire [7:0] t_r39_c60_2;
  wire [7:0] t_r39_c60_3;
  wire [7:0] t_r39_c60_4;
  wire [7:0] t_r39_c60_5;
  wire [7:0] t_r39_c60_6;
  wire [7:0] t_r39_c60_7;
  wire [7:0] t_r39_c60_8;
  wire [7:0] t_r39_c60_9;
  wire [7:0] t_r39_c60_10;
  wire [7:0] t_r39_c60_11;
  wire [7:0] t_r39_c60_12;
  wire [7:0] t_r39_c61_0;
  wire [7:0] t_r39_c61_1;
  wire [7:0] t_r39_c61_2;
  wire [7:0] t_r39_c61_3;
  wire [7:0] t_r39_c61_4;
  wire [7:0] t_r39_c61_5;
  wire [7:0] t_r39_c61_6;
  wire [7:0] t_r39_c61_7;
  wire [7:0] t_r39_c61_8;
  wire [7:0] t_r39_c61_9;
  wire [7:0] t_r39_c61_10;
  wire [7:0] t_r39_c61_11;
  wire [7:0] t_r39_c61_12;
  wire [7:0] t_r39_c62_0;
  wire [7:0] t_r39_c62_1;
  wire [7:0] t_r39_c62_2;
  wire [7:0] t_r39_c62_3;
  wire [7:0] t_r39_c62_4;
  wire [7:0] t_r39_c62_5;
  wire [7:0] t_r39_c62_6;
  wire [7:0] t_r39_c62_7;
  wire [7:0] t_r39_c62_8;
  wire [7:0] t_r39_c62_9;
  wire [7:0] t_r39_c62_10;
  wire [7:0] t_r39_c62_11;
  wire [7:0] t_r39_c62_12;
  wire [7:0] t_r39_c63_0;
  wire [7:0] t_r39_c63_1;
  wire [7:0] t_r39_c63_2;
  wire [7:0] t_r39_c63_3;
  wire [7:0] t_r39_c63_4;
  wire [7:0] t_r39_c63_5;
  wire [7:0] t_r39_c63_6;
  wire [7:0] t_r39_c63_7;
  wire [7:0] t_r39_c63_8;
  wire [7:0] t_r39_c63_9;
  wire [7:0] t_r39_c63_10;
  wire [7:0] t_r39_c63_11;
  wire [7:0] t_r39_c63_12;
  wire [7:0] t_r39_c64_0;
  wire [7:0] t_r39_c64_1;
  wire [7:0] t_r39_c64_2;
  wire [7:0] t_r39_c64_3;
  wire [7:0] t_r39_c64_4;
  wire [7:0] t_r39_c64_5;
  wire [7:0] t_r39_c64_6;
  wire [7:0] t_r39_c64_7;
  wire [7:0] t_r39_c64_8;
  wire [7:0] t_r39_c64_9;
  wire [7:0] t_r39_c64_10;
  wire [7:0] t_r39_c64_11;
  wire [7:0] t_r39_c64_12;
  wire [7:0] t_r39_c65_0;
  wire [7:0] t_r39_c65_1;
  wire [7:0] t_r39_c65_2;
  wire [7:0] t_r39_c65_3;
  wire [7:0] t_r39_c65_4;
  wire [7:0] t_r39_c65_5;
  wire [7:0] t_r39_c65_6;
  wire [7:0] t_r39_c65_7;
  wire [7:0] t_r39_c65_8;
  wire [7:0] t_r39_c65_9;
  wire [7:0] t_r39_c65_10;
  wire [7:0] t_r39_c65_11;
  wire [7:0] t_r39_c65_12;
  wire [7:0] t_r40_c0_0;
  wire [7:0] t_r40_c0_1;
  wire [7:0] t_r40_c0_2;
  wire [7:0] t_r40_c0_3;
  wire [7:0] t_r40_c0_4;
  wire [7:0] t_r40_c0_5;
  wire [7:0] t_r40_c0_6;
  wire [7:0] t_r40_c0_7;
  wire [7:0] t_r40_c0_8;
  wire [7:0] t_r40_c0_9;
  wire [7:0] t_r40_c0_10;
  wire [7:0] t_r40_c0_11;
  wire [7:0] t_r40_c0_12;
  wire [7:0] t_r40_c1_0;
  wire [7:0] t_r40_c1_1;
  wire [7:0] t_r40_c1_2;
  wire [7:0] t_r40_c1_3;
  wire [7:0] t_r40_c1_4;
  wire [7:0] t_r40_c1_5;
  wire [7:0] t_r40_c1_6;
  wire [7:0] t_r40_c1_7;
  wire [7:0] t_r40_c1_8;
  wire [7:0] t_r40_c1_9;
  wire [7:0] t_r40_c1_10;
  wire [7:0] t_r40_c1_11;
  wire [7:0] t_r40_c1_12;
  wire [7:0] t_r40_c2_0;
  wire [7:0] t_r40_c2_1;
  wire [7:0] t_r40_c2_2;
  wire [7:0] t_r40_c2_3;
  wire [7:0] t_r40_c2_4;
  wire [7:0] t_r40_c2_5;
  wire [7:0] t_r40_c2_6;
  wire [7:0] t_r40_c2_7;
  wire [7:0] t_r40_c2_8;
  wire [7:0] t_r40_c2_9;
  wire [7:0] t_r40_c2_10;
  wire [7:0] t_r40_c2_11;
  wire [7:0] t_r40_c2_12;
  wire [7:0] t_r40_c3_0;
  wire [7:0] t_r40_c3_1;
  wire [7:0] t_r40_c3_2;
  wire [7:0] t_r40_c3_3;
  wire [7:0] t_r40_c3_4;
  wire [7:0] t_r40_c3_5;
  wire [7:0] t_r40_c3_6;
  wire [7:0] t_r40_c3_7;
  wire [7:0] t_r40_c3_8;
  wire [7:0] t_r40_c3_9;
  wire [7:0] t_r40_c3_10;
  wire [7:0] t_r40_c3_11;
  wire [7:0] t_r40_c3_12;
  wire [7:0] t_r40_c4_0;
  wire [7:0] t_r40_c4_1;
  wire [7:0] t_r40_c4_2;
  wire [7:0] t_r40_c4_3;
  wire [7:0] t_r40_c4_4;
  wire [7:0] t_r40_c4_5;
  wire [7:0] t_r40_c4_6;
  wire [7:0] t_r40_c4_7;
  wire [7:0] t_r40_c4_8;
  wire [7:0] t_r40_c4_9;
  wire [7:0] t_r40_c4_10;
  wire [7:0] t_r40_c4_11;
  wire [7:0] t_r40_c4_12;
  wire [7:0] t_r40_c5_0;
  wire [7:0] t_r40_c5_1;
  wire [7:0] t_r40_c5_2;
  wire [7:0] t_r40_c5_3;
  wire [7:0] t_r40_c5_4;
  wire [7:0] t_r40_c5_5;
  wire [7:0] t_r40_c5_6;
  wire [7:0] t_r40_c5_7;
  wire [7:0] t_r40_c5_8;
  wire [7:0] t_r40_c5_9;
  wire [7:0] t_r40_c5_10;
  wire [7:0] t_r40_c5_11;
  wire [7:0] t_r40_c5_12;
  wire [7:0] t_r40_c6_0;
  wire [7:0] t_r40_c6_1;
  wire [7:0] t_r40_c6_2;
  wire [7:0] t_r40_c6_3;
  wire [7:0] t_r40_c6_4;
  wire [7:0] t_r40_c6_5;
  wire [7:0] t_r40_c6_6;
  wire [7:0] t_r40_c6_7;
  wire [7:0] t_r40_c6_8;
  wire [7:0] t_r40_c6_9;
  wire [7:0] t_r40_c6_10;
  wire [7:0] t_r40_c6_11;
  wire [7:0] t_r40_c6_12;
  wire [7:0] t_r40_c7_0;
  wire [7:0] t_r40_c7_1;
  wire [7:0] t_r40_c7_2;
  wire [7:0] t_r40_c7_3;
  wire [7:0] t_r40_c7_4;
  wire [7:0] t_r40_c7_5;
  wire [7:0] t_r40_c7_6;
  wire [7:0] t_r40_c7_7;
  wire [7:0] t_r40_c7_8;
  wire [7:0] t_r40_c7_9;
  wire [7:0] t_r40_c7_10;
  wire [7:0] t_r40_c7_11;
  wire [7:0] t_r40_c7_12;
  wire [7:0] t_r40_c8_0;
  wire [7:0] t_r40_c8_1;
  wire [7:0] t_r40_c8_2;
  wire [7:0] t_r40_c8_3;
  wire [7:0] t_r40_c8_4;
  wire [7:0] t_r40_c8_5;
  wire [7:0] t_r40_c8_6;
  wire [7:0] t_r40_c8_7;
  wire [7:0] t_r40_c8_8;
  wire [7:0] t_r40_c8_9;
  wire [7:0] t_r40_c8_10;
  wire [7:0] t_r40_c8_11;
  wire [7:0] t_r40_c8_12;
  wire [7:0] t_r40_c9_0;
  wire [7:0] t_r40_c9_1;
  wire [7:0] t_r40_c9_2;
  wire [7:0] t_r40_c9_3;
  wire [7:0] t_r40_c9_4;
  wire [7:0] t_r40_c9_5;
  wire [7:0] t_r40_c9_6;
  wire [7:0] t_r40_c9_7;
  wire [7:0] t_r40_c9_8;
  wire [7:0] t_r40_c9_9;
  wire [7:0] t_r40_c9_10;
  wire [7:0] t_r40_c9_11;
  wire [7:0] t_r40_c9_12;
  wire [7:0] t_r40_c10_0;
  wire [7:0] t_r40_c10_1;
  wire [7:0] t_r40_c10_2;
  wire [7:0] t_r40_c10_3;
  wire [7:0] t_r40_c10_4;
  wire [7:0] t_r40_c10_5;
  wire [7:0] t_r40_c10_6;
  wire [7:0] t_r40_c10_7;
  wire [7:0] t_r40_c10_8;
  wire [7:0] t_r40_c10_9;
  wire [7:0] t_r40_c10_10;
  wire [7:0] t_r40_c10_11;
  wire [7:0] t_r40_c10_12;
  wire [7:0] t_r40_c11_0;
  wire [7:0] t_r40_c11_1;
  wire [7:0] t_r40_c11_2;
  wire [7:0] t_r40_c11_3;
  wire [7:0] t_r40_c11_4;
  wire [7:0] t_r40_c11_5;
  wire [7:0] t_r40_c11_6;
  wire [7:0] t_r40_c11_7;
  wire [7:0] t_r40_c11_8;
  wire [7:0] t_r40_c11_9;
  wire [7:0] t_r40_c11_10;
  wire [7:0] t_r40_c11_11;
  wire [7:0] t_r40_c11_12;
  wire [7:0] t_r40_c12_0;
  wire [7:0] t_r40_c12_1;
  wire [7:0] t_r40_c12_2;
  wire [7:0] t_r40_c12_3;
  wire [7:0] t_r40_c12_4;
  wire [7:0] t_r40_c12_5;
  wire [7:0] t_r40_c12_6;
  wire [7:0] t_r40_c12_7;
  wire [7:0] t_r40_c12_8;
  wire [7:0] t_r40_c12_9;
  wire [7:0] t_r40_c12_10;
  wire [7:0] t_r40_c12_11;
  wire [7:0] t_r40_c12_12;
  wire [7:0] t_r40_c13_0;
  wire [7:0] t_r40_c13_1;
  wire [7:0] t_r40_c13_2;
  wire [7:0] t_r40_c13_3;
  wire [7:0] t_r40_c13_4;
  wire [7:0] t_r40_c13_5;
  wire [7:0] t_r40_c13_6;
  wire [7:0] t_r40_c13_7;
  wire [7:0] t_r40_c13_8;
  wire [7:0] t_r40_c13_9;
  wire [7:0] t_r40_c13_10;
  wire [7:0] t_r40_c13_11;
  wire [7:0] t_r40_c13_12;
  wire [7:0] t_r40_c14_0;
  wire [7:0] t_r40_c14_1;
  wire [7:0] t_r40_c14_2;
  wire [7:0] t_r40_c14_3;
  wire [7:0] t_r40_c14_4;
  wire [7:0] t_r40_c14_5;
  wire [7:0] t_r40_c14_6;
  wire [7:0] t_r40_c14_7;
  wire [7:0] t_r40_c14_8;
  wire [7:0] t_r40_c14_9;
  wire [7:0] t_r40_c14_10;
  wire [7:0] t_r40_c14_11;
  wire [7:0] t_r40_c14_12;
  wire [7:0] t_r40_c15_0;
  wire [7:0] t_r40_c15_1;
  wire [7:0] t_r40_c15_2;
  wire [7:0] t_r40_c15_3;
  wire [7:0] t_r40_c15_4;
  wire [7:0] t_r40_c15_5;
  wire [7:0] t_r40_c15_6;
  wire [7:0] t_r40_c15_7;
  wire [7:0] t_r40_c15_8;
  wire [7:0] t_r40_c15_9;
  wire [7:0] t_r40_c15_10;
  wire [7:0] t_r40_c15_11;
  wire [7:0] t_r40_c15_12;
  wire [7:0] t_r40_c16_0;
  wire [7:0] t_r40_c16_1;
  wire [7:0] t_r40_c16_2;
  wire [7:0] t_r40_c16_3;
  wire [7:0] t_r40_c16_4;
  wire [7:0] t_r40_c16_5;
  wire [7:0] t_r40_c16_6;
  wire [7:0] t_r40_c16_7;
  wire [7:0] t_r40_c16_8;
  wire [7:0] t_r40_c16_9;
  wire [7:0] t_r40_c16_10;
  wire [7:0] t_r40_c16_11;
  wire [7:0] t_r40_c16_12;
  wire [7:0] t_r40_c17_0;
  wire [7:0] t_r40_c17_1;
  wire [7:0] t_r40_c17_2;
  wire [7:0] t_r40_c17_3;
  wire [7:0] t_r40_c17_4;
  wire [7:0] t_r40_c17_5;
  wire [7:0] t_r40_c17_6;
  wire [7:0] t_r40_c17_7;
  wire [7:0] t_r40_c17_8;
  wire [7:0] t_r40_c17_9;
  wire [7:0] t_r40_c17_10;
  wire [7:0] t_r40_c17_11;
  wire [7:0] t_r40_c17_12;
  wire [7:0] t_r40_c18_0;
  wire [7:0] t_r40_c18_1;
  wire [7:0] t_r40_c18_2;
  wire [7:0] t_r40_c18_3;
  wire [7:0] t_r40_c18_4;
  wire [7:0] t_r40_c18_5;
  wire [7:0] t_r40_c18_6;
  wire [7:0] t_r40_c18_7;
  wire [7:0] t_r40_c18_8;
  wire [7:0] t_r40_c18_9;
  wire [7:0] t_r40_c18_10;
  wire [7:0] t_r40_c18_11;
  wire [7:0] t_r40_c18_12;
  wire [7:0] t_r40_c19_0;
  wire [7:0] t_r40_c19_1;
  wire [7:0] t_r40_c19_2;
  wire [7:0] t_r40_c19_3;
  wire [7:0] t_r40_c19_4;
  wire [7:0] t_r40_c19_5;
  wire [7:0] t_r40_c19_6;
  wire [7:0] t_r40_c19_7;
  wire [7:0] t_r40_c19_8;
  wire [7:0] t_r40_c19_9;
  wire [7:0] t_r40_c19_10;
  wire [7:0] t_r40_c19_11;
  wire [7:0] t_r40_c19_12;
  wire [7:0] t_r40_c20_0;
  wire [7:0] t_r40_c20_1;
  wire [7:0] t_r40_c20_2;
  wire [7:0] t_r40_c20_3;
  wire [7:0] t_r40_c20_4;
  wire [7:0] t_r40_c20_5;
  wire [7:0] t_r40_c20_6;
  wire [7:0] t_r40_c20_7;
  wire [7:0] t_r40_c20_8;
  wire [7:0] t_r40_c20_9;
  wire [7:0] t_r40_c20_10;
  wire [7:0] t_r40_c20_11;
  wire [7:0] t_r40_c20_12;
  wire [7:0] t_r40_c21_0;
  wire [7:0] t_r40_c21_1;
  wire [7:0] t_r40_c21_2;
  wire [7:0] t_r40_c21_3;
  wire [7:0] t_r40_c21_4;
  wire [7:0] t_r40_c21_5;
  wire [7:0] t_r40_c21_6;
  wire [7:0] t_r40_c21_7;
  wire [7:0] t_r40_c21_8;
  wire [7:0] t_r40_c21_9;
  wire [7:0] t_r40_c21_10;
  wire [7:0] t_r40_c21_11;
  wire [7:0] t_r40_c21_12;
  wire [7:0] t_r40_c22_0;
  wire [7:0] t_r40_c22_1;
  wire [7:0] t_r40_c22_2;
  wire [7:0] t_r40_c22_3;
  wire [7:0] t_r40_c22_4;
  wire [7:0] t_r40_c22_5;
  wire [7:0] t_r40_c22_6;
  wire [7:0] t_r40_c22_7;
  wire [7:0] t_r40_c22_8;
  wire [7:0] t_r40_c22_9;
  wire [7:0] t_r40_c22_10;
  wire [7:0] t_r40_c22_11;
  wire [7:0] t_r40_c22_12;
  wire [7:0] t_r40_c23_0;
  wire [7:0] t_r40_c23_1;
  wire [7:0] t_r40_c23_2;
  wire [7:0] t_r40_c23_3;
  wire [7:0] t_r40_c23_4;
  wire [7:0] t_r40_c23_5;
  wire [7:0] t_r40_c23_6;
  wire [7:0] t_r40_c23_7;
  wire [7:0] t_r40_c23_8;
  wire [7:0] t_r40_c23_9;
  wire [7:0] t_r40_c23_10;
  wire [7:0] t_r40_c23_11;
  wire [7:0] t_r40_c23_12;
  wire [7:0] t_r40_c24_0;
  wire [7:0] t_r40_c24_1;
  wire [7:0] t_r40_c24_2;
  wire [7:0] t_r40_c24_3;
  wire [7:0] t_r40_c24_4;
  wire [7:0] t_r40_c24_5;
  wire [7:0] t_r40_c24_6;
  wire [7:0] t_r40_c24_7;
  wire [7:0] t_r40_c24_8;
  wire [7:0] t_r40_c24_9;
  wire [7:0] t_r40_c24_10;
  wire [7:0] t_r40_c24_11;
  wire [7:0] t_r40_c24_12;
  wire [7:0] t_r40_c25_0;
  wire [7:0] t_r40_c25_1;
  wire [7:0] t_r40_c25_2;
  wire [7:0] t_r40_c25_3;
  wire [7:0] t_r40_c25_4;
  wire [7:0] t_r40_c25_5;
  wire [7:0] t_r40_c25_6;
  wire [7:0] t_r40_c25_7;
  wire [7:0] t_r40_c25_8;
  wire [7:0] t_r40_c25_9;
  wire [7:0] t_r40_c25_10;
  wire [7:0] t_r40_c25_11;
  wire [7:0] t_r40_c25_12;
  wire [7:0] t_r40_c26_0;
  wire [7:0] t_r40_c26_1;
  wire [7:0] t_r40_c26_2;
  wire [7:0] t_r40_c26_3;
  wire [7:0] t_r40_c26_4;
  wire [7:0] t_r40_c26_5;
  wire [7:0] t_r40_c26_6;
  wire [7:0] t_r40_c26_7;
  wire [7:0] t_r40_c26_8;
  wire [7:0] t_r40_c26_9;
  wire [7:0] t_r40_c26_10;
  wire [7:0] t_r40_c26_11;
  wire [7:0] t_r40_c26_12;
  wire [7:0] t_r40_c27_0;
  wire [7:0] t_r40_c27_1;
  wire [7:0] t_r40_c27_2;
  wire [7:0] t_r40_c27_3;
  wire [7:0] t_r40_c27_4;
  wire [7:0] t_r40_c27_5;
  wire [7:0] t_r40_c27_6;
  wire [7:0] t_r40_c27_7;
  wire [7:0] t_r40_c27_8;
  wire [7:0] t_r40_c27_9;
  wire [7:0] t_r40_c27_10;
  wire [7:0] t_r40_c27_11;
  wire [7:0] t_r40_c27_12;
  wire [7:0] t_r40_c28_0;
  wire [7:0] t_r40_c28_1;
  wire [7:0] t_r40_c28_2;
  wire [7:0] t_r40_c28_3;
  wire [7:0] t_r40_c28_4;
  wire [7:0] t_r40_c28_5;
  wire [7:0] t_r40_c28_6;
  wire [7:0] t_r40_c28_7;
  wire [7:0] t_r40_c28_8;
  wire [7:0] t_r40_c28_9;
  wire [7:0] t_r40_c28_10;
  wire [7:0] t_r40_c28_11;
  wire [7:0] t_r40_c28_12;
  wire [7:0] t_r40_c29_0;
  wire [7:0] t_r40_c29_1;
  wire [7:0] t_r40_c29_2;
  wire [7:0] t_r40_c29_3;
  wire [7:0] t_r40_c29_4;
  wire [7:0] t_r40_c29_5;
  wire [7:0] t_r40_c29_6;
  wire [7:0] t_r40_c29_7;
  wire [7:0] t_r40_c29_8;
  wire [7:0] t_r40_c29_9;
  wire [7:0] t_r40_c29_10;
  wire [7:0] t_r40_c29_11;
  wire [7:0] t_r40_c29_12;
  wire [7:0] t_r40_c30_0;
  wire [7:0] t_r40_c30_1;
  wire [7:0] t_r40_c30_2;
  wire [7:0] t_r40_c30_3;
  wire [7:0] t_r40_c30_4;
  wire [7:0] t_r40_c30_5;
  wire [7:0] t_r40_c30_6;
  wire [7:0] t_r40_c30_7;
  wire [7:0] t_r40_c30_8;
  wire [7:0] t_r40_c30_9;
  wire [7:0] t_r40_c30_10;
  wire [7:0] t_r40_c30_11;
  wire [7:0] t_r40_c30_12;
  wire [7:0] t_r40_c31_0;
  wire [7:0] t_r40_c31_1;
  wire [7:0] t_r40_c31_2;
  wire [7:0] t_r40_c31_3;
  wire [7:0] t_r40_c31_4;
  wire [7:0] t_r40_c31_5;
  wire [7:0] t_r40_c31_6;
  wire [7:0] t_r40_c31_7;
  wire [7:0] t_r40_c31_8;
  wire [7:0] t_r40_c31_9;
  wire [7:0] t_r40_c31_10;
  wire [7:0] t_r40_c31_11;
  wire [7:0] t_r40_c31_12;
  wire [7:0] t_r40_c32_0;
  wire [7:0] t_r40_c32_1;
  wire [7:0] t_r40_c32_2;
  wire [7:0] t_r40_c32_3;
  wire [7:0] t_r40_c32_4;
  wire [7:0] t_r40_c32_5;
  wire [7:0] t_r40_c32_6;
  wire [7:0] t_r40_c32_7;
  wire [7:0] t_r40_c32_8;
  wire [7:0] t_r40_c32_9;
  wire [7:0] t_r40_c32_10;
  wire [7:0] t_r40_c32_11;
  wire [7:0] t_r40_c32_12;
  wire [7:0] t_r40_c33_0;
  wire [7:0] t_r40_c33_1;
  wire [7:0] t_r40_c33_2;
  wire [7:0] t_r40_c33_3;
  wire [7:0] t_r40_c33_4;
  wire [7:0] t_r40_c33_5;
  wire [7:0] t_r40_c33_6;
  wire [7:0] t_r40_c33_7;
  wire [7:0] t_r40_c33_8;
  wire [7:0] t_r40_c33_9;
  wire [7:0] t_r40_c33_10;
  wire [7:0] t_r40_c33_11;
  wire [7:0] t_r40_c33_12;
  wire [7:0] t_r40_c34_0;
  wire [7:0] t_r40_c34_1;
  wire [7:0] t_r40_c34_2;
  wire [7:0] t_r40_c34_3;
  wire [7:0] t_r40_c34_4;
  wire [7:0] t_r40_c34_5;
  wire [7:0] t_r40_c34_6;
  wire [7:0] t_r40_c34_7;
  wire [7:0] t_r40_c34_8;
  wire [7:0] t_r40_c34_9;
  wire [7:0] t_r40_c34_10;
  wire [7:0] t_r40_c34_11;
  wire [7:0] t_r40_c34_12;
  wire [7:0] t_r40_c35_0;
  wire [7:0] t_r40_c35_1;
  wire [7:0] t_r40_c35_2;
  wire [7:0] t_r40_c35_3;
  wire [7:0] t_r40_c35_4;
  wire [7:0] t_r40_c35_5;
  wire [7:0] t_r40_c35_6;
  wire [7:0] t_r40_c35_7;
  wire [7:0] t_r40_c35_8;
  wire [7:0] t_r40_c35_9;
  wire [7:0] t_r40_c35_10;
  wire [7:0] t_r40_c35_11;
  wire [7:0] t_r40_c35_12;
  wire [7:0] t_r40_c36_0;
  wire [7:0] t_r40_c36_1;
  wire [7:0] t_r40_c36_2;
  wire [7:0] t_r40_c36_3;
  wire [7:0] t_r40_c36_4;
  wire [7:0] t_r40_c36_5;
  wire [7:0] t_r40_c36_6;
  wire [7:0] t_r40_c36_7;
  wire [7:0] t_r40_c36_8;
  wire [7:0] t_r40_c36_9;
  wire [7:0] t_r40_c36_10;
  wire [7:0] t_r40_c36_11;
  wire [7:0] t_r40_c36_12;
  wire [7:0] t_r40_c37_0;
  wire [7:0] t_r40_c37_1;
  wire [7:0] t_r40_c37_2;
  wire [7:0] t_r40_c37_3;
  wire [7:0] t_r40_c37_4;
  wire [7:0] t_r40_c37_5;
  wire [7:0] t_r40_c37_6;
  wire [7:0] t_r40_c37_7;
  wire [7:0] t_r40_c37_8;
  wire [7:0] t_r40_c37_9;
  wire [7:0] t_r40_c37_10;
  wire [7:0] t_r40_c37_11;
  wire [7:0] t_r40_c37_12;
  wire [7:0] t_r40_c38_0;
  wire [7:0] t_r40_c38_1;
  wire [7:0] t_r40_c38_2;
  wire [7:0] t_r40_c38_3;
  wire [7:0] t_r40_c38_4;
  wire [7:0] t_r40_c38_5;
  wire [7:0] t_r40_c38_6;
  wire [7:0] t_r40_c38_7;
  wire [7:0] t_r40_c38_8;
  wire [7:0] t_r40_c38_9;
  wire [7:0] t_r40_c38_10;
  wire [7:0] t_r40_c38_11;
  wire [7:0] t_r40_c38_12;
  wire [7:0] t_r40_c39_0;
  wire [7:0] t_r40_c39_1;
  wire [7:0] t_r40_c39_2;
  wire [7:0] t_r40_c39_3;
  wire [7:0] t_r40_c39_4;
  wire [7:0] t_r40_c39_5;
  wire [7:0] t_r40_c39_6;
  wire [7:0] t_r40_c39_7;
  wire [7:0] t_r40_c39_8;
  wire [7:0] t_r40_c39_9;
  wire [7:0] t_r40_c39_10;
  wire [7:0] t_r40_c39_11;
  wire [7:0] t_r40_c39_12;
  wire [7:0] t_r40_c40_0;
  wire [7:0] t_r40_c40_1;
  wire [7:0] t_r40_c40_2;
  wire [7:0] t_r40_c40_3;
  wire [7:0] t_r40_c40_4;
  wire [7:0] t_r40_c40_5;
  wire [7:0] t_r40_c40_6;
  wire [7:0] t_r40_c40_7;
  wire [7:0] t_r40_c40_8;
  wire [7:0] t_r40_c40_9;
  wire [7:0] t_r40_c40_10;
  wire [7:0] t_r40_c40_11;
  wire [7:0] t_r40_c40_12;
  wire [7:0] t_r40_c41_0;
  wire [7:0] t_r40_c41_1;
  wire [7:0] t_r40_c41_2;
  wire [7:0] t_r40_c41_3;
  wire [7:0] t_r40_c41_4;
  wire [7:0] t_r40_c41_5;
  wire [7:0] t_r40_c41_6;
  wire [7:0] t_r40_c41_7;
  wire [7:0] t_r40_c41_8;
  wire [7:0] t_r40_c41_9;
  wire [7:0] t_r40_c41_10;
  wire [7:0] t_r40_c41_11;
  wire [7:0] t_r40_c41_12;
  wire [7:0] t_r40_c42_0;
  wire [7:0] t_r40_c42_1;
  wire [7:0] t_r40_c42_2;
  wire [7:0] t_r40_c42_3;
  wire [7:0] t_r40_c42_4;
  wire [7:0] t_r40_c42_5;
  wire [7:0] t_r40_c42_6;
  wire [7:0] t_r40_c42_7;
  wire [7:0] t_r40_c42_8;
  wire [7:0] t_r40_c42_9;
  wire [7:0] t_r40_c42_10;
  wire [7:0] t_r40_c42_11;
  wire [7:0] t_r40_c42_12;
  wire [7:0] t_r40_c43_0;
  wire [7:0] t_r40_c43_1;
  wire [7:0] t_r40_c43_2;
  wire [7:0] t_r40_c43_3;
  wire [7:0] t_r40_c43_4;
  wire [7:0] t_r40_c43_5;
  wire [7:0] t_r40_c43_6;
  wire [7:0] t_r40_c43_7;
  wire [7:0] t_r40_c43_8;
  wire [7:0] t_r40_c43_9;
  wire [7:0] t_r40_c43_10;
  wire [7:0] t_r40_c43_11;
  wire [7:0] t_r40_c43_12;
  wire [7:0] t_r40_c44_0;
  wire [7:0] t_r40_c44_1;
  wire [7:0] t_r40_c44_2;
  wire [7:0] t_r40_c44_3;
  wire [7:0] t_r40_c44_4;
  wire [7:0] t_r40_c44_5;
  wire [7:0] t_r40_c44_6;
  wire [7:0] t_r40_c44_7;
  wire [7:0] t_r40_c44_8;
  wire [7:0] t_r40_c44_9;
  wire [7:0] t_r40_c44_10;
  wire [7:0] t_r40_c44_11;
  wire [7:0] t_r40_c44_12;
  wire [7:0] t_r40_c45_0;
  wire [7:0] t_r40_c45_1;
  wire [7:0] t_r40_c45_2;
  wire [7:0] t_r40_c45_3;
  wire [7:0] t_r40_c45_4;
  wire [7:0] t_r40_c45_5;
  wire [7:0] t_r40_c45_6;
  wire [7:0] t_r40_c45_7;
  wire [7:0] t_r40_c45_8;
  wire [7:0] t_r40_c45_9;
  wire [7:0] t_r40_c45_10;
  wire [7:0] t_r40_c45_11;
  wire [7:0] t_r40_c45_12;
  wire [7:0] t_r40_c46_0;
  wire [7:0] t_r40_c46_1;
  wire [7:0] t_r40_c46_2;
  wire [7:0] t_r40_c46_3;
  wire [7:0] t_r40_c46_4;
  wire [7:0] t_r40_c46_5;
  wire [7:0] t_r40_c46_6;
  wire [7:0] t_r40_c46_7;
  wire [7:0] t_r40_c46_8;
  wire [7:0] t_r40_c46_9;
  wire [7:0] t_r40_c46_10;
  wire [7:0] t_r40_c46_11;
  wire [7:0] t_r40_c46_12;
  wire [7:0] t_r40_c47_0;
  wire [7:0] t_r40_c47_1;
  wire [7:0] t_r40_c47_2;
  wire [7:0] t_r40_c47_3;
  wire [7:0] t_r40_c47_4;
  wire [7:0] t_r40_c47_5;
  wire [7:0] t_r40_c47_6;
  wire [7:0] t_r40_c47_7;
  wire [7:0] t_r40_c47_8;
  wire [7:0] t_r40_c47_9;
  wire [7:0] t_r40_c47_10;
  wire [7:0] t_r40_c47_11;
  wire [7:0] t_r40_c47_12;
  wire [7:0] t_r40_c48_0;
  wire [7:0] t_r40_c48_1;
  wire [7:0] t_r40_c48_2;
  wire [7:0] t_r40_c48_3;
  wire [7:0] t_r40_c48_4;
  wire [7:0] t_r40_c48_5;
  wire [7:0] t_r40_c48_6;
  wire [7:0] t_r40_c48_7;
  wire [7:0] t_r40_c48_8;
  wire [7:0] t_r40_c48_9;
  wire [7:0] t_r40_c48_10;
  wire [7:0] t_r40_c48_11;
  wire [7:0] t_r40_c48_12;
  wire [7:0] t_r40_c49_0;
  wire [7:0] t_r40_c49_1;
  wire [7:0] t_r40_c49_2;
  wire [7:0] t_r40_c49_3;
  wire [7:0] t_r40_c49_4;
  wire [7:0] t_r40_c49_5;
  wire [7:0] t_r40_c49_6;
  wire [7:0] t_r40_c49_7;
  wire [7:0] t_r40_c49_8;
  wire [7:0] t_r40_c49_9;
  wire [7:0] t_r40_c49_10;
  wire [7:0] t_r40_c49_11;
  wire [7:0] t_r40_c49_12;
  wire [7:0] t_r40_c50_0;
  wire [7:0] t_r40_c50_1;
  wire [7:0] t_r40_c50_2;
  wire [7:0] t_r40_c50_3;
  wire [7:0] t_r40_c50_4;
  wire [7:0] t_r40_c50_5;
  wire [7:0] t_r40_c50_6;
  wire [7:0] t_r40_c50_7;
  wire [7:0] t_r40_c50_8;
  wire [7:0] t_r40_c50_9;
  wire [7:0] t_r40_c50_10;
  wire [7:0] t_r40_c50_11;
  wire [7:0] t_r40_c50_12;
  wire [7:0] t_r40_c51_0;
  wire [7:0] t_r40_c51_1;
  wire [7:0] t_r40_c51_2;
  wire [7:0] t_r40_c51_3;
  wire [7:0] t_r40_c51_4;
  wire [7:0] t_r40_c51_5;
  wire [7:0] t_r40_c51_6;
  wire [7:0] t_r40_c51_7;
  wire [7:0] t_r40_c51_8;
  wire [7:0] t_r40_c51_9;
  wire [7:0] t_r40_c51_10;
  wire [7:0] t_r40_c51_11;
  wire [7:0] t_r40_c51_12;
  wire [7:0] t_r40_c52_0;
  wire [7:0] t_r40_c52_1;
  wire [7:0] t_r40_c52_2;
  wire [7:0] t_r40_c52_3;
  wire [7:0] t_r40_c52_4;
  wire [7:0] t_r40_c52_5;
  wire [7:0] t_r40_c52_6;
  wire [7:0] t_r40_c52_7;
  wire [7:0] t_r40_c52_8;
  wire [7:0] t_r40_c52_9;
  wire [7:0] t_r40_c52_10;
  wire [7:0] t_r40_c52_11;
  wire [7:0] t_r40_c52_12;
  wire [7:0] t_r40_c53_0;
  wire [7:0] t_r40_c53_1;
  wire [7:0] t_r40_c53_2;
  wire [7:0] t_r40_c53_3;
  wire [7:0] t_r40_c53_4;
  wire [7:0] t_r40_c53_5;
  wire [7:0] t_r40_c53_6;
  wire [7:0] t_r40_c53_7;
  wire [7:0] t_r40_c53_8;
  wire [7:0] t_r40_c53_9;
  wire [7:0] t_r40_c53_10;
  wire [7:0] t_r40_c53_11;
  wire [7:0] t_r40_c53_12;
  wire [7:0] t_r40_c54_0;
  wire [7:0] t_r40_c54_1;
  wire [7:0] t_r40_c54_2;
  wire [7:0] t_r40_c54_3;
  wire [7:0] t_r40_c54_4;
  wire [7:0] t_r40_c54_5;
  wire [7:0] t_r40_c54_6;
  wire [7:0] t_r40_c54_7;
  wire [7:0] t_r40_c54_8;
  wire [7:0] t_r40_c54_9;
  wire [7:0] t_r40_c54_10;
  wire [7:0] t_r40_c54_11;
  wire [7:0] t_r40_c54_12;
  wire [7:0] t_r40_c55_0;
  wire [7:0] t_r40_c55_1;
  wire [7:0] t_r40_c55_2;
  wire [7:0] t_r40_c55_3;
  wire [7:0] t_r40_c55_4;
  wire [7:0] t_r40_c55_5;
  wire [7:0] t_r40_c55_6;
  wire [7:0] t_r40_c55_7;
  wire [7:0] t_r40_c55_8;
  wire [7:0] t_r40_c55_9;
  wire [7:0] t_r40_c55_10;
  wire [7:0] t_r40_c55_11;
  wire [7:0] t_r40_c55_12;
  wire [7:0] t_r40_c56_0;
  wire [7:0] t_r40_c56_1;
  wire [7:0] t_r40_c56_2;
  wire [7:0] t_r40_c56_3;
  wire [7:0] t_r40_c56_4;
  wire [7:0] t_r40_c56_5;
  wire [7:0] t_r40_c56_6;
  wire [7:0] t_r40_c56_7;
  wire [7:0] t_r40_c56_8;
  wire [7:0] t_r40_c56_9;
  wire [7:0] t_r40_c56_10;
  wire [7:0] t_r40_c56_11;
  wire [7:0] t_r40_c56_12;
  wire [7:0] t_r40_c57_0;
  wire [7:0] t_r40_c57_1;
  wire [7:0] t_r40_c57_2;
  wire [7:0] t_r40_c57_3;
  wire [7:0] t_r40_c57_4;
  wire [7:0] t_r40_c57_5;
  wire [7:0] t_r40_c57_6;
  wire [7:0] t_r40_c57_7;
  wire [7:0] t_r40_c57_8;
  wire [7:0] t_r40_c57_9;
  wire [7:0] t_r40_c57_10;
  wire [7:0] t_r40_c57_11;
  wire [7:0] t_r40_c57_12;
  wire [7:0] t_r40_c58_0;
  wire [7:0] t_r40_c58_1;
  wire [7:0] t_r40_c58_2;
  wire [7:0] t_r40_c58_3;
  wire [7:0] t_r40_c58_4;
  wire [7:0] t_r40_c58_5;
  wire [7:0] t_r40_c58_6;
  wire [7:0] t_r40_c58_7;
  wire [7:0] t_r40_c58_8;
  wire [7:0] t_r40_c58_9;
  wire [7:0] t_r40_c58_10;
  wire [7:0] t_r40_c58_11;
  wire [7:0] t_r40_c58_12;
  wire [7:0] t_r40_c59_0;
  wire [7:0] t_r40_c59_1;
  wire [7:0] t_r40_c59_2;
  wire [7:0] t_r40_c59_3;
  wire [7:0] t_r40_c59_4;
  wire [7:0] t_r40_c59_5;
  wire [7:0] t_r40_c59_6;
  wire [7:0] t_r40_c59_7;
  wire [7:0] t_r40_c59_8;
  wire [7:0] t_r40_c59_9;
  wire [7:0] t_r40_c59_10;
  wire [7:0] t_r40_c59_11;
  wire [7:0] t_r40_c59_12;
  wire [7:0] t_r40_c60_0;
  wire [7:0] t_r40_c60_1;
  wire [7:0] t_r40_c60_2;
  wire [7:0] t_r40_c60_3;
  wire [7:0] t_r40_c60_4;
  wire [7:0] t_r40_c60_5;
  wire [7:0] t_r40_c60_6;
  wire [7:0] t_r40_c60_7;
  wire [7:0] t_r40_c60_8;
  wire [7:0] t_r40_c60_9;
  wire [7:0] t_r40_c60_10;
  wire [7:0] t_r40_c60_11;
  wire [7:0] t_r40_c60_12;
  wire [7:0] t_r40_c61_0;
  wire [7:0] t_r40_c61_1;
  wire [7:0] t_r40_c61_2;
  wire [7:0] t_r40_c61_3;
  wire [7:0] t_r40_c61_4;
  wire [7:0] t_r40_c61_5;
  wire [7:0] t_r40_c61_6;
  wire [7:0] t_r40_c61_7;
  wire [7:0] t_r40_c61_8;
  wire [7:0] t_r40_c61_9;
  wire [7:0] t_r40_c61_10;
  wire [7:0] t_r40_c61_11;
  wire [7:0] t_r40_c61_12;
  wire [7:0] t_r40_c62_0;
  wire [7:0] t_r40_c62_1;
  wire [7:0] t_r40_c62_2;
  wire [7:0] t_r40_c62_3;
  wire [7:0] t_r40_c62_4;
  wire [7:0] t_r40_c62_5;
  wire [7:0] t_r40_c62_6;
  wire [7:0] t_r40_c62_7;
  wire [7:0] t_r40_c62_8;
  wire [7:0] t_r40_c62_9;
  wire [7:0] t_r40_c62_10;
  wire [7:0] t_r40_c62_11;
  wire [7:0] t_r40_c62_12;
  wire [7:0] t_r40_c63_0;
  wire [7:0] t_r40_c63_1;
  wire [7:0] t_r40_c63_2;
  wire [7:0] t_r40_c63_3;
  wire [7:0] t_r40_c63_4;
  wire [7:0] t_r40_c63_5;
  wire [7:0] t_r40_c63_6;
  wire [7:0] t_r40_c63_7;
  wire [7:0] t_r40_c63_8;
  wire [7:0] t_r40_c63_9;
  wire [7:0] t_r40_c63_10;
  wire [7:0] t_r40_c63_11;
  wire [7:0] t_r40_c63_12;
  wire [7:0] t_r40_c64_0;
  wire [7:0] t_r40_c64_1;
  wire [7:0] t_r40_c64_2;
  wire [7:0] t_r40_c64_3;
  wire [7:0] t_r40_c64_4;
  wire [7:0] t_r40_c64_5;
  wire [7:0] t_r40_c64_6;
  wire [7:0] t_r40_c64_7;
  wire [7:0] t_r40_c64_8;
  wire [7:0] t_r40_c64_9;
  wire [7:0] t_r40_c64_10;
  wire [7:0] t_r40_c64_11;
  wire [7:0] t_r40_c64_12;
  wire [7:0] t_r40_c65_0;
  wire [7:0] t_r40_c65_1;
  wire [7:0] t_r40_c65_2;
  wire [7:0] t_r40_c65_3;
  wire [7:0] t_r40_c65_4;
  wire [7:0] t_r40_c65_5;
  wire [7:0] t_r40_c65_6;
  wire [7:0] t_r40_c65_7;
  wire [7:0] t_r40_c65_8;
  wire [7:0] t_r40_c65_9;
  wire [7:0] t_r40_c65_10;
  wire [7:0] t_r40_c65_11;
  wire [7:0] t_r40_c65_12;
  wire [7:0] t_r41_c0_0;
  wire [7:0] t_r41_c0_1;
  wire [7:0] t_r41_c0_2;
  wire [7:0] t_r41_c0_3;
  wire [7:0] t_r41_c0_4;
  wire [7:0] t_r41_c0_5;
  wire [7:0] t_r41_c0_6;
  wire [7:0] t_r41_c0_7;
  wire [7:0] t_r41_c0_8;
  wire [7:0] t_r41_c0_9;
  wire [7:0] t_r41_c0_10;
  wire [7:0] t_r41_c0_11;
  wire [7:0] t_r41_c0_12;
  wire [7:0] t_r41_c1_0;
  wire [7:0] t_r41_c1_1;
  wire [7:0] t_r41_c1_2;
  wire [7:0] t_r41_c1_3;
  wire [7:0] t_r41_c1_4;
  wire [7:0] t_r41_c1_5;
  wire [7:0] t_r41_c1_6;
  wire [7:0] t_r41_c1_7;
  wire [7:0] t_r41_c1_8;
  wire [7:0] t_r41_c1_9;
  wire [7:0] t_r41_c1_10;
  wire [7:0] t_r41_c1_11;
  wire [7:0] t_r41_c1_12;
  wire [7:0] t_r41_c2_0;
  wire [7:0] t_r41_c2_1;
  wire [7:0] t_r41_c2_2;
  wire [7:0] t_r41_c2_3;
  wire [7:0] t_r41_c2_4;
  wire [7:0] t_r41_c2_5;
  wire [7:0] t_r41_c2_6;
  wire [7:0] t_r41_c2_7;
  wire [7:0] t_r41_c2_8;
  wire [7:0] t_r41_c2_9;
  wire [7:0] t_r41_c2_10;
  wire [7:0] t_r41_c2_11;
  wire [7:0] t_r41_c2_12;
  wire [7:0] t_r41_c3_0;
  wire [7:0] t_r41_c3_1;
  wire [7:0] t_r41_c3_2;
  wire [7:0] t_r41_c3_3;
  wire [7:0] t_r41_c3_4;
  wire [7:0] t_r41_c3_5;
  wire [7:0] t_r41_c3_6;
  wire [7:0] t_r41_c3_7;
  wire [7:0] t_r41_c3_8;
  wire [7:0] t_r41_c3_9;
  wire [7:0] t_r41_c3_10;
  wire [7:0] t_r41_c3_11;
  wire [7:0] t_r41_c3_12;
  wire [7:0] t_r41_c4_0;
  wire [7:0] t_r41_c4_1;
  wire [7:0] t_r41_c4_2;
  wire [7:0] t_r41_c4_3;
  wire [7:0] t_r41_c4_4;
  wire [7:0] t_r41_c4_5;
  wire [7:0] t_r41_c4_6;
  wire [7:0] t_r41_c4_7;
  wire [7:0] t_r41_c4_8;
  wire [7:0] t_r41_c4_9;
  wire [7:0] t_r41_c4_10;
  wire [7:0] t_r41_c4_11;
  wire [7:0] t_r41_c4_12;
  wire [7:0] t_r41_c5_0;
  wire [7:0] t_r41_c5_1;
  wire [7:0] t_r41_c5_2;
  wire [7:0] t_r41_c5_3;
  wire [7:0] t_r41_c5_4;
  wire [7:0] t_r41_c5_5;
  wire [7:0] t_r41_c5_6;
  wire [7:0] t_r41_c5_7;
  wire [7:0] t_r41_c5_8;
  wire [7:0] t_r41_c5_9;
  wire [7:0] t_r41_c5_10;
  wire [7:0] t_r41_c5_11;
  wire [7:0] t_r41_c5_12;
  wire [7:0] t_r41_c6_0;
  wire [7:0] t_r41_c6_1;
  wire [7:0] t_r41_c6_2;
  wire [7:0] t_r41_c6_3;
  wire [7:0] t_r41_c6_4;
  wire [7:0] t_r41_c6_5;
  wire [7:0] t_r41_c6_6;
  wire [7:0] t_r41_c6_7;
  wire [7:0] t_r41_c6_8;
  wire [7:0] t_r41_c6_9;
  wire [7:0] t_r41_c6_10;
  wire [7:0] t_r41_c6_11;
  wire [7:0] t_r41_c6_12;
  wire [7:0] t_r41_c7_0;
  wire [7:0] t_r41_c7_1;
  wire [7:0] t_r41_c7_2;
  wire [7:0] t_r41_c7_3;
  wire [7:0] t_r41_c7_4;
  wire [7:0] t_r41_c7_5;
  wire [7:0] t_r41_c7_6;
  wire [7:0] t_r41_c7_7;
  wire [7:0] t_r41_c7_8;
  wire [7:0] t_r41_c7_9;
  wire [7:0] t_r41_c7_10;
  wire [7:0] t_r41_c7_11;
  wire [7:0] t_r41_c7_12;
  wire [7:0] t_r41_c8_0;
  wire [7:0] t_r41_c8_1;
  wire [7:0] t_r41_c8_2;
  wire [7:0] t_r41_c8_3;
  wire [7:0] t_r41_c8_4;
  wire [7:0] t_r41_c8_5;
  wire [7:0] t_r41_c8_6;
  wire [7:0] t_r41_c8_7;
  wire [7:0] t_r41_c8_8;
  wire [7:0] t_r41_c8_9;
  wire [7:0] t_r41_c8_10;
  wire [7:0] t_r41_c8_11;
  wire [7:0] t_r41_c8_12;
  wire [7:0] t_r41_c9_0;
  wire [7:0] t_r41_c9_1;
  wire [7:0] t_r41_c9_2;
  wire [7:0] t_r41_c9_3;
  wire [7:0] t_r41_c9_4;
  wire [7:0] t_r41_c9_5;
  wire [7:0] t_r41_c9_6;
  wire [7:0] t_r41_c9_7;
  wire [7:0] t_r41_c9_8;
  wire [7:0] t_r41_c9_9;
  wire [7:0] t_r41_c9_10;
  wire [7:0] t_r41_c9_11;
  wire [7:0] t_r41_c9_12;
  wire [7:0] t_r41_c10_0;
  wire [7:0] t_r41_c10_1;
  wire [7:0] t_r41_c10_2;
  wire [7:0] t_r41_c10_3;
  wire [7:0] t_r41_c10_4;
  wire [7:0] t_r41_c10_5;
  wire [7:0] t_r41_c10_6;
  wire [7:0] t_r41_c10_7;
  wire [7:0] t_r41_c10_8;
  wire [7:0] t_r41_c10_9;
  wire [7:0] t_r41_c10_10;
  wire [7:0] t_r41_c10_11;
  wire [7:0] t_r41_c10_12;
  wire [7:0] t_r41_c11_0;
  wire [7:0] t_r41_c11_1;
  wire [7:0] t_r41_c11_2;
  wire [7:0] t_r41_c11_3;
  wire [7:0] t_r41_c11_4;
  wire [7:0] t_r41_c11_5;
  wire [7:0] t_r41_c11_6;
  wire [7:0] t_r41_c11_7;
  wire [7:0] t_r41_c11_8;
  wire [7:0] t_r41_c11_9;
  wire [7:0] t_r41_c11_10;
  wire [7:0] t_r41_c11_11;
  wire [7:0] t_r41_c11_12;
  wire [7:0] t_r41_c12_0;
  wire [7:0] t_r41_c12_1;
  wire [7:0] t_r41_c12_2;
  wire [7:0] t_r41_c12_3;
  wire [7:0] t_r41_c12_4;
  wire [7:0] t_r41_c12_5;
  wire [7:0] t_r41_c12_6;
  wire [7:0] t_r41_c12_7;
  wire [7:0] t_r41_c12_8;
  wire [7:0] t_r41_c12_9;
  wire [7:0] t_r41_c12_10;
  wire [7:0] t_r41_c12_11;
  wire [7:0] t_r41_c12_12;
  wire [7:0] t_r41_c13_0;
  wire [7:0] t_r41_c13_1;
  wire [7:0] t_r41_c13_2;
  wire [7:0] t_r41_c13_3;
  wire [7:0] t_r41_c13_4;
  wire [7:0] t_r41_c13_5;
  wire [7:0] t_r41_c13_6;
  wire [7:0] t_r41_c13_7;
  wire [7:0] t_r41_c13_8;
  wire [7:0] t_r41_c13_9;
  wire [7:0] t_r41_c13_10;
  wire [7:0] t_r41_c13_11;
  wire [7:0] t_r41_c13_12;
  wire [7:0] t_r41_c14_0;
  wire [7:0] t_r41_c14_1;
  wire [7:0] t_r41_c14_2;
  wire [7:0] t_r41_c14_3;
  wire [7:0] t_r41_c14_4;
  wire [7:0] t_r41_c14_5;
  wire [7:0] t_r41_c14_6;
  wire [7:0] t_r41_c14_7;
  wire [7:0] t_r41_c14_8;
  wire [7:0] t_r41_c14_9;
  wire [7:0] t_r41_c14_10;
  wire [7:0] t_r41_c14_11;
  wire [7:0] t_r41_c14_12;
  wire [7:0] t_r41_c15_0;
  wire [7:0] t_r41_c15_1;
  wire [7:0] t_r41_c15_2;
  wire [7:0] t_r41_c15_3;
  wire [7:0] t_r41_c15_4;
  wire [7:0] t_r41_c15_5;
  wire [7:0] t_r41_c15_6;
  wire [7:0] t_r41_c15_7;
  wire [7:0] t_r41_c15_8;
  wire [7:0] t_r41_c15_9;
  wire [7:0] t_r41_c15_10;
  wire [7:0] t_r41_c15_11;
  wire [7:0] t_r41_c15_12;
  wire [7:0] t_r41_c16_0;
  wire [7:0] t_r41_c16_1;
  wire [7:0] t_r41_c16_2;
  wire [7:0] t_r41_c16_3;
  wire [7:0] t_r41_c16_4;
  wire [7:0] t_r41_c16_5;
  wire [7:0] t_r41_c16_6;
  wire [7:0] t_r41_c16_7;
  wire [7:0] t_r41_c16_8;
  wire [7:0] t_r41_c16_9;
  wire [7:0] t_r41_c16_10;
  wire [7:0] t_r41_c16_11;
  wire [7:0] t_r41_c16_12;
  wire [7:0] t_r41_c17_0;
  wire [7:0] t_r41_c17_1;
  wire [7:0] t_r41_c17_2;
  wire [7:0] t_r41_c17_3;
  wire [7:0] t_r41_c17_4;
  wire [7:0] t_r41_c17_5;
  wire [7:0] t_r41_c17_6;
  wire [7:0] t_r41_c17_7;
  wire [7:0] t_r41_c17_8;
  wire [7:0] t_r41_c17_9;
  wire [7:0] t_r41_c17_10;
  wire [7:0] t_r41_c17_11;
  wire [7:0] t_r41_c17_12;
  wire [7:0] t_r41_c18_0;
  wire [7:0] t_r41_c18_1;
  wire [7:0] t_r41_c18_2;
  wire [7:0] t_r41_c18_3;
  wire [7:0] t_r41_c18_4;
  wire [7:0] t_r41_c18_5;
  wire [7:0] t_r41_c18_6;
  wire [7:0] t_r41_c18_7;
  wire [7:0] t_r41_c18_8;
  wire [7:0] t_r41_c18_9;
  wire [7:0] t_r41_c18_10;
  wire [7:0] t_r41_c18_11;
  wire [7:0] t_r41_c18_12;
  wire [7:0] t_r41_c19_0;
  wire [7:0] t_r41_c19_1;
  wire [7:0] t_r41_c19_2;
  wire [7:0] t_r41_c19_3;
  wire [7:0] t_r41_c19_4;
  wire [7:0] t_r41_c19_5;
  wire [7:0] t_r41_c19_6;
  wire [7:0] t_r41_c19_7;
  wire [7:0] t_r41_c19_8;
  wire [7:0] t_r41_c19_9;
  wire [7:0] t_r41_c19_10;
  wire [7:0] t_r41_c19_11;
  wire [7:0] t_r41_c19_12;
  wire [7:0] t_r41_c20_0;
  wire [7:0] t_r41_c20_1;
  wire [7:0] t_r41_c20_2;
  wire [7:0] t_r41_c20_3;
  wire [7:0] t_r41_c20_4;
  wire [7:0] t_r41_c20_5;
  wire [7:0] t_r41_c20_6;
  wire [7:0] t_r41_c20_7;
  wire [7:0] t_r41_c20_8;
  wire [7:0] t_r41_c20_9;
  wire [7:0] t_r41_c20_10;
  wire [7:0] t_r41_c20_11;
  wire [7:0] t_r41_c20_12;
  wire [7:0] t_r41_c21_0;
  wire [7:0] t_r41_c21_1;
  wire [7:0] t_r41_c21_2;
  wire [7:0] t_r41_c21_3;
  wire [7:0] t_r41_c21_4;
  wire [7:0] t_r41_c21_5;
  wire [7:0] t_r41_c21_6;
  wire [7:0] t_r41_c21_7;
  wire [7:0] t_r41_c21_8;
  wire [7:0] t_r41_c21_9;
  wire [7:0] t_r41_c21_10;
  wire [7:0] t_r41_c21_11;
  wire [7:0] t_r41_c21_12;
  wire [7:0] t_r41_c22_0;
  wire [7:0] t_r41_c22_1;
  wire [7:0] t_r41_c22_2;
  wire [7:0] t_r41_c22_3;
  wire [7:0] t_r41_c22_4;
  wire [7:0] t_r41_c22_5;
  wire [7:0] t_r41_c22_6;
  wire [7:0] t_r41_c22_7;
  wire [7:0] t_r41_c22_8;
  wire [7:0] t_r41_c22_9;
  wire [7:0] t_r41_c22_10;
  wire [7:0] t_r41_c22_11;
  wire [7:0] t_r41_c22_12;
  wire [7:0] t_r41_c23_0;
  wire [7:0] t_r41_c23_1;
  wire [7:0] t_r41_c23_2;
  wire [7:0] t_r41_c23_3;
  wire [7:0] t_r41_c23_4;
  wire [7:0] t_r41_c23_5;
  wire [7:0] t_r41_c23_6;
  wire [7:0] t_r41_c23_7;
  wire [7:0] t_r41_c23_8;
  wire [7:0] t_r41_c23_9;
  wire [7:0] t_r41_c23_10;
  wire [7:0] t_r41_c23_11;
  wire [7:0] t_r41_c23_12;
  wire [7:0] t_r41_c24_0;
  wire [7:0] t_r41_c24_1;
  wire [7:0] t_r41_c24_2;
  wire [7:0] t_r41_c24_3;
  wire [7:0] t_r41_c24_4;
  wire [7:0] t_r41_c24_5;
  wire [7:0] t_r41_c24_6;
  wire [7:0] t_r41_c24_7;
  wire [7:0] t_r41_c24_8;
  wire [7:0] t_r41_c24_9;
  wire [7:0] t_r41_c24_10;
  wire [7:0] t_r41_c24_11;
  wire [7:0] t_r41_c24_12;
  wire [7:0] t_r41_c25_0;
  wire [7:0] t_r41_c25_1;
  wire [7:0] t_r41_c25_2;
  wire [7:0] t_r41_c25_3;
  wire [7:0] t_r41_c25_4;
  wire [7:0] t_r41_c25_5;
  wire [7:0] t_r41_c25_6;
  wire [7:0] t_r41_c25_7;
  wire [7:0] t_r41_c25_8;
  wire [7:0] t_r41_c25_9;
  wire [7:0] t_r41_c25_10;
  wire [7:0] t_r41_c25_11;
  wire [7:0] t_r41_c25_12;
  wire [7:0] t_r41_c26_0;
  wire [7:0] t_r41_c26_1;
  wire [7:0] t_r41_c26_2;
  wire [7:0] t_r41_c26_3;
  wire [7:0] t_r41_c26_4;
  wire [7:0] t_r41_c26_5;
  wire [7:0] t_r41_c26_6;
  wire [7:0] t_r41_c26_7;
  wire [7:0] t_r41_c26_8;
  wire [7:0] t_r41_c26_9;
  wire [7:0] t_r41_c26_10;
  wire [7:0] t_r41_c26_11;
  wire [7:0] t_r41_c26_12;
  wire [7:0] t_r41_c27_0;
  wire [7:0] t_r41_c27_1;
  wire [7:0] t_r41_c27_2;
  wire [7:0] t_r41_c27_3;
  wire [7:0] t_r41_c27_4;
  wire [7:0] t_r41_c27_5;
  wire [7:0] t_r41_c27_6;
  wire [7:0] t_r41_c27_7;
  wire [7:0] t_r41_c27_8;
  wire [7:0] t_r41_c27_9;
  wire [7:0] t_r41_c27_10;
  wire [7:0] t_r41_c27_11;
  wire [7:0] t_r41_c27_12;
  wire [7:0] t_r41_c28_0;
  wire [7:0] t_r41_c28_1;
  wire [7:0] t_r41_c28_2;
  wire [7:0] t_r41_c28_3;
  wire [7:0] t_r41_c28_4;
  wire [7:0] t_r41_c28_5;
  wire [7:0] t_r41_c28_6;
  wire [7:0] t_r41_c28_7;
  wire [7:0] t_r41_c28_8;
  wire [7:0] t_r41_c28_9;
  wire [7:0] t_r41_c28_10;
  wire [7:0] t_r41_c28_11;
  wire [7:0] t_r41_c28_12;
  wire [7:0] t_r41_c29_0;
  wire [7:0] t_r41_c29_1;
  wire [7:0] t_r41_c29_2;
  wire [7:0] t_r41_c29_3;
  wire [7:0] t_r41_c29_4;
  wire [7:0] t_r41_c29_5;
  wire [7:0] t_r41_c29_6;
  wire [7:0] t_r41_c29_7;
  wire [7:0] t_r41_c29_8;
  wire [7:0] t_r41_c29_9;
  wire [7:0] t_r41_c29_10;
  wire [7:0] t_r41_c29_11;
  wire [7:0] t_r41_c29_12;
  wire [7:0] t_r41_c30_0;
  wire [7:0] t_r41_c30_1;
  wire [7:0] t_r41_c30_2;
  wire [7:0] t_r41_c30_3;
  wire [7:0] t_r41_c30_4;
  wire [7:0] t_r41_c30_5;
  wire [7:0] t_r41_c30_6;
  wire [7:0] t_r41_c30_7;
  wire [7:0] t_r41_c30_8;
  wire [7:0] t_r41_c30_9;
  wire [7:0] t_r41_c30_10;
  wire [7:0] t_r41_c30_11;
  wire [7:0] t_r41_c30_12;
  wire [7:0] t_r41_c31_0;
  wire [7:0] t_r41_c31_1;
  wire [7:0] t_r41_c31_2;
  wire [7:0] t_r41_c31_3;
  wire [7:0] t_r41_c31_4;
  wire [7:0] t_r41_c31_5;
  wire [7:0] t_r41_c31_6;
  wire [7:0] t_r41_c31_7;
  wire [7:0] t_r41_c31_8;
  wire [7:0] t_r41_c31_9;
  wire [7:0] t_r41_c31_10;
  wire [7:0] t_r41_c31_11;
  wire [7:0] t_r41_c31_12;
  wire [7:0] t_r41_c32_0;
  wire [7:0] t_r41_c32_1;
  wire [7:0] t_r41_c32_2;
  wire [7:0] t_r41_c32_3;
  wire [7:0] t_r41_c32_4;
  wire [7:0] t_r41_c32_5;
  wire [7:0] t_r41_c32_6;
  wire [7:0] t_r41_c32_7;
  wire [7:0] t_r41_c32_8;
  wire [7:0] t_r41_c32_9;
  wire [7:0] t_r41_c32_10;
  wire [7:0] t_r41_c32_11;
  wire [7:0] t_r41_c32_12;
  wire [7:0] t_r41_c33_0;
  wire [7:0] t_r41_c33_1;
  wire [7:0] t_r41_c33_2;
  wire [7:0] t_r41_c33_3;
  wire [7:0] t_r41_c33_4;
  wire [7:0] t_r41_c33_5;
  wire [7:0] t_r41_c33_6;
  wire [7:0] t_r41_c33_7;
  wire [7:0] t_r41_c33_8;
  wire [7:0] t_r41_c33_9;
  wire [7:0] t_r41_c33_10;
  wire [7:0] t_r41_c33_11;
  wire [7:0] t_r41_c33_12;
  wire [7:0] t_r41_c34_0;
  wire [7:0] t_r41_c34_1;
  wire [7:0] t_r41_c34_2;
  wire [7:0] t_r41_c34_3;
  wire [7:0] t_r41_c34_4;
  wire [7:0] t_r41_c34_5;
  wire [7:0] t_r41_c34_6;
  wire [7:0] t_r41_c34_7;
  wire [7:0] t_r41_c34_8;
  wire [7:0] t_r41_c34_9;
  wire [7:0] t_r41_c34_10;
  wire [7:0] t_r41_c34_11;
  wire [7:0] t_r41_c34_12;
  wire [7:0] t_r41_c35_0;
  wire [7:0] t_r41_c35_1;
  wire [7:0] t_r41_c35_2;
  wire [7:0] t_r41_c35_3;
  wire [7:0] t_r41_c35_4;
  wire [7:0] t_r41_c35_5;
  wire [7:0] t_r41_c35_6;
  wire [7:0] t_r41_c35_7;
  wire [7:0] t_r41_c35_8;
  wire [7:0] t_r41_c35_9;
  wire [7:0] t_r41_c35_10;
  wire [7:0] t_r41_c35_11;
  wire [7:0] t_r41_c35_12;
  wire [7:0] t_r41_c36_0;
  wire [7:0] t_r41_c36_1;
  wire [7:0] t_r41_c36_2;
  wire [7:0] t_r41_c36_3;
  wire [7:0] t_r41_c36_4;
  wire [7:0] t_r41_c36_5;
  wire [7:0] t_r41_c36_6;
  wire [7:0] t_r41_c36_7;
  wire [7:0] t_r41_c36_8;
  wire [7:0] t_r41_c36_9;
  wire [7:0] t_r41_c36_10;
  wire [7:0] t_r41_c36_11;
  wire [7:0] t_r41_c36_12;
  wire [7:0] t_r41_c37_0;
  wire [7:0] t_r41_c37_1;
  wire [7:0] t_r41_c37_2;
  wire [7:0] t_r41_c37_3;
  wire [7:0] t_r41_c37_4;
  wire [7:0] t_r41_c37_5;
  wire [7:0] t_r41_c37_6;
  wire [7:0] t_r41_c37_7;
  wire [7:0] t_r41_c37_8;
  wire [7:0] t_r41_c37_9;
  wire [7:0] t_r41_c37_10;
  wire [7:0] t_r41_c37_11;
  wire [7:0] t_r41_c37_12;
  wire [7:0] t_r41_c38_0;
  wire [7:0] t_r41_c38_1;
  wire [7:0] t_r41_c38_2;
  wire [7:0] t_r41_c38_3;
  wire [7:0] t_r41_c38_4;
  wire [7:0] t_r41_c38_5;
  wire [7:0] t_r41_c38_6;
  wire [7:0] t_r41_c38_7;
  wire [7:0] t_r41_c38_8;
  wire [7:0] t_r41_c38_9;
  wire [7:0] t_r41_c38_10;
  wire [7:0] t_r41_c38_11;
  wire [7:0] t_r41_c38_12;
  wire [7:0] t_r41_c39_0;
  wire [7:0] t_r41_c39_1;
  wire [7:0] t_r41_c39_2;
  wire [7:0] t_r41_c39_3;
  wire [7:0] t_r41_c39_4;
  wire [7:0] t_r41_c39_5;
  wire [7:0] t_r41_c39_6;
  wire [7:0] t_r41_c39_7;
  wire [7:0] t_r41_c39_8;
  wire [7:0] t_r41_c39_9;
  wire [7:0] t_r41_c39_10;
  wire [7:0] t_r41_c39_11;
  wire [7:0] t_r41_c39_12;
  wire [7:0] t_r41_c40_0;
  wire [7:0] t_r41_c40_1;
  wire [7:0] t_r41_c40_2;
  wire [7:0] t_r41_c40_3;
  wire [7:0] t_r41_c40_4;
  wire [7:0] t_r41_c40_5;
  wire [7:0] t_r41_c40_6;
  wire [7:0] t_r41_c40_7;
  wire [7:0] t_r41_c40_8;
  wire [7:0] t_r41_c40_9;
  wire [7:0] t_r41_c40_10;
  wire [7:0] t_r41_c40_11;
  wire [7:0] t_r41_c40_12;
  wire [7:0] t_r41_c41_0;
  wire [7:0] t_r41_c41_1;
  wire [7:0] t_r41_c41_2;
  wire [7:0] t_r41_c41_3;
  wire [7:0] t_r41_c41_4;
  wire [7:0] t_r41_c41_5;
  wire [7:0] t_r41_c41_6;
  wire [7:0] t_r41_c41_7;
  wire [7:0] t_r41_c41_8;
  wire [7:0] t_r41_c41_9;
  wire [7:0] t_r41_c41_10;
  wire [7:0] t_r41_c41_11;
  wire [7:0] t_r41_c41_12;
  wire [7:0] t_r41_c42_0;
  wire [7:0] t_r41_c42_1;
  wire [7:0] t_r41_c42_2;
  wire [7:0] t_r41_c42_3;
  wire [7:0] t_r41_c42_4;
  wire [7:0] t_r41_c42_5;
  wire [7:0] t_r41_c42_6;
  wire [7:0] t_r41_c42_7;
  wire [7:0] t_r41_c42_8;
  wire [7:0] t_r41_c42_9;
  wire [7:0] t_r41_c42_10;
  wire [7:0] t_r41_c42_11;
  wire [7:0] t_r41_c42_12;
  wire [7:0] t_r41_c43_0;
  wire [7:0] t_r41_c43_1;
  wire [7:0] t_r41_c43_2;
  wire [7:0] t_r41_c43_3;
  wire [7:0] t_r41_c43_4;
  wire [7:0] t_r41_c43_5;
  wire [7:0] t_r41_c43_6;
  wire [7:0] t_r41_c43_7;
  wire [7:0] t_r41_c43_8;
  wire [7:0] t_r41_c43_9;
  wire [7:0] t_r41_c43_10;
  wire [7:0] t_r41_c43_11;
  wire [7:0] t_r41_c43_12;
  wire [7:0] t_r41_c44_0;
  wire [7:0] t_r41_c44_1;
  wire [7:0] t_r41_c44_2;
  wire [7:0] t_r41_c44_3;
  wire [7:0] t_r41_c44_4;
  wire [7:0] t_r41_c44_5;
  wire [7:0] t_r41_c44_6;
  wire [7:0] t_r41_c44_7;
  wire [7:0] t_r41_c44_8;
  wire [7:0] t_r41_c44_9;
  wire [7:0] t_r41_c44_10;
  wire [7:0] t_r41_c44_11;
  wire [7:0] t_r41_c44_12;
  wire [7:0] t_r41_c45_0;
  wire [7:0] t_r41_c45_1;
  wire [7:0] t_r41_c45_2;
  wire [7:0] t_r41_c45_3;
  wire [7:0] t_r41_c45_4;
  wire [7:0] t_r41_c45_5;
  wire [7:0] t_r41_c45_6;
  wire [7:0] t_r41_c45_7;
  wire [7:0] t_r41_c45_8;
  wire [7:0] t_r41_c45_9;
  wire [7:0] t_r41_c45_10;
  wire [7:0] t_r41_c45_11;
  wire [7:0] t_r41_c45_12;
  wire [7:0] t_r41_c46_0;
  wire [7:0] t_r41_c46_1;
  wire [7:0] t_r41_c46_2;
  wire [7:0] t_r41_c46_3;
  wire [7:0] t_r41_c46_4;
  wire [7:0] t_r41_c46_5;
  wire [7:0] t_r41_c46_6;
  wire [7:0] t_r41_c46_7;
  wire [7:0] t_r41_c46_8;
  wire [7:0] t_r41_c46_9;
  wire [7:0] t_r41_c46_10;
  wire [7:0] t_r41_c46_11;
  wire [7:0] t_r41_c46_12;
  wire [7:0] t_r41_c47_0;
  wire [7:0] t_r41_c47_1;
  wire [7:0] t_r41_c47_2;
  wire [7:0] t_r41_c47_3;
  wire [7:0] t_r41_c47_4;
  wire [7:0] t_r41_c47_5;
  wire [7:0] t_r41_c47_6;
  wire [7:0] t_r41_c47_7;
  wire [7:0] t_r41_c47_8;
  wire [7:0] t_r41_c47_9;
  wire [7:0] t_r41_c47_10;
  wire [7:0] t_r41_c47_11;
  wire [7:0] t_r41_c47_12;
  wire [7:0] t_r41_c48_0;
  wire [7:0] t_r41_c48_1;
  wire [7:0] t_r41_c48_2;
  wire [7:0] t_r41_c48_3;
  wire [7:0] t_r41_c48_4;
  wire [7:0] t_r41_c48_5;
  wire [7:0] t_r41_c48_6;
  wire [7:0] t_r41_c48_7;
  wire [7:0] t_r41_c48_8;
  wire [7:0] t_r41_c48_9;
  wire [7:0] t_r41_c48_10;
  wire [7:0] t_r41_c48_11;
  wire [7:0] t_r41_c48_12;
  wire [7:0] t_r41_c49_0;
  wire [7:0] t_r41_c49_1;
  wire [7:0] t_r41_c49_2;
  wire [7:0] t_r41_c49_3;
  wire [7:0] t_r41_c49_4;
  wire [7:0] t_r41_c49_5;
  wire [7:0] t_r41_c49_6;
  wire [7:0] t_r41_c49_7;
  wire [7:0] t_r41_c49_8;
  wire [7:0] t_r41_c49_9;
  wire [7:0] t_r41_c49_10;
  wire [7:0] t_r41_c49_11;
  wire [7:0] t_r41_c49_12;
  wire [7:0] t_r41_c50_0;
  wire [7:0] t_r41_c50_1;
  wire [7:0] t_r41_c50_2;
  wire [7:0] t_r41_c50_3;
  wire [7:0] t_r41_c50_4;
  wire [7:0] t_r41_c50_5;
  wire [7:0] t_r41_c50_6;
  wire [7:0] t_r41_c50_7;
  wire [7:0] t_r41_c50_8;
  wire [7:0] t_r41_c50_9;
  wire [7:0] t_r41_c50_10;
  wire [7:0] t_r41_c50_11;
  wire [7:0] t_r41_c50_12;
  wire [7:0] t_r41_c51_0;
  wire [7:0] t_r41_c51_1;
  wire [7:0] t_r41_c51_2;
  wire [7:0] t_r41_c51_3;
  wire [7:0] t_r41_c51_4;
  wire [7:0] t_r41_c51_5;
  wire [7:0] t_r41_c51_6;
  wire [7:0] t_r41_c51_7;
  wire [7:0] t_r41_c51_8;
  wire [7:0] t_r41_c51_9;
  wire [7:0] t_r41_c51_10;
  wire [7:0] t_r41_c51_11;
  wire [7:0] t_r41_c51_12;
  wire [7:0] t_r41_c52_0;
  wire [7:0] t_r41_c52_1;
  wire [7:0] t_r41_c52_2;
  wire [7:0] t_r41_c52_3;
  wire [7:0] t_r41_c52_4;
  wire [7:0] t_r41_c52_5;
  wire [7:0] t_r41_c52_6;
  wire [7:0] t_r41_c52_7;
  wire [7:0] t_r41_c52_8;
  wire [7:0] t_r41_c52_9;
  wire [7:0] t_r41_c52_10;
  wire [7:0] t_r41_c52_11;
  wire [7:0] t_r41_c52_12;
  wire [7:0] t_r41_c53_0;
  wire [7:0] t_r41_c53_1;
  wire [7:0] t_r41_c53_2;
  wire [7:0] t_r41_c53_3;
  wire [7:0] t_r41_c53_4;
  wire [7:0] t_r41_c53_5;
  wire [7:0] t_r41_c53_6;
  wire [7:0] t_r41_c53_7;
  wire [7:0] t_r41_c53_8;
  wire [7:0] t_r41_c53_9;
  wire [7:0] t_r41_c53_10;
  wire [7:0] t_r41_c53_11;
  wire [7:0] t_r41_c53_12;
  wire [7:0] t_r41_c54_0;
  wire [7:0] t_r41_c54_1;
  wire [7:0] t_r41_c54_2;
  wire [7:0] t_r41_c54_3;
  wire [7:0] t_r41_c54_4;
  wire [7:0] t_r41_c54_5;
  wire [7:0] t_r41_c54_6;
  wire [7:0] t_r41_c54_7;
  wire [7:0] t_r41_c54_8;
  wire [7:0] t_r41_c54_9;
  wire [7:0] t_r41_c54_10;
  wire [7:0] t_r41_c54_11;
  wire [7:0] t_r41_c54_12;
  wire [7:0] t_r41_c55_0;
  wire [7:0] t_r41_c55_1;
  wire [7:0] t_r41_c55_2;
  wire [7:0] t_r41_c55_3;
  wire [7:0] t_r41_c55_4;
  wire [7:0] t_r41_c55_5;
  wire [7:0] t_r41_c55_6;
  wire [7:0] t_r41_c55_7;
  wire [7:0] t_r41_c55_8;
  wire [7:0] t_r41_c55_9;
  wire [7:0] t_r41_c55_10;
  wire [7:0] t_r41_c55_11;
  wire [7:0] t_r41_c55_12;
  wire [7:0] t_r41_c56_0;
  wire [7:0] t_r41_c56_1;
  wire [7:0] t_r41_c56_2;
  wire [7:0] t_r41_c56_3;
  wire [7:0] t_r41_c56_4;
  wire [7:0] t_r41_c56_5;
  wire [7:0] t_r41_c56_6;
  wire [7:0] t_r41_c56_7;
  wire [7:0] t_r41_c56_8;
  wire [7:0] t_r41_c56_9;
  wire [7:0] t_r41_c56_10;
  wire [7:0] t_r41_c56_11;
  wire [7:0] t_r41_c56_12;
  wire [7:0] t_r41_c57_0;
  wire [7:0] t_r41_c57_1;
  wire [7:0] t_r41_c57_2;
  wire [7:0] t_r41_c57_3;
  wire [7:0] t_r41_c57_4;
  wire [7:0] t_r41_c57_5;
  wire [7:0] t_r41_c57_6;
  wire [7:0] t_r41_c57_7;
  wire [7:0] t_r41_c57_8;
  wire [7:0] t_r41_c57_9;
  wire [7:0] t_r41_c57_10;
  wire [7:0] t_r41_c57_11;
  wire [7:0] t_r41_c57_12;
  wire [7:0] t_r41_c58_0;
  wire [7:0] t_r41_c58_1;
  wire [7:0] t_r41_c58_2;
  wire [7:0] t_r41_c58_3;
  wire [7:0] t_r41_c58_4;
  wire [7:0] t_r41_c58_5;
  wire [7:0] t_r41_c58_6;
  wire [7:0] t_r41_c58_7;
  wire [7:0] t_r41_c58_8;
  wire [7:0] t_r41_c58_9;
  wire [7:0] t_r41_c58_10;
  wire [7:0] t_r41_c58_11;
  wire [7:0] t_r41_c58_12;
  wire [7:0] t_r41_c59_0;
  wire [7:0] t_r41_c59_1;
  wire [7:0] t_r41_c59_2;
  wire [7:0] t_r41_c59_3;
  wire [7:0] t_r41_c59_4;
  wire [7:0] t_r41_c59_5;
  wire [7:0] t_r41_c59_6;
  wire [7:0] t_r41_c59_7;
  wire [7:0] t_r41_c59_8;
  wire [7:0] t_r41_c59_9;
  wire [7:0] t_r41_c59_10;
  wire [7:0] t_r41_c59_11;
  wire [7:0] t_r41_c59_12;
  wire [7:0] t_r41_c60_0;
  wire [7:0] t_r41_c60_1;
  wire [7:0] t_r41_c60_2;
  wire [7:0] t_r41_c60_3;
  wire [7:0] t_r41_c60_4;
  wire [7:0] t_r41_c60_5;
  wire [7:0] t_r41_c60_6;
  wire [7:0] t_r41_c60_7;
  wire [7:0] t_r41_c60_8;
  wire [7:0] t_r41_c60_9;
  wire [7:0] t_r41_c60_10;
  wire [7:0] t_r41_c60_11;
  wire [7:0] t_r41_c60_12;
  wire [7:0] t_r41_c61_0;
  wire [7:0] t_r41_c61_1;
  wire [7:0] t_r41_c61_2;
  wire [7:0] t_r41_c61_3;
  wire [7:0] t_r41_c61_4;
  wire [7:0] t_r41_c61_5;
  wire [7:0] t_r41_c61_6;
  wire [7:0] t_r41_c61_7;
  wire [7:0] t_r41_c61_8;
  wire [7:0] t_r41_c61_9;
  wire [7:0] t_r41_c61_10;
  wire [7:0] t_r41_c61_11;
  wire [7:0] t_r41_c61_12;
  wire [7:0] t_r41_c62_0;
  wire [7:0] t_r41_c62_1;
  wire [7:0] t_r41_c62_2;
  wire [7:0] t_r41_c62_3;
  wire [7:0] t_r41_c62_4;
  wire [7:0] t_r41_c62_5;
  wire [7:0] t_r41_c62_6;
  wire [7:0] t_r41_c62_7;
  wire [7:0] t_r41_c62_8;
  wire [7:0] t_r41_c62_9;
  wire [7:0] t_r41_c62_10;
  wire [7:0] t_r41_c62_11;
  wire [7:0] t_r41_c62_12;
  wire [7:0] t_r41_c63_0;
  wire [7:0] t_r41_c63_1;
  wire [7:0] t_r41_c63_2;
  wire [7:0] t_r41_c63_3;
  wire [7:0] t_r41_c63_4;
  wire [7:0] t_r41_c63_5;
  wire [7:0] t_r41_c63_6;
  wire [7:0] t_r41_c63_7;
  wire [7:0] t_r41_c63_8;
  wire [7:0] t_r41_c63_9;
  wire [7:0] t_r41_c63_10;
  wire [7:0] t_r41_c63_11;
  wire [7:0] t_r41_c63_12;
  wire [7:0] t_r41_c64_0;
  wire [7:0] t_r41_c64_1;
  wire [7:0] t_r41_c64_2;
  wire [7:0] t_r41_c64_3;
  wire [7:0] t_r41_c64_4;
  wire [7:0] t_r41_c64_5;
  wire [7:0] t_r41_c64_6;
  wire [7:0] t_r41_c64_7;
  wire [7:0] t_r41_c64_8;
  wire [7:0] t_r41_c64_9;
  wire [7:0] t_r41_c64_10;
  wire [7:0] t_r41_c64_11;
  wire [7:0] t_r41_c64_12;
  wire [7:0] t_r41_c65_0;
  wire [7:0] t_r41_c65_1;
  wire [7:0] t_r41_c65_2;
  wire [7:0] t_r41_c65_3;
  wire [7:0] t_r41_c65_4;
  wire [7:0] t_r41_c65_5;
  wire [7:0] t_r41_c65_6;
  wire [7:0] t_r41_c65_7;
  wire [7:0] t_r41_c65_8;
  wire [7:0] t_r41_c65_9;
  wire [7:0] t_r41_c65_10;
  wire [7:0] t_r41_c65_11;
  wire [7:0] t_r41_c65_12;
  wire [7:0] t_r42_c0_0;
  wire [7:0] t_r42_c0_1;
  wire [7:0] t_r42_c0_2;
  wire [7:0] t_r42_c0_3;
  wire [7:0] t_r42_c0_4;
  wire [7:0] t_r42_c0_5;
  wire [7:0] t_r42_c0_6;
  wire [7:0] t_r42_c0_7;
  wire [7:0] t_r42_c0_8;
  wire [7:0] t_r42_c0_9;
  wire [7:0] t_r42_c0_10;
  wire [7:0] t_r42_c0_11;
  wire [7:0] t_r42_c0_12;
  wire [7:0] t_r42_c1_0;
  wire [7:0] t_r42_c1_1;
  wire [7:0] t_r42_c1_2;
  wire [7:0] t_r42_c1_3;
  wire [7:0] t_r42_c1_4;
  wire [7:0] t_r42_c1_5;
  wire [7:0] t_r42_c1_6;
  wire [7:0] t_r42_c1_7;
  wire [7:0] t_r42_c1_8;
  wire [7:0] t_r42_c1_9;
  wire [7:0] t_r42_c1_10;
  wire [7:0] t_r42_c1_11;
  wire [7:0] t_r42_c1_12;
  wire [7:0] t_r42_c2_0;
  wire [7:0] t_r42_c2_1;
  wire [7:0] t_r42_c2_2;
  wire [7:0] t_r42_c2_3;
  wire [7:0] t_r42_c2_4;
  wire [7:0] t_r42_c2_5;
  wire [7:0] t_r42_c2_6;
  wire [7:0] t_r42_c2_7;
  wire [7:0] t_r42_c2_8;
  wire [7:0] t_r42_c2_9;
  wire [7:0] t_r42_c2_10;
  wire [7:0] t_r42_c2_11;
  wire [7:0] t_r42_c2_12;
  wire [7:0] t_r42_c3_0;
  wire [7:0] t_r42_c3_1;
  wire [7:0] t_r42_c3_2;
  wire [7:0] t_r42_c3_3;
  wire [7:0] t_r42_c3_4;
  wire [7:0] t_r42_c3_5;
  wire [7:0] t_r42_c3_6;
  wire [7:0] t_r42_c3_7;
  wire [7:0] t_r42_c3_8;
  wire [7:0] t_r42_c3_9;
  wire [7:0] t_r42_c3_10;
  wire [7:0] t_r42_c3_11;
  wire [7:0] t_r42_c3_12;
  wire [7:0] t_r42_c4_0;
  wire [7:0] t_r42_c4_1;
  wire [7:0] t_r42_c4_2;
  wire [7:0] t_r42_c4_3;
  wire [7:0] t_r42_c4_4;
  wire [7:0] t_r42_c4_5;
  wire [7:0] t_r42_c4_6;
  wire [7:0] t_r42_c4_7;
  wire [7:0] t_r42_c4_8;
  wire [7:0] t_r42_c4_9;
  wire [7:0] t_r42_c4_10;
  wire [7:0] t_r42_c4_11;
  wire [7:0] t_r42_c4_12;
  wire [7:0] t_r42_c5_0;
  wire [7:0] t_r42_c5_1;
  wire [7:0] t_r42_c5_2;
  wire [7:0] t_r42_c5_3;
  wire [7:0] t_r42_c5_4;
  wire [7:0] t_r42_c5_5;
  wire [7:0] t_r42_c5_6;
  wire [7:0] t_r42_c5_7;
  wire [7:0] t_r42_c5_8;
  wire [7:0] t_r42_c5_9;
  wire [7:0] t_r42_c5_10;
  wire [7:0] t_r42_c5_11;
  wire [7:0] t_r42_c5_12;
  wire [7:0] t_r42_c6_0;
  wire [7:0] t_r42_c6_1;
  wire [7:0] t_r42_c6_2;
  wire [7:0] t_r42_c6_3;
  wire [7:0] t_r42_c6_4;
  wire [7:0] t_r42_c6_5;
  wire [7:0] t_r42_c6_6;
  wire [7:0] t_r42_c6_7;
  wire [7:0] t_r42_c6_8;
  wire [7:0] t_r42_c6_9;
  wire [7:0] t_r42_c6_10;
  wire [7:0] t_r42_c6_11;
  wire [7:0] t_r42_c6_12;
  wire [7:0] t_r42_c7_0;
  wire [7:0] t_r42_c7_1;
  wire [7:0] t_r42_c7_2;
  wire [7:0] t_r42_c7_3;
  wire [7:0] t_r42_c7_4;
  wire [7:0] t_r42_c7_5;
  wire [7:0] t_r42_c7_6;
  wire [7:0] t_r42_c7_7;
  wire [7:0] t_r42_c7_8;
  wire [7:0] t_r42_c7_9;
  wire [7:0] t_r42_c7_10;
  wire [7:0] t_r42_c7_11;
  wire [7:0] t_r42_c7_12;
  wire [7:0] t_r42_c8_0;
  wire [7:0] t_r42_c8_1;
  wire [7:0] t_r42_c8_2;
  wire [7:0] t_r42_c8_3;
  wire [7:0] t_r42_c8_4;
  wire [7:0] t_r42_c8_5;
  wire [7:0] t_r42_c8_6;
  wire [7:0] t_r42_c8_7;
  wire [7:0] t_r42_c8_8;
  wire [7:0] t_r42_c8_9;
  wire [7:0] t_r42_c8_10;
  wire [7:0] t_r42_c8_11;
  wire [7:0] t_r42_c8_12;
  wire [7:0] t_r42_c9_0;
  wire [7:0] t_r42_c9_1;
  wire [7:0] t_r42_c9_2;
  wire [7:0] t_r42_c9_3;
  wire [7:0] t_r42_c9_4;
  wire [7:0] t_r42_c9_5;
  wire [7:0] t_r42_c9_6;
  wire [7:0] t_r42_c9_7;
  wire [7:0] t_r42_c9_8;
  wire [7:0] t_r42_c9_9;
  wire [7:0] t_r42_c9_10;
  wire [7:0] t_r42_c9_11;
  wire [7:0] t_r42_c9_12;
  wire [7:0] t_r42_c10_0;
  wire [7:0] t_r42_c10_1;
  wire [7:0] t_r42_c10_2;
  wire [7:0] t_r42_c10_3;
  wire [7:0] t_r42_c10_4;
  wire [7:0] t_r42_c10_5;
  wire [7:0] t_r42_c10_6;
  wire [7:0] t_r42_c10_7;
  wire [7:0] t_r42_c10_8;
  wire [7:0] t_r42_c10_9;
  wire [7:0] t_r42_c10_10;
  wire [7:0] t_r42_c10_11;
  wire [7:0] t_r42_c10_12;
  wire [7:0] t_r42_c11_0;
  wire [7:0] t_r42_c11_1;
  wire [7:0] t_r42_c11_2;
  wire [7:0] t_r42_c11_3;
  wire [7:0] t_r42_c11_4;
  wire [7:0] t_r42_c11_5;
  wire [7:0] t_r42_c11_6;
  wire [7:0] t_r42_c11_7;
  wire [7:0] t_r42_c11_8;
  wire [7:0] t_r42_c11_9;
  wire [7:0] t_r42_c11_10;
  wire [7:0] t_r42_c11_11;
  wire [7:0] t_r42_c11_12;
  wire [7:0] t_r42_c12_0;
  wire [7:0] t_r42_c12_1;
  wire [7:0] t_r42_c12_2;
  wire [7:0] t_r42_c12_3;
  wire [7:0] t_r42_c12_4;
  wire [7:0] t_r42_c12_5;
  wire [7:0] t_r42_c12_6;
  wire [7:0] t_r42_c12_7;
  wire [7:0] t_r42_c12_8;
  wire [7:0] t_r42_c12_9;
  wire [7:0] t_r42_c12_10;
  wire [7:0] t_r42_c12_11;
  wire [7:0] t_r42_c12_12;
  wire [7:0] t_r42_c13_0;
  wire [7:0] t_r42_c13_1;
  wire [7:0] t_r42_c13_2;
  wire [7:0] t_r42_c13_3;
  wire [7:0] t_r42_c13_4;
  wire [7:0] t_r42_c13_5;
  wire [7:0] t_r42_c13_6;
  wire [7:0] t_r42_c13_7;
  wire [7:0] t_r42_c13_8;
  wire [7:0] t_r42_c13_9;
  wire [7:0] t_r42_c13_10;
  wire [7:0] t_r42_c13_11;
  wire [7:0] t_r42_c13_12;
  wire [7:0] t_r42_c14_0;
  wire [7:0] t_r42_c14_1;
  wire [7:0] t_r42_c14_2;
  wire [7:0] t_r42_c14_3;
  wire [7:0] t_r42_c14_4;
  wire [7:0] t_r42_c14_5;
  wire [7:0] t_r42_c14_6;
  wire [7:0] t_r42_c14_7;
  wire [7:0] t_r42_c14_8;
  wire [7:0] t_r42_c14_9;
  wire [7:0] t_r42_c14_10;
  wire [7:0] t_r42_c14_11;
  wire [7:0] t_r42_c14_12;
  wire [7:0] t_r42_c15_0;
  wire [7:0] t_r42_c15_1;
  wire [7:0] t_r42_c15_2;
  wire [7:0] t_r42_c15_3;
  wire [7:0] t_r42_c15_4;
  wire [7:0] t_r42_c15_5;
  wire [7:0] t_r42_c15_6;
  wire [7:0] t_r42_c15_7;
  wire [7:0] t_r42_c15_8;
  wire [7:0] t_r42_c15_9;
  wire [7:0] t_r42_c15_10;
  wire [7:0] t_r42_c15_11;
  wire [7:0] t_r42_c15_12;
  wire [7:0] t_r42_c16_0;
  wire [7:0] t_r42_c16_1;
  wire [7:0] t_r42_c16_2;
  wire [7:0] t_r42_c16_3;
  wire [7:0] t_r42_c16_4;
  wire [7:0] t_r42_c16_5;
  wire [7:0] t_r42_c16_6;
  wire [7:0] t_r42_c16_7;
  wire [7:0] t_r42_c16_8;
  wire [7:0] t_r42_c16_9;
  wire [7:0] t_r42_c16_10;
  wire [7:0] t_r42_c16_11;
  wire [7:0] t_r42_c16_12;
  wire [7:0] t_r42_c17_0;
  wire [7:0] t_r42_c17_1;
  wire [7:0] t_r42_c17_2;
  wire [7:0] t_r42_c17_3;
  wire [7:0] t_r42_c17_4;
  wire [7:0] t_r42_c17_5;
  wire [7:0] t_r42_c17_6;
  wire [7:0] t_r42_c17_7;
  wire [7:0] t_r42_c17_8;
  wire [7:0] t_r42_c17_9;
  wire [7:0] t_r42_c17_10;
  wire [7:0] t_r42_c17_11;
  wire [7:0] t_r42_c17_12;
  wire [7:0] t_r42_c18_0;
  wire [7:0] t_r42_c18_1;
  wire [7:0] t_r42_c18_2;
  wire [7:0] t_r42_c18_3;
  wire [7:0] t_r42_c18_4;
  wire [7:0] t_r42_c18_5;
  wire [7:0] t_r42_c18_6;
  wire [7:0] t_r42_c18_7;
  wire [7:0] t_r42_c18_8;
  wire [7:0] t_r42_c18_9;
  wire [7:0] t_r42_c18_10;
  wire [7:0] t_r42_c18_11;
  wire [7:0] t_r42_c18_12;
  wire [7:0] t_r42_c19_0;
  wire [7:0] t_r42_c19_1;
  wire [7:0] t_r42_c19_2;
  wire [7:0] t_r42_c19_3;
  wire [7:0] t_r42_c19_4;
  wire [7:0] t_r42_c19_5;
  wire [7:0] t_r42_c19_6;
  wire [7:0] t_r42_c19_7;
  wire [7:0] t_r42_c19_8;
  wire [7:0] t_r42_c19_9;
  wire [7:0] t_r42_c19_10;
  wire [7:0] t_r42_c19_11;
  wire [7:0] t_r42_c19_12;
  wire [7:0] t_r42_c20_0;
  wire [7:0] t_r42_c20_1;
  wire [7:0] t_r42_c20_2;
  wire [7:0] t_r42_c20_3;
  wire [7:0] t_r42_c20_4;
  wire [7:0] t_r42_c20_5;
  wire [7:0] t_r42_c20_6;
  wire [7:0] t_r42_c20_7;
  wire [7:0] t_r42_c20_8;
  wire [7:0] t_r42_c20_9;
  wire [7:0] t_r42_c20_10;
  wire [7:0] t_r42_c20_11;
  wire [7:0] t_r42_c20_12;
  wire [7:0] t_r42_c21_0;
  wire [7:0] t_r42_c21_1;
  wire [7:0] t_r42_c21_2;
  wire [7:0] t_r42_c21_3;
  wire [7:0] t_r42_c21_4;
  wire [7:0] t_r42_c21_5;
  wire [7:0] t_r42_c21_6;
  wire [7:0] t_r42_c21_7;
  wire [7:0] t_r42_c21_8;
  wire [7:0] t_r42_c21_9;
  wire [7:0] t_r42_c21_10;
  wire [7:0] t_r42_c21_11;
  wire [7:0] t_r42_c21_12;
  wire [7:0] t_r42_c22_0;
  wire [7:0] t_r42_c22_1;
  wire [7:0] t_r42_c22_2;
  wire [7:0] t_r42_c22_3;
  wire [7:0] t_r42_c22_4;
  wire [7:0] t_r42_c22_5;
  wire [7:0] t_r42_c22_6;
  wire [7:0] t_r42_c22_7;
  wire [7:0] t_r42_c22_8;
  wire [7:0] t_r42_c22_9;
  wire [7:0] t_r42_c22_10;
  wire [7:0] t_r42_c22_11;
  wire [7:0] t_r42_c22_12;
  wire [7:0] t_r42_c23_0;
  wire [7:0] t_r42_c23_1;
  wire [7:0] t_r42_c23_2;
  wire [7:0] t_r42_c23_3;
  wire [7:0] t_r42_c23_4;
  wire [7:0] t_r42_c23_5;
  wire [7:0] t_r42_c23_6;
  wire [7:0] t_r42_c23_7;
  wire [7:0] t_r42_c23_8;
  wire [7:0] t_r42_c23_9;
  wire [7:0] t_r42_c23_10;
  wire [7:0] t_r42_c23_11;
  wire [7:0] t_r42_c23_12;
  wire [7:0] t_r42_c24_0;
  wire [7:0] t_r42_c24_1;
  wire [7:0] t_r42_c24_2;
  wire [7:0] t_r42_c24_3;
  wire [7:0] t_r42_c24_4;
  wire [7:0] t_r42_c24_5;
  wire [7:0] t_r42_c24_6;
  wire [7:0] t_r42_c24_7;
  wire [7:0] t_r42_c24_8;
  wire [7:0] t_r42_c24_9;
  wire [7:0] t_r42_c24_10;
  wire [7:0] t_r42_c24_11;
  wire [7:0] t_r42_c24_12;
  wire [7:0] t_r42_c25_0;
  wire [7:0] t_r42_c25_1;
  wire [7:0] t_r42_c25_2;
  wire [7:0] t_r42_c25_3;
  wire [7:0] t_r42_c25_4;
  wire [7:0] t_r42_c25_5;
  wire [7:0] t_r42_c25_6;
  wire [7:0] t_r42_c25_7;
  wire [7:0] t_r42_c25_8;
  wire [7:0] t_r42_c25_9;
  wire [7:0] t_r42_c25_10;
  wire [7:0] t_r42_c25_11;
  wire [7:0] t_r42_c25_12;
  wire [7:0] t_r42_c26_0;
  wire [7:0] t_r42_c26_1;
  wire [7:0] t_r42_c26_2;
  wire [7:0] t_r42_c26_3;
  wire [7:0] t_r42_c26_4;
  wire [7:0] t_r42_c26_5;
  wire [7:0] t_r42_c26_6;
  wire [7:0] t_r42_c26_7;
  wire [7:0] t_r42_c26_8;
  wire [7:0] t_r42_c26_9;
  wire [7:0] t_r42_c26_10;
  wire [7:0] t_r42_c26_11;
  wire [7:0] t_r42_c26_12;
  wire [7:0] t_r42_c27_0;
  wire [7:0] t_r42_c27_1;
  wire [7:0] t_r42_c27_2;
  wire [7:0] t_r42_c27_3;
  wire [7:0] t_r42_c27_4;
  wire [7:0] t_r42_c27_5;
  wire [7:0] t_r42_c27_6;
  wire [7:0] t_r42_c27_7;
  wire [7:0] t_r42_c27_8;
  wire [7:0] t_r42_c27_9;
  wire [7:0] t_r42_c27_10;
  wire [7:0] t_r42_c27_11;
  wire [7:0] t_r42_c27_12;
  wire [7:0] t_r42_c28_0;
  wire [7:0] t_r42_c28_1;
  wire [7:0] t_r42_c28_2;
  wire [7:0] t_r42_c28_3;
  wire [7:0] t_r42_c28_4;
  wire [7:0] t_r42_c28_5;
  wire [7:0] t_r42_c28_6;
  wire [7:0] t_r42_c28_7;
  wire [7:0] t_r42_c28_8;
  wire [7:0] t_r42_c28_9;
  wire [7:0] t_r42_c28_10;
  wire [7:0] t_r42_c28_11;
  wire [7:0] t_r42_c28_12;
  wire [7:0] t_r42_c29_0;
  wire [7:0] t_r42_c29_1;
  wire [7:0] t_r42_c29_2;
  wire [7:0] t_r42_c29_3;
  wire [7:0] t_r42_c29_4;
  wire [7:0] t_r42_c29_5;
  wire [7:0] t_r42_c29_6;
  wire [7:0] t_r42_c29_7;
  wire [7:0] t_r42_c29_8;
  wire [7:0] t_r42_c29_9;
  wire [7:0] t_r42_c29_10;
  wire [7:0] t_r42_c29_11;
  wire [7:0] t_r42_c29_12;
  wire [7:0] t_r42_c30_0;
  wire [7:0] t_r42_c30_1;
  wire [7:0] t_r42_c30_2;
  wire [7:0] t_r42_c30_3;
  wire [7:0] t_r42_c30_4;
  wire [7:0] t_r42_c30_5;
  wire [7:0] t_r42_c30_6;
  wire [7:0] t_r42_c30_7;
  wire [7:0] t_r42_c30_8;
  wire [7:0] t_r42_c30_9;
  wire [7:0] t_r42_c30_10;
  wire [7:0] t_r42_c30_11;
  wire [7:0] t_r42_c30_12;
  wire [7:0] t_r42_c31_0;
  wire [7:0] t_r42_c31_1;
  wire [7:0] t_r42_c31_2;
  wire [7:0] t_r42_c31_3;
  wire [7:0] t_r42_c31_4;
  wire [7:0] t_r42_c31_5;
  wire [7:0] t_r42_c31_6;
  wire [7:0] t_r42_c31_7;
  wire [7:0] t_r42_c31_8;
  wire [7:0] t_r42_c31_9;
  wire [7:0] t_r42_c31_10;
  wire [7:0] t_r42_c31_11;
  wire [7:0] t_r42_c31_12;
  wire [7:0] t_r42_c32_0;
  wire [7:0] t_r42_c32_1;
  wire [7:0] t_r42_c32_2;
  wire [7:0] t_r42_c32_3;
  wire [7:0] t_r42_c32_4;
  wire [7:0] t_r42_c32_5;
  wire [7:0] t_r42_c32_6;
  wire [7:0] t_r42_c32_7;
  wire [7:0] t_r42_c32_8;
  wire [7:0] t_r42_c32_9;
  wire [7:0] t_r42_c32_10;
  wire [7:0] t_r42_c32_11;
  wire [7:0] t_r42_c32_12;
  wire [7:0] t_r42_c33_0;
  wire [7:0] t_r42_c33_1;
  wire [7:0] t_r42_c33_2;
  wire [7:0] t_r42_c33_3;
  wire [7:0] t_r42_c33_4;
  wire [7:0] t_r42_c33_5;
  wire [7:0] t_r42_c33_6;
  wire [7:0] t_r42_c33_7;
  wire [7:0] t_r42_c33_8;
  wire [7:0] t_r42_c33_9;
  wire [7:0] t_r42_c33_10;
  wire [7:0] t_r42_c33_11;
  wire [7:0] t_r42_c33_12;
  wire [7:0] t_r42_c34_0;
  wire [7:0] t_r42_c34_1;
  wire [7:0] t_r42_c34_2;
  wire [7:0] t_r42_c34_3;
  wire [7:0] t_r42_c34_4;
  wire [7:0] t_r42_c34_5;
  wire [7:0] t_r42_c34_6;
  wire [7:0] t_r42_c34_7;
  wire [7:0] t_r42_c34_8;
  wire [7:0] t_r42_c34_9;
  wire [7:0] t_r42_c34_10;
  wire [7:0] t_r42_c34_11;
  wire [7:0] t_r42_c34_12;
  wire [7:0] t_r42_c35_0;
  wire [7:0] t_r42_c35_1;
  wire [7:0] t_r42_c35_2;
  wire [7:0] t_r42_c35_3;
  wire [7:0] t_r42_c35_4;
  wire [7:0] t_r42_c35_5;
  wire [7:0] t_r42_c35_6;
  wire [7:0] t_r42_c35_7;
  wire [7:0] t_r42_c35_8;
  wire [7:0] t_r42_c35_9;
  wire [7:0] t_r42_c35_10;
  wire [7:0] t_r42_c35_11;
  wire [7:0] t_r42_c35_12;
  wire [7:0] t_r42_c36_0;
  wire [7:0] t_r42_c36_1;
  wire [7:0] t_r42_c36_2;
  wire [7:0] t_r42_c36_3;
  wire [7:0] t_r42_c36_4;
  wire [7:0] t_r42_c36_5;
  wire [7:0] t_r42_c36_6;
  wire [7:0] t_r42_c36_7;
  wire [7:0] t_r42_c36_8;
  wire [7:0] t_r42_c36_9;
  wire [7:0] t_r42_c36_10;
  wire [7:0] t_r42_c36_11;
  wire [7:0] t_r42_c36_12;
  wire [7:0] t_r42_c37_0;
  wire [7:0] t_r42_c37_1;
  wire [7:0] t_r42_c37_2;
  wire [7:0] t_r42_c37_3;
  wire [7:0] t_r42_c37_4;
  wire [7:0] t_r42_c37_5;
  wire [7:0] t_r42_c37_6;
  wire [7:0] t_r42_c37_7;
  wire [7:0] t_r42_c37_8;
  wire [7:0] t_r42_c37_9;
  wire [7:0] t_r42_c37_10;
  wire [7:0] t_r42_c37_11;
  wire [7:0] t_r42_c37_12;
  wire [7:0] t_r42_c38_0;
  wire [7:0] t_r42_c38_1;
  wire [7:0] t_r42_c38_2;
  wire [7:0] t_r42_c38_3;
  wire [7:0] t_r42_c38_4;
  wire [7:0] t_r42_c38_5;
  wire [7:0] t_r42_c38_6;
  wire [7:0] t_r42_c38_7;
  wire [7:0] t_r42_c38_8;
  wire [7:0] t_r42_c38_9;
  wire [7:0] t_r42_c38_10;
  wire [7:0] t_r42_c38_11;
  wire [7:0] t_r42_c38_12;
  wire [7:0] t_r42_c39_0;
  wire [7:0] t_r42_c39_1;
  wire [7:0] t_r42_c39_2;
  wire [7:0] t_r42_c39_3;
  wire [7:0] t_r42_c39_4;
  wire [7:0] t_r42_c39_5;
  wire [7:0] t_r42_c39_6;
  wire [7:0] t_r42_c39_7;
  wire [7:0] t_r42_c39_8;
  wire [7:0] t_r42_c39_9;
  wire [7:0] t_r42_c39_10;
  wire [7:0] t_r42_c39_11;
  wire [7:0] t_r42_c39_12;
  wire [7:0] t_r42_c40_0;
  wire [7:0] t_r42_c40_1;
  wire [7:0] t_r42_c40_2;
  wire [7:0] t_r42_c40_3;
  wire [7:0] t_r42_c40_4;
  wire [7:0] t_r42_c40_5;
  wire [7:0] t_r42_c40_6;
  wire [7:0] t_r42_c40_7;
  wire [7:0] t_r42_c40_8;
  wire [7:0] t_r42_c40_9;
  wire [7:0] t_r42_c40_10;
  wire [7:0] t_r42_c40_11;
  wire [7:0] t_r42_c40_12;
  wire [7:0] t_r42_c41_0;
  wire [7:0] t_r42_c41_1;
  wire [7:0] t_r42_c41_2;
  wire [7:0] t_r42_c41_3;
  wire [7:0] t_r42_c41_4;
  wire [7:0] t_r42_c41_5;
  wire [7:0] t_r42_c41_6;
  wire [7:0] t_r42_c41_7;
  wire [7:0] t_r42_c41_8;
  wire [7:0] t_r42_c41_9;
  wire [7:0] t_r42_c41_10;
  wire [7:0] t_r42_c41_11;
  wire [7:0] t_r42_c41_12;
  wire [7:0] t_r42_c42_0;
  wire [7:0] t_r42_c42_1;
  wire [7:0] t_r42_c42_2;
  wire [7:0] t_r42_c42_3;
  wire [7:0] t_r42_c42_4;
  wire [7:0] t_r42_c42_5;
  wire [7:0] t_r42_c42_6;
  wire [7:0] t_r42_c42_7;
  wire [7:0] t_r42_c42_8;
  wire [7:0] t_r42_c42_9;
  wire [7:0] t_r42_c42_10;
  wire [7:0] t_r42_c42_11;
  wire [7:0] t_r42_c42_12;
  wire [7:0] t_r42_c43_0;
  wire [7:0] t_r42_c43_1;
  wire [7:0] t_r42_c43_2;
  wire [7:0] t_r42_c43_3;
  wire [7:0] t_r42_c43_4;
  wire [7:0] t_r42_c43_5;
  wire [7:0] t_r42_c43_6;
  wire [7:0] t_r42_c43_7;
  wire [7:0] t_r42_c43_8;
  wire [7:0] t_r42_c43_9;
  wire [7:0] t_r42_c43_10;
  wire [7:0] t_r42_c43_11;
  wire [7:0] t_r42_c43_12;
  wire [7:0] t_r42_c44_0;
  wire [7:0] t_r42_c44_1;
  wire [7:0] t_r42_c44_2;
  wire [7:0] t_r42_c44_3;
  wire [7:0] t_r42_c44_4;
  wire [7:0] t_r42_c44_5;
  wire [7:0] t_r42_c44_6;
  wire [7:0] t_r42_c44_7;
  wire [7:0] t_r42_c44_8;
  wire [7:0] t_r42_c44_9;
  wire [7:0] t_r42_c44_10;
  wire [7:0] t_r42_c44_11;
  wire [7:0] t_r42_c44_12;
  wire [7:0] t_r42_c45_0;
  wire [7:0] t_r42_c45_1;
  wire [7:0] t_r42_c45_2;
  wire [7:0] t_r42_c45_3;
  wire [7:0] t_r42_c45_4;
  wire [7:0] t_r42_c45_5;
  wire [7:0] t_r42_c45_6;
  wire [7:0] t_r42_c45_7;
  wire [7:0] t_r42_c45_8;
  wire [7:0] t_r42_c45_9;
  wire [7:0] t_r42_c45_10;
  wire [7:0] t_r42_c45_11;
  wire [7:0] t_r42_c45_12;
  wire [7:0] t_r42_c46_0;
  wire [7:0] t_r42_c46_1;
  wire [7:0] t_r42_c46_2;
  wire [7:0] t_r42_c46_3;
  wire [7:0] t_r42_c46_4;
  wire [7:0] t_r42_c46_5;
  wire [7:0] t_r42_c46_6;
  wire [7:0] t_r42_c46_7;
  wire [7:0] t_r42_c46_8;
  wire [7:0] t_r42_c46_9;
  wire [7:0] t_r42_c46_10;
  wire [7:0] t_r42_c46_11;
  wire [7:0] t_r42_c46_12;
  wire [7:0] t_r42_c47_0;
  wire [7:0] t_r42_c47_1;
  wire [7:0] t_r42_c47_2;
  wire [7:0] t_r42_c47_3;
  wire [7:0] t_r42_c47_4;
  wire [7:0] t_r42_c47_5;
  wire [7:0] t_r42_c47_6;
  wire [7:0] t_r42_c47_7;
  wire [7:0] t_r42_c47_8;
  wire [7:0] t_r42_c47_9;
  wire [7:0] t_r42_c47_10;
  wire [7:0] t_r42_c47_11;
  wire [7:0] t_r42_c47_12;
  wire [7:0] t_r42_c48_0;
  wire [7:0] t_r42_c48_1;
  wire [7:0] t_r42_c48_2;
  wire [7:0] t_r42_c48_3;
  wire [7:0] t_r42_c48_4;
  wire [7:0] t_r42_c48_5;
  wire [7:0] t_r42_c48_6;
  wire [7:0] t_r42_c48_7;
  wire [7:0] t_r42_c48_8;
  wire [7:0] t_r42_c48_9;
  wire [7:0] t_r42_c48_10;
  wire [7:0] t_r42_c48_11;
  wire [7:0] t_r42_c48_12;
  wire [7:0] t_r42_c49_0;
  wire [7:0] t_r42_c49_1;
  wire [7:0] t_r42_c49_2;
  wire [7:0] t_r42_c49_3;
  wire [7:0] t_r42_c49_4;
  wire [7:0] t_r42_c49_5;
  wire [7:0] t_r42_c49_6;
  wire [7:0] t_r42_c49_7;
  wire [7:0] t_r42_c49_8;
  wire [7:0] t_r42_c49_9;
  wire [7:0] t_r42_c49_10;
  wire [7:0] t_r42_c49_11;
  wire [7:0] t_r42_c49_12;
  wire [7:0] t_r42_c50_0;
  wire [7:0] t_r42_c50_1;
  wire [7:0] t_r42_c50_2;
  wire [7:0] t_r42_c50_3;
  wire [7:0] t_r42_c50_4;
  wire [7:0] t_r42_c50_5;
  wire [7:0] t_r42_c50_6;
  wire [7:0] t_r42_c50_7;
  wire [7:0] t_r42_c50_8;
  wire [7:0] t_r42_c50_9;
  wire [7:0] t_r42_c50_10;
  wire [7:0] t_r42_c50_11;
  wire [7:0] t_r42_c50_12;
  wire [7:0] t_r42_c51_0;
  wire [7:0] t_r42_c51_1;
  wire [7:0] t_r42_c51_2;
  wire [7:0] t_r42_c51_3;
  wire [7:0] t_r42_c51_4;
  wire [7:0] t_r42_c51_5;
  wire [7:0] t_r42_c51_6;
  wire [7:0] t_r42_c51_7;
  wire [7:0] t_r42_c51_8;
  wire [7:0] t_r42_c51_9;
  wire [7:0] t_r42_c51_10;
  wire [7:0] t_r42_c51_11;
  wire [7:0] t_r42_c51_12;
  wire [7:0] t_r42_c52_0;
  wire [7:0] t_r42_c52_1;
  wire [7:0] t_r42_c52_2;
  wire [7:0] t_r42_c52_3;
  wire [7:0] t_r42_c52_4;
  wire [7:0] t_r42_c52_5;
  wire [7:0] t_r42_c52_6;
  wire [7:0] t_r42_c52_7;
  wire [7:0] t_r42_c52_8;
  wire [7:0] t_r42_c52_9;
  wire [7:0] t_r42_c52_10;
  wire [7:0] t_r42_c52_11;
  wire [7:0] t_r42_c52_12;
  wire [7:0] t_r42_c53_0;
  wire [7:0] t_r42_c53_1;
  wire [7:0] t_r42_c53_2;
  wire [7:0] t_r42_c53_3;
  wire [7:0] t_r42_c53_4;
  wire [7:0] t_r42_c53_5;
  wire [7:0] t_r42_c53_6;
  wire [7:0] t_r42_c53_7;
  wire [7:0] t_r42_c53_8;
  wire [7:0] t_r42_c53_9;
  wire [7:0] t_r42_c53_10;
  wire [7:0] t_r42_c53_11;
  wire [7:0] t_r42_c53_12;
  wire [7:0] t_r42_c54_0;
  wire [7:0] t_r42_c54_1;
  wire [7:0] t_r42_c54_2;
  wire [7:0] t_r42_c54_3;
  wire [7:0] t_r42_c54_4;
  wire [7:0] t_r42_c54_5;
  wire [7:0] t_r42_c54_6;
  wire [7:0] t_r42_c54_7;
  wire [7:0] t_r42_c54_8;
  wire [7:0] t_r42_c54_9;
  wire [7:0] t_r42_c54_10;
  wire [7:0] t_r42_c54_11;
  wire [7:0] t_r42_c54_12;
  wire [7:0] t_r42_c55_0;
  wire [7:0] t_r42_c55_1;
  wire [7:0] t_r42_c55_2;
  wire [7:0] t_r42_c55_3;
  wire [7:0] t_r42_c55_4;
  wire [7:0] t_r42_c55_5;
  wire [7:0] t_r42_c55_6;
  wire [7:0] t_r42_c55_7;
  wire [7:0] t_r42_c55_8;
  wire [7:0] t_r42_c55_9;
  wire [7:0] t_r42_c55_10;
  wire [7:0] t_r42_c55_11;
  wire [7:0] t_r42_c55_12;
  wire [7:0] t_r42_c56_0;
  wire [7:0] t_r42_c56_1;
  wire [7:0] t_r42_c56_2;
  wire [7:0] t_r42_c56_3;
  wire [7:0] t_r42_c56_4;
  wire [7:0] t_r42_c56_5;
  wire [7:0] t_r42_c56_6;
  wire [7:0] t_r42_c56_7;
  wire [7:0] t_r42_c56_8;
  wire [7:0] t_r42_c56_9;
  wire [7:0] t_r42_c56_10;
  wire [7:0] t_r42_c56_11;
  wire [7:0] t_r42_c56_12;
  wire [7:0] t_r42_c57_0;
  wire [7:0] t_r42_c57_1;
  wire [7:0] t_r42_c57_2;
  wire [7:0] t_r42_c57_3;
  wire [7:0] t_r42_c57_4;
  wire [7:0] t_r42_c57_5;
  wire [7:0] t_r42_c57_6;
  wire [7:0] t_r42_c57_7;
  wire [7:0] t_r42_c57_8;
  wire [7:0] t_r42_c57_9;
  wire [7:0] t_r42_c57_10;
  wire [7:0] t_r42_c57_11;
  wire [7:0] t_r42_c57_12;
  wire [7:0] t_r42_c58_0;
  wire [7:0] t_r42_c58_1;
  wire [7:0] t_r42_c58_2;
  wire [7:0] t_r42_c58_3;
  wire [7:0] t_r42_c58_4;
  wire [7:0] t_r42_c58_5;
  wire [7:0] t_r42_c58_6;
  wire [7:0] t_r42_c58_7;
  wire [7:0] t_r42_c58_8;
  wire [7:0] t_r42_c58_9;
  wire [7:0] t_r42_c58_10;
  wire [7:0] t_r42_c58_11;
  wire [7:0] t_r42_c58_12;
  wire [7:0] t_r42_c59_0;
  wire [7:0] t_r42_c59_1;
  wire [7:0] t_r42_c59_2;
  wire [7:0] t_r42_c59_3;
  wire [7:0] t_r42_c59_4;
  wire [7:0] t_r42_c59_5;
  wire [7:0] t_r42_c59_6;
  wire [7:0] t_r42_c59_7;
  wire [7:0] t_r42_c59_8;
  wire [7:0] t_r42_c59_9;
  wire [7:0] t_r42_c59_10;
  wire [7:0] t_r42_c59_11;
  wire [7:0] t_r42_c59_12;
  wire [7:0] t_r42_c60_0;
  wire [7:0] t_r42_c60_1;
  wire [7:0] t_r42_c60_2;
  wire [7:0] t_r42_c60_3;
  wire [7:0] t_r42_c60_4;
  wire [7:0] t_r42_c60_5;
  wire [7:0] t_r42_c60_6;
  wire [7:0] t_r42_c60_7;
  wire [7:0] t_r42_c60_8;
  wire [7:0] t_r42_c60_9;
  wire [7:0] t_r42_c60_10;
  wire [7:0] t_r42_c60_11;
  wire [7:0] t_r42_c60_12;
  wire [7:0] t_r42_c61_0;
  wire [7:0] t_r42_c61_1;
  wire [7:0] t_r42_c61_2;
  wire [7:0] t_r42_c61_3;
  wire [7:0] t_r42_c61_4;
  wire [7:0] t_r42_c61_5;
  wire [7:0] t_r42_c61_6;
  wire [7:0] t_r42_c61_7;
  wire [7:0] t_r42_c61_8;
  wire [7:0] t_r42_c61_9;
  wire [7:0] t_r42_c61_10;
  wire [7:0] t_r42_c61_11;
  wire [7:0] t_r42_c61_12;
  wire [7:0] t_r42_c62_0;
  wire [7:0] t_r42_c62_1;
  wire [7:0] t_r42_c62_2;
  wire [7:0] t_r42_c62_3;
  wire [7:0] t_r42_c62_4;
  wire [7:0] t_r42_c62_5;
  wire [7:0] t_r42_c62_6;
  wire [7:0] t_r42_c62_7;
  wire [7:0] t_r42_c62_8;
  wire [7:0] t_r42_c62_9;
  wire [7:0] t_r42_c62_10;
  wire [7:0] t_r42_c62_11;
  wire [7:0] t_r42_c62_12;
  wire [7:0] t_r42_c63_0;
  wire [7:0] t_r42_c63_1;
  wire [7:0] t_r42_c63_2;
  wire [7:0] t_r42_c63_3;
  wire [7:0] t_r42_c63_4;
  wire [7:0] t_r42_c63_5;
  wire [7:0] t_r42_c63_6;
  wire [7:0] t_r42_c63_7;
  wire [7:0] t_r42_c63_8;
  wire [7:0] t_r42_c63_9;
  wire [7:0] t_r42_c63_10;
  wire [7:0] t_r42_c63_11;
  wire [7:0] t_r42_c63_12;
  wire [7:0] t_r42_c64_0;
  wire [7:0] t_r42_c64_1;
  wire [7:0] t_r42_c64_2;
  wire [7:0] t_r42_c64_3;
  wire [7:0] t_r42_c64_4;
  wire [7:0] t_r42_c64_5;
  wire [7:0] t_r42_c64_6;
  wire [7:0] t_r42_c64_7;
  wire [7:0] t_r42_c64_8;
  wire [7:0] t_r42_c64_9;
  wire [7:0] t_r42_c64_10;
  wire [7:0] t_r42_c64_11;
  wire [7:0] t_r42_c64_12;
  wire [7:0] t_r42_c65_0;
  wire [7:0] t_r42_c65_1;
  wire [7:0] t_r42_c65_2;
  wire [7:0] t_r42_c65_3;
  wire [7:0] t_r42_c65_4;
  wire [7:0] t_r42_c65_5;
  wire [7:0] t_r42_c65_6;
  wire [7:0] t_r42_c65_7;
  wire [7:0] t_r42_c65_8;
  wire [7:0] t_r42_c65_9;
  wire [7:0] t_r42_c65_10;
  wire [7:0] t_r42_c65_11;
  wire [7:0] t_r42_c65_12;
  wire [7:0] t_r43_c0_0;
  wire [7:0] t_r43_c0_1;
  wire [7:0] t_r43_c0_2;
  wire [7:0] t_r43_c0_3;
  wire [7:0] t_r43_c0_4;
  wire [7:0] t_r43_c0_5;
  wire [7:0] t_r43_c0_6;
  wire [7:0] t_r43_c0_7;
  wire [7:0] t_r43_c0_8;
  wire [7:0] t_r43_c0_9;
  wire [7:0] t_r43_c0_10;
  wire [7:0] t_r43_c0_11;
  wire [7:0] t_r43_c0_12;
  wire [7:0] t_r43_c1_0;
  wire [7:0] t_r43_c1_1;
  wire [7:0] t_r43_c1_2;
  wire [7:0] t_r43_c1_3;
  wire [7:0] t_r43_c1_4;
  wire [7:0] t_r43_c1_5;
  wire [7:0] t_r43_c1_6;
  wire [7:0] t_r43_c1_7;
  wire [7:0] t_r43_c1_8;
  wire [7:0] t_r43_c1_9;
  wire [7:0] t_r43_c1_10;
  wire [7:0] t_r43_c1_11;
  wire [7:0] t_r43_c1_12;
  wire [7:0] t_r43_c2_0;
  wire [7:0] t_r43_c2_1;
  wire [7:0] t_r43_c2_2;
  wire [7:0] t_r43_c2_3;
  wire [7:0] t_r43_c2_4;
  wire [7:0] t_r43_c2_5;
  wire [7:0] t_r43_c2_6;
  wire [7:0] t_r43_c2_7;
  wire [7:0] t_r43_c2_8;
  wire [7:0] t_r43_c2_9;
  wire [7:0] t_r43_c2_10;
  wire [7:0] t_r43_c2_11;
  wire [7:0] t_r43_c2_12;
  wire [7:0] t_r43_c3_0;
  wire [7:0] t_r43_c3_1;
  wire [7:0] t_r43_c3_2;
  wire [7:0] t_r43_c3_3;
  wire [7:0] t_r43_c3_4;
  wire [7:0] t_r43_c3_5;
  wire [7:0] t_r43_c3_6;
  wire [7:0] t_r43_c3_7;
  wire [7:0] t_r43_c3_8;
  wire [7:0] t_r43_c3_9;
  wire [7:0] t_r43_c3_10;
  wire [7:0] t_r43_c3_11;
  wire [7:0] t_r43_c3_12;
  wire [7:0] t_r43_c4_0;
  wire [7:0] t_r43_c4_1;
  wire [7:0] t_r43_c4_2;
  wire [7:0] t_r43_c4_3;
  wire [7:0] t_r43_c4_4;
  wire [7:0] t_r43_c4_5;
  wire [7:0] t_r43_c4_6;
  wire [7:0] t_r43_c4_7;
  wire [7:0] t_r43_c4_8;
  wire [7:0] t_r43_c4_9;
  wire [7:0] t_r43_c4_10;
  wire [7:0] t_r43_c4_11;
  wire [7:0] t_r43_c4_12;
  wire [7:0] t_r43_c5_0;
  wire [7:0] t_r43_c5_1;
  wire [7:0] t_r43_c5_2;
  wire [7:0] t_r43_c5_3;
  wire [7:0] t_r43_c5_4;
  wire [7:0] t_r43_c5_5;
  wire [7:0] t_r43_c5_6;
  wire [7:0] t_r43_c5_7;
  wire [7:0] t_r43_c5_8;
  wire [7:0] t_r43_c5_9;
  wire [7:0] t_r43_c5_10;
  wire [7:0] t_r43_c5_11;
  wire [7:0] t_r43_c5_12;
  wire [7:0] t_r43_c6_0;
  wire [7:0] t_r43_c6_1;
  wire [7:0] t_r43_c6_2;
  wire [7:0] t_r43_c6_3;
  wire [7:0] t_r43_c6_4;
  wire [7:0] t_r43_c6_5;
  wire [7:0] t_r43_c6_6;
  wire [7:0] t_r43_c6_7;
  wire [7:0] t_r43_c6_8;
  wire [7:0] t_r43_c6_9;
  wire [7:0] t_r43_c6_10;
  wire [7:0] t_r43_c6_11;
  wire [7:0] t_r43_c6_12;
  wire [7:0] t_r43_c7_0;
  wire [7:0] t_r43_c7_1;
  wire [7:0] t_r43_c7_2;
  wire [7:0] t_r43_c7_3;
  wire [7:0] t_r43_c7_4;
  wire [7:0] t_r43_c7_5;
  wire [7:0] t_r43_c7_6;
  wire [7:0] t_r43_c7_7;
  wire [7:0] t_r43_c7_8;
  wire [7:0] t_r43_c7_9;
  wire [7:0] t_r43_c7_10;
  wire [7:0] t_r43_c7_11;
  wire [7:0] t_r43_c7_12;
  wire [7:0] t_r43_c8_0;
  wire [7:0] t_r43_c8_1;
  wire [7:0] t_r43_c8_2;
  wire [7:0] t_r43_c8_3;
  wire [7:0] t_r43_c8_4;
  wire [7:0] t_r43_c8_5;
  wire [7:0] t_r43_c8_6;
  wire [7:0] t_r43_c8_7;
  wire [7:0] t_r43_c8_8;
  wire [7:0] t_r43_c8_9;
  wire [7:0] t_r43_c8_10;
  wire [7:0] t_r43_c8_11;
  wire [7:0] t_r43_c8_12;
  wire [7:0] t_r43_c9_0;
  wire [7:0] t_r43_c9_1;
  wire [7:0] t_r43_c9_2;
  wire [7:0] t_r43_c9_3;
  wire [7:0] t_r43_c9_4;
  wire [7:0] t_r43_c9_5;
  wire [7:0] t_r43_c9_6;
  wire [7:0] t_r43_c9_7;
  wire [7:0] t_r43_c9_8;
  wire [7:0] t_r43_c9_9;
  wire [7:0] t_r43_c9_10;
  wire [7:0] t_r43_c9_11;
  wire [7:0] t_r43_c9_12;
  wire [7:0] t_r43_c10_0;
  wire [7:0] t_r43_c10_1;
  wire [7:0] t_r43_c10_2;
  wire [7:0] t_r43_c10_3;
  wire [7:0] t_r43_c10_4;
  wire [7:0] t_r43_c10_5;
  wire [7:0] t_r43_c10_6;
  wire [7:0] t_r43_c10_7;
  wire [7:0] t_r43_c10_8;
  wire [7:0] t_r43_c10_9;
  wire [7:0] t_r43_c10_10;
  wire [7:0] t_r43_c10_11;
  wire [7:0] t_r43_c10_12;
  wire [7:0] t_r43_c11_0;
  wire [7:0] t_r43_c11_1;
  wire [7:0] t_r43_c11_2;
  wire [7:0] t_r43_c11_3;
  wire [7:0] t_r43_c11_4;
  wire [7:0] t_r43_c11_5;
  wire [7:0] t_r43_c11_6;
  wire [7:0] t_r43_c11_7;
  wire [7:0] t_r43_c11_8;
  wire [7:0] t_r43_c11_9;
  wire [7:0] t_r43_c11_10;
  wire [7:0] t_r43_c11_11;
  wire [7:0] t_r43_c11_12;
  wire [7:0] t_r43_c12_0;
  wire [7:0] t_r43_c12_1;
  wire [7:0] t_r43_c12_2;
  wire [7:0] t_r43_c12_3;
  wire [7:0] t_r43_c12_4;
  wire [7:0] t_r43_c12_5;
  wire [7:0] t_r43_c12_6;
  wire [7:0] t_r43_c12_7;
  wire [7:0] t_r43_c12_8;
  wire [7:0] t_r43_c12_9;
  wire [7:0] t_r43_c12_10;
  wire [7:0] t_r43_c12_11;
  wire [7:0] t_r43_c12_12;
  wire [7:0] t_r43_c13_0;
  wire [7:0] t_r43_c13_1;
  wire [7:0] t_r43_c13_2;
  wire [7:0] t_r43_c13_3;
  wire [7:0] t_r43_c13_4;
  wire [7:0] t_r43_c13_5;
  wire [7:0] t_r43_c13_6;
  wire [7:0] t_r43_c13_7;
  wire [7:0] t_r43_c13_8;
  wire [7:0] t_r43_c13_9;
  wire [7:0] t_r43_c13_10;
  wire [7:0] t_r43_c13_11;
  wire [7:0] t_r43_c13_12;
  wire [7:0] t_r43_c14_0;
  wire [7:0] t_r43_c14_1;
  wire [7:0] t_r43_c14_2;
  wire [7:0] t_r43_c14_3;
  wire [7:0] t_r43_c14_4;
  wire [7:0] t_r43_c14_5;
  wire [7:0] t_r43_c14_6;
  wire [7:0] t_r43_c14_7;
  wire [7:0] t_r43_c14_8;
  wire [7:0] t_r43_c14_9;
  wire [7:0] t_r43_c14_10;
  wire [7:0] t_r43_c14_11;
  wire [7:0] t_r43_c14_12;
  wire [7:0] t_r43_c15_0;
  wire [7:0] t_r43_c15_1;
  wire [7:0] t_r43_c15_2;
  wire [7:0] t_r43_c15_3;
  wire [7:0] t_r43_c15_4;
  wire [7:0] t_r43_c15_5;
  wire [7:0] t_r43_c15_6;
  wire [7:0] t_r43_c15_7;
  wire [7:0] t_r43_c15_8;
  wire [7:0] t_r43_c15_9;
  wire [7:0] t_r43_c15_10;
  wire [7:0] t_r43_c15_11;
  wire [7:0] t_r43_c15_12;
  wire [7:0] t_r43_c16_0;
  wire [7:0] t_r43_c16_1;
  wire [7:0] t_r43_c16_2;
  wire [7:0] t_r43_c16_3;
  wire [7:0] t_r43_c16_4;
  wire [7:0] t_r43_c16_5;
  wire [7:0] t_r43_c16_6;
  wire [7:0] t_r43_c16_7;
  wire [7:0] t_r43_c16_8;
  wire [7:0] t_r43_c16_9;
  wire [7:0] t_r43_c16_10;
  wire [7:0] t_r43_c16_11;
  wire [7:0] t_r43_c16_12;
  wire [7:0] t_r43_c17_0;
  wire [7:0] t_r43_c17_1;
  wire [7:0] t_r43_c17_2;
  wire [7:0] t_r43_c17_3;
  wire [7:0] t_r43_c17_4;
  wire [7:0] t_r43_c17_5;
  wire [7:0] t_r43_c17_6;
  wire [7:0] t_r43_c17_7;
  wire [7:0] t_r43_c17_8;
  wire [7:0] t_r43_c17_9;
  wire [7:0] t_r43_c17_10;
  wire [7:0] t_r43_c17_11;
  wire [7:0] t_r43_c17_12;
  wire [7:0] t_r43_c18_0;
  wire [7:0] t_r43_c18_1;
  wire [7:0] t_r43_c18_2;
  wire [7:0] t_r43_c18_3;
  wire [7:0] t_r43_c18_4;
  wire [7:0] t_r43_c18_5;
  wire [7:0] t_r43_c18_6;
  wire [7:0] t_r43_c18_7;
  wire [7:0] t_r43_c18_8;
  wire [7:0] t_r43_c18_9;
  wire [7:0] t_r43_c18_10;
  wire [7:0] t_r43_c18_11;
  wire [7:0] t_r43_c18_12;
  wire [7:0] t_r43_c19_0;
  wire [7:0] t_r43_c19_1;
  wire [7:0] t_r43_c19_2;
  wire [7:0] t_r43_c19_3;
  wire [7:0] t_r43_c19_4;
  wire [7:0] t_r43_c19_5;
  wire [7:0] t_r43_c19_6;
  wire [7:0] t_r43_c19_7;
  wire [7:0] t_r43_c19_8;
  wire [7:0] t_r43_c19_9;
  wire [7:0] t_r43_c19_10;
  wire [7:0] t_r43_c19_11;
  wire [7:0] t_r43_c19_12;
  wire [7:0] t_r43_c20_0;
  wire [7:0] t_r43_c20_1;
  wire [7:0] t_r43_c20_2;
  wire [7:0] t_r43_c20_3;
  wire [7:0] t_r43_c20_4;
  wire [7:0] t_r43_c20_5;
  wire [7:0] t_r43_c20_6;
  wire [7:0] t_r43_c20_7;
  wire [7:0] t_r43_c20_8;
  wire [7:0] t_r43_c20_9;
  wire [7:0] t_r43_c20_10;
  wire [7:0] t_r43_c20_11;
  wire [7:0] t_r43_c20_12;
  wire [7:0] t_r43_c21_0;
  wire [7:0] t_r43_c21_1;
  wire [7:0] t_r43_c21_2;
  wire [7:0] t_r43_c21_3;
  wire [7:0] t_r43_c21_4;
  wire [7:0] t_r43_c21_5;
  wire [7:0] t_r43_c21_6;
  wire [7:0] t_r43_c21_7;
  wire [7:0] t_r43_c21_8;
  wire [7:0] t_r43_c21_9;
  wire [7:0] t_r43_c21_10;
  wire [7:0] t_r43_c21_11;
  wire [7:0] t_r43_c21_12;
  wire [7:0] t_r43_c22_0;
  wire [7:0] t_r43_c22_1;
  wire [7:0] t_r43_c22_2;
  wire [7:0] t_r43_c22_3;
  wire [7:0] t_r43_c22_4;
  wire [7:0] t_r43_c22_5;
  wire [7:0] t_r43_c22_6;
  wire [7:0] t_r43_c22_7;
  wire [7:0] t_r43_c22_8;
  wire [7:0] t_r43_c22_9;
  wire [7:0] t_r43_c22_10;
  wire [7:0] t_r43_c22_11;
  wire [7:0] t_r43_c22_12;
  wire [7:0] t_r43_c23_0;
  wire [7:0] t_r43_c23_1;
  wire [7:0] t_r43_c23_2;
  wire [7:0] t_r43_c23_3;
  wire [7:0] t_r43_c23_4;
  wire [7:0] t_r43_c23_5;
  wire [7:0] t_r43_c23_6;
  wire [7:0] t_r43_c23_7;
  wire [7:0] t_r43_c23_8;
  wire [7:0] t_r43_c23_9;
  wire [7:0] t_r43_c23_10;
  wire [7:0] t_r43_c23_11;
  wire [7:0] t_r43_c23_12;
  wire [7:0] t_r43_c24_0;
  wire [7:0] t_r43_c24_1;
  wire [7:0] t_r43_c24_2;
  wire [7:0] t_r43_c24_3;
  wire [7:0] t_r43_c24_4;
  wire [7:0] t_r43_c24_5;
  wire [7:0] t_r43_c24_6;
  wire [7:0] t_r43_c24_7;
  wire [7:0] t_r43_c24_8;
  wire [7:0] t_r43_c24_9;
  wire [7:0] t_r43_c24_10;
  wire [7:0] t_r43_c24_11;
  wire [7:0] t_r43_c24_12;
  wire [7:0] t_r43_c25_0;
  wire [7:0] t_r43_c25_1;
  wire [7:0] t_r43_c25_2;
  wire [7:0] t_r43_c25_3;
  wire [7:0] t_r43_c25_4;
  wire [7:0] t_r43_c25_5;
  wire [7:0] t_r43_c25_6;
  wire [7:0] t_r43_c25_7;
  wire [7:0] t_r43_c25_8;
  wire [7:0] t_r43_c25_9;
  wire [7:0] t_r43_c25_10;
  wire [7:0] t_r43_c25_11;
  wire [7:0] t_r43_c25_12;
  wire [7:0] t_r43_c26_0;
  wire [7:0] t_r43_c26_1;
  wire [7:0] t_r43_c26_2;
  wire [7:0] t_r43_c26_3;
  wire [7:0] t_r43_c26_4;
  wire [7:0] t_r43_c26_5;
  wire [7:0] t_r43_c26_6;
  wire [7:0] t_r43_c26_7;
  wire [7:0] t_r43_c26_8;
  wire [7:0] t_r43_c26_9;
  wire [7:0] t_r43_c26_10;
  wire [7:0] t_r43_c26_11;
  wire [7:0] t_r43_c26_12;
  wire [7:0] t_r43_c27_0;
  wire [7:0] t_r43_c27_1;
  wire [7:0] t_r43_c27_2;
  wire [7:0] t_r43_c27_3;
  wire [7:0] t_r43_c27_4;
  wire [7:0] t_r43_c27_5;
  wire [7:0] t_r43_c27_6;
  wire [7:0] t_r43_c27_7;
  wire [7:0] t_r43_c27_8;
  wire [7:0] t_r43_c27_9;
  wire [7:0] t_r43_c27_10;
  wire [7:0] t_r43_c27_11;
  wire [7:0] t_r43_c27_12;
  wire [7:0] t_r43_c28_0;
  wire [7:0] t_r43_c28_1;
  wire [7:0] t_r43_c28_2;
  wire [7:0] t_r43_c28_3;
  wire [7:0] t_r43_c28_4;
  wire [7:0] t_r43_c28_5;
  wire [7:0] t_r43_c28_6;
  wire [7:0] t_r43_c28_7;
  wire [7:0] t_r43_c28_8;
  wire [7:0] t_r43_c28_9;
  wire [7:0] t_r43_c28_10;
  wire [7:0] t_r43_c28_11;
  wire [7:0] t_r43_c28_12;
  wire [7:0] t_r43_c29_0;
  wire [7:0] t_r43_c29_1;
  wire [7:0] t_r43_c29_2;
  wire [7:0] t_r43_c29_3;
  wire [7:0] t_r43_c29_4;
  wire [7:0] t_r43_c29_5;
  wire [7:0] t_r43_c29_6;
  wire [7:0] t_r43_c29_7;
  wire [7:0] t_r43_c29_8;
  wire [7:0] t_r43_c29_9;
  wire [7:0] t_r43_c29_10;
  wire [7:0] t_r43_c29_11;
  wire [7:0] t_r43_c29_12;
  wire [7:0] t_r43_c30_0;
  wire [7:0] t_r43_c30_1;
  wire [7:0] t_r43_c30_2;
  wire [7:0] t_r43_c30_3;
  wire [7:0] t_r43_c30_4;
  wire [7:0] t_r43_c30_5;
  wire [7:0] t_r43_c30_6;
  wire [7:0] t_r43_c30_7;
  wire [7:0] t_r43_c30_8;
  wire [7:0] t_r43_c30_9;
  wire [7:0] t_r43_c30_10;
  wire [7:0] t_r43_c30_11;
  wire [7:0] t_r43_c30_12;
  wire [7:0] t_r43_c31_0;
  wire [7:0] t_r43_c31_1;
  wire [7:0] t_r43_c31_2;
  wire [7:0] t_r43_c31_3;
  wire [7:0] t_r43_c31_4;
  wire [7:0] t_r43_c31_5;
  wire [7:0] t_r43_c31_6;
  wire [7:0] t_r43_c31_7;
  wire [7:0] t_r43_c31_8;
  wire [7:0] t_r43_c31_9;
  wire [7:0] t_r43_c31_10;
  wire [7:0] t_r43_c31_11;
  wire [7:0] t_r43_c31_12;
  wire [7:0] t_r43_c32_0;
  wire [7:0] t_r43_c32_1;
  wire [7:0] t_r43_c32_2;
  wire [7:0] t_r43_c32_3;
  wire [7:0] t_r43_c32_4;
  wire [7:0] t_r43_c32_5;
  wire [7:0] t_r43_c32_6;
  wire [7:0] t_r43_c32_7;
  wire [7:0] t_r43_c32_8;
  wire [7:0] t_r43_c32_9;
  wire [7:0] t_r43_c32_10;
  wire [7:0] t_r43_c32_11;
  wire [7:0] t_r43_c32_12;
  wire [7:0] t_r43_c33_0;
  wire [7:0] t_r43_c33_1;
  wire [7:0] t_r43_c33_2;
  wire [7:0] t_r43_c33_3;
  wire [7:0] t_r43_c33_4;
  wire [7:0] t_r43_c33_5;
  wire [7:0] t_r43_c33_6;
  wire [7:0] t_r43_c33_7;
  wire [7:0] t_r43_c33_8;
  wire [7:0] t_r43_c33_9;
  wire [7:0] t_r43_c33_10;
  wire [7:0] t_r43_c33_11;
  wire [7:0] t_r43_c33_12;
  wire [7:0] t_r43_c34_0;
  wire [7:0] t_r43_c34_1;
  wire [7:0] t_r43_c34_2;
  wire [7:0] t_r43_c34_3;
  wire [7:0] t_r43_c34_4;
  wire [7:0] t_r43_c34_5;
  wire [7:0] t_r43_c34_6;
  wire [7:0] t_r43_c34_7;
  wire [7:0] t_r43_c34_8;
  wire [7:0] t_r43_c34_9;
  wire [7:0] t_r43_c34_10;
  wire [7:0] t_r43_c34_11;
  wire [7:0] t_r43_c34_12;
  wire [7:0] t_r43_c35_0;
  wire [7:0] t_r43_c35_1;
  wire [7:0] t_r43_c35_2;
  wire [7:0] t_r43_c35_3;
  wire [7:0] t_r43_c35_4;
  wire [7:0] t_r43_c35_5;
  wire [7:0] t_r43_c35_6;
  wire [7:0] t_r43_c35_7;
  wire [7:0] t_r43_c35_8;
  wire [7:0] t_r43_c35_9;
  wire [7:0] t_r43_c35_10;
  wire [7:0] t_r43_c35_11;
  wire [7:0] t_r43_c35_12;
  wire [7:0] t_r43_c36_0;
  wire [7:0] t_r43_c36_1;
  wire [7:0] t_r43_c36_2;
  wire [7:0] t_r43_c36_3;
  wire [7:0] t_r43_c36_4;
  wire [7:0] t_r43_c36_5;
  wire [7:0] t_r43_c36_6;
  wire [7:0] t_r43_c36_7;
  wire [7:0] t_r43_c36_8;
  wire [7:0] t_r43_c36_9;
  wire [7:0] t_r43_c36_10;
  wire [7:0] t_r43_c36_11;
  wire [7:0] t_r43_c36_12;
  wire [7:0] t_r43_c37_0;
  wire [7:0] t_r43_c37_1;
  wire [7:0] t_r43_c37_2;
  wire [7:0] t_r43_c37_3;
  wire [7:0] t_r43_c37_4;
  wire [7:0] t_r43_c37_5;
  wire [7:0] t_r43_c37_6;
  wire [7:0] t_r43_c37_7;
  wire [7:0] t_r43_c37_8;
  wire [7:0] t_r43_c37_9;
  wire [7:0] t_r43_c37_10;
  wire [7:0] t_r43_c37_11;
  wire [7:0] t_r43_c37_12;
  wire [7:0] t_r43_c38_0;
  wire [7:0] t_r43_c38_1;
  wire [7:0] t_r43_c38_2;
  wire [7:0] t_r43_c38_3;
  wire [7:0] t_r43_c38_4;
  wire [7:0] t_r43_c38_5;
  wire [7:0] t_r43_c38_6;
  wire [7:0] t_r43_c38_7;
  wire [7:0] t_r43_c38_8;
  wire [7:0] t_r43_c38_9;
  wire [7:0] t_r43_c38_10;
  wire [7:0] t_r43_c38_11;
  wire [7:0] t_r43_c38_12;
  wire [7:0] t_r43_c39_0;
  wire [7:0] t_r43_c39_1;
  wire [7:0] t_r43_c39_2;
  wire [7:0] t_r43_c39_3;
  wire [7:0] t_r43_c39_4;
  wire [7:0] t_r43_c39_5;
  wire [7:0] t_r43_c39_6;
  wire [7:0] t_r43_c39_7;
  wire [7:0] t_r43_c39_8;
  wire [7:0] t_r43_c39_9;
  wire [7:0] t_r43_c39_10;
  wire [7:0] t_r43_c39_11;
  wire [7:0] t_r43_c39_12;
  wire [7:0] t_r43_c40_0;
  wire [7:0] t_r43_c40_1;
  wire [7:0] t_r43_c40_2;
  wire [7:0] t_r43_c40_3;
  wire [7:0] t_r43_c40_4;
  wire [7:0] t_r43_c40_5;
  wire [7:0] t_r43_c40_6;
  wire [7:0] t_r43_c40_7;
  wire [7:0] t_r43_c40_8;
  wire [7:0] t_r43_c40_9;
  wire [7:0] t_r43_c40_10;
  wire [7:0] t_r43_c40_11;
  wire [7:0] t_r43_c40_12;
  wire [7:0] t_r43_c41_0;
  wire [7:0] t_r43_c41_1;
  wire [7:0] t_r43_c41_2;
  wire [7:0] t_r43_c41_3;
  wire [7:0] t_r43_c41_4;
  wire [7:0] t_r43_c41_5;
  wire [7:0] t_r43_c41_6;
  wire [7:0] t_r43_c41_7;
  wire [7:0] t_r43_c41_8;
  wire [7:0] t_r43_c41_9;
  wire [7:0] t_r43_c41_10;
  wire [7:0] t_r43_c41_11;
  wire [7:0] t_r43_c41_12;
  wire [7:0] t_r43_c42_0;
  wire [7:0] t_r43_c42_1;
  wire [7:0] t_r43_c42_2;
  wire [7:0] t_r43_c42_3;
  wire [7:0] t_r43_c42_4;
  wire [7:0] t_r43_c42_5;
  wire [7:0] t_r43_c42_6;
  wire [7:0] t_r43_c42_7;
  wire [7:0] t_r43_c42_8;
  wire [7:0] t_r43_c42_9;
  wire [7:0] t_r43_c42_10;
  wire [7:0] t_r43_c42_11;
  wire [7:0] t_r43_c42_12;
  wire [7:0] t_r43_c43_0;
  wire [7:0] t_r43_c43_1;
  wire [7:0] t_r43_c43_2;
  wire [7:0] t_r43_c43_3;
  wire [7:0] t_r43_c43_4;
  wire [7:0] t_r43_c43_5;
  wire [7:0] t_r43_c43_6;
  wire [7:0] t_r43_c43_7;
  wire [7:0] t_r43_c43_8;
  wire [7:0] t_r43_c43_9;
  wire [7:0] t_r43_c43_10;
  wire [7:0] t_r43_c43_11;
  wire [7:0] t_r43_c43_12;
  wire [7:0] t_r43_c44_0;
  wire [7:0] t_r43_c44_1;
  wire [7:0] t_r43_c44_2;
  wire [7:0] t_r43_c44_3;
  wire [7:0] t_r43_c44_4;
  wire [7:0] t_r43_c44_5;
  wire [7:0] t_r43_c44_6;
  wire [7:0] t_r43_c44_7;
  wire [7:0] t_r43_c44_8;
  wire [7:0] t_r43_c44_9;
  wire [7:0] t_r43_c44_10;
  wire [7:0] t_r43_c44_11;
  wire [7:0] t_r43_c44_12;
  wire [7:0] t_r43_c45_0;
  wire [7:0] t_r43_c45_1;
  wire [7:0] t_r43_c45_2;
  wire [7:0] t_r43_c45_3;
  wire [7:0] t_r43_c45_4;
  wire [7:0] t_r43_c45_5;
  wire [7:0] t_r43_c45_6;
  wire [7:0] t_r43_c45_7;
  wire [7:0] t_r43_c45_8;
  wire [7:0] t_r43_c45_9;
  wire [7:0] t_r43_c45_10;
  wire [7:0] t_r43_c45_11;
  wire [7:0] t_r43_c45_12;
  wire [7:0] t_r43_c46_0;
  wire [7:0] t_r43_c46_1;
  wire [7:0] t_r43_c46_2;
  wire [7:0] t_r43_c46_3;
  wire [7:0] t_r43_c46_4;
  wire [7:0] t_r43_c46_5;
  wire [7:0] t_r43_c46_6;
  wire [7:0] t_r43_c46_7;
  wire [7:0] t_r43_c46_8;
  wire [7:0] t_r43_c46_9;
  wire [7:0] t_r43_c46_10;
  wire [7:0] t_r43_c46_11;
  wire [7:0] t_r43_c46_12;
  wire [7:0] t_r43_c47_0;
  wire [7:0] t_r43_c47_1;
  wire [7:0] t_r43_c47_2;
  wire [7:0] t_r43_c47_3;
  wire [7:0] t_r43_c47_4;
  wire [7:0] t_r43_c47_5;
  wire [7:0] t_r43_c47_6;
  wire [7:0] t_r43_c47_7;
  wire [7:0] t_r43_c47_8;
  wire [7:0] t_r43_c47_9;
  wire [7:0] t_r43_c47_10;
  wire [7:0] t_r43_c47_11;
  wire [7:0] t_r43_c47_12;
  wire [7:0] t_r43_c48_0;
  wire [7:0] t_r43_c48_1;
  wire [7:0] t_r43_c48_2;
  wire [7:0] t_r43_c48_3;
  wire [7:0] t_r43_c48_4;
  wire [7:0] t_r43_c48_5;
  wire [7:0] t_r43_c48_6;
  wire [7:0] t_r43_c48_7;
  wire [7:0] t_r43_c48_8;
  wire [7:0] t_r43_c48_9;
  wire [7:0] t_r43_c48_10;
  wire [7:0] t_r43_c48_11;
  wire [7:0] t_r43_c48_12;
  wire [7:0] t_r43_c49_0;
  wire [7:0] t_r43_c49_1;
  wire [7:0] t_r43_c49_2;
  wire [7:0] t_r43_c49_3;
  wire [7:0] t_r43_c49_4;
  wire [7:0] t_r43_c49_5;
  wire [7:0] t_r43_c49_6;
  wire [7:0] t_r43_c49_7;
  wire [7:0] t_r43_c49_8;
  wire [7:0] t_r43_c49_9;
  wire [7:0] t_r43_c49_10;
  wire [7:0] t_r43_c49_11;
  wire [7:0] t_r43_c49_12;
  wire [7:0] t_r43_c50_0;
  wire [7:0] t_r43_c50_1;
  wire [7:0] t_r43_c50_2;
  wire [7:0] t_r43_c50_3;
  wire [7:0] t_r43_c50_4;
  wire [7:0] t_r43_c50_5;
  wire [7:0] t_r43_c50_6;
  wire [7:0] t_r43_c50_7;
  wire [7:0] t_r43_c50_8;
  wire [7:0] t_r43_c50_9;
  wire [7:0] t_r43_c50_10;
  wire [7:0] t_r43_c50_11;
  wire [7:0] t_r43_c50_12;
  wire [7:0] t_r43_c51_0;
  wire [7:0] t_r43_c51_1;
  wire [7:0] t_r43_c51_2;
  wire [7:0] t_r43_c51_3;
  wire [7:0] t_r43_c51_4;
  wire [7:0] t_r43_c51_5;
  wire [7:0] t_r43_c51_6;
  wire [7:0] t_r43_c51_7;
  wire [7:0] t_r43_c51_8;
  wire [7:0] t_r43_c51_9;
  wire [7:0] t_r43_c51_10;
  wire [7:0] t_r43_c51_11;
  wire [7:0] t_r43_c51_12;
  wire [7:0] t_r43_c52_0;
  wire [7:0] t_r43_c52_1;
  wire [7:0] t_r43_c52_2;
  wire [7:0] t_r43_c52_3;
  wire [7:0] t_r43_c52_4;
  wire [7:0] t_r43_c52_5;
  wire [7:0] t_r43_c52_6;
  wire [7:0] t_r43_c52_7;
  wire [7:0] t_r43_c52_8;
  wire [7:0] t_r43_c52_9;
  wire [7:0] t_r43_c52_10;
  wire [7:0] t_r43_c52_11;
  wire [7:0] t_r43_c52_12;
  wire [7:0] t_r43_c53_0;
  wire [7:0] t_r43_c53_1;
  wire [7:0] t_r43_c53_2;
  wire [7:0] t_r43_c53_3;
  wire [7:0] t_r43_c53_4;
  wire [7:0] t_r43_c53_5;
  wire [7:0] t_r43_c53_6;
  wire [7:0] t_r43_c53_7;
  wire [7:0] t_r43_c53_8;
  wire [7:0] t_r43_c53_9;
  wire [7:0] t_r43_c53_10;
  wire [7:0] t_r43_c53_11;
  wire [7:0] t_r43_c53_12;
  wire [7:0] t_r43_c54_0;
  wire [7:0] t_r43_c54_1;
  wire [7:0] t_r43_c54_2;
  wire [7:0] t_r43_c54_3;
  wire [7:0] t_r43_c54_4;
  wire [7:0] t_r43_c54_5;
  wire [7:0] t_r43_c54_6;
  wire [7:0] t_r43_c54_7;
  wire [7:0] t_r43_c54_8;
  wire [7:0] t_r43_c54_9;
  wire [7:0] t_r43_c54_10;
  wire [7:0] t_r43_c54_11;
  wire [7:0] t_r43_c54_12;
  wire [7:0] t_r43_c55_0;
  wire [7:0] t_r43_c55_1;
  wire [7:0] t_r43_c55_2;
  wire [7:0] t_r43_c55_3;
  wire [7:0] t_r43_c55_4;
  wire [7:0] t_r43_c55_5;
  wire [7:0] t_r43_c55_6;
  wire [7:0] t_r43_c55_7;
  wire [7:0] t_r43_c55_8;
  wire [7:0] t_r43_c55_9;
  wire [7:0] t_r43_c55_10;
  wire [7:0] t_r43_c55_11;
  wire [7:0] t_r43_c55_12;
  wire [7:0] t_r43_c56_0;
  wire [7:0] t_r43_c56_1;
  wire [7:0] t_r43_c56_2;
  wire [7:0] t_r43_c56_3;
  wire [7:0] t_r43_c56_4;
  wire [7:0] t_r43_c56_5;
  wire [7:0] t_r43_c56_6;
  wire [7:0] t_r43_c56_7;
  wire [7:0] t_r43_c56_8;
  wire [7:0] t_r43_c56_9;
  wire [7:0] t_r43_c56_10;
  wire [7:0] t_r43_c56_11;
  wire [7:0] t_r43_c56_12;
  wire [7:0] t_r43_c57_0;
  wire [7:0] t_r43_c57_1;
  wire [7:0] t_r43_c57_2;
  wire [7:0] t_r43_c57_3;
  wire [7:0] t_r43_c57_4;
  wire [7:0] t_r43_c57_5;
  wire [7:0] t_r43_c57_6;
  wire [7:0] t_r43_c57_7;
  wire [7:0] t_r43_c57_8;
  wire [7:0] t_r43_c57_9;
  wire [7:0] t_r43_c57_10;
  wire [7:0] t_r43_c57_11;
  wire [7:0] t_r43_c57_12;
  wire [7:0] t_r43_c58_0;
  wire [7:0] t_r43_c58_1;
  wire [7:0] t_r43_c58_2;
  wire [7:0] t_r43_c58_3;
  wire [7:0] t_r43_c58_4;
  wire [7:0] t_r43_c58_5;
  wire [7:0] t_r43_c58_6;
  wire [7:0] t_r43_c58_7;
  wire [7:0] t_r43_c58_8;
  wire [7:0] t_r43_c58_9;
  wire [7:0] t_r43_c58_10;
  wire [7:0] t_r43_c58_11;
  wire [7:0] t_r43_c58_12;
  wire [7:0] t_r43_c59_0;
  wire [7:0] t_r43_c59_1;
  wire [7:0] t_r43_c59_2;
  wire [7:0] t_r43_c59_3;
  wire [7:0] t_r43_c59_4;
  wire [7:0] t_r43_c59_5;
  wire [7:0] t_r43_c59_6;
  wire [7:0] t_r43_c59_7;
  wire [7:0] t_r43_c59_8;
  wire [7:0] t_r43_c59_9;
  wire [7:0] t_r43_c59_10;
  wire [7:0] t_r43_c59_11;
  wire [7:0] t_r43_c59_12;
  wire [7:0] t_r43_c60_0;
  wire [7:0] t_r43_c60_1;
  wire [7:0] t_r43_c60_2;
  wire [7:0] t_r43_c60_3;
  wire [7:0] t_r43_c60_4;
  wire [7:0] t_r43_c60_5;
  wire [7:0] t_r43_c60_6;
  wire [7:0] t_r43_c60_7;
  wire [7:0] t_r43_c60_8;
  wire [7:0] t_r43_c60_9;
  wire [7:0] t_r43_c60_10;
  wire [7:0] t_r43_c60_11;
  wire [7:0] t_r43_c60_12;
  wire [7:0] t_r43_c61_0;
  wire [7:0] t_r43_c61_1;
  wire [7:0] t_r43_c61_2;
  wire [7:0] t_r43_c61_3;
  wire [7:0] t_r43_c61_4;
  wire [7:0] t_r43_c61_5;
  wire [7:0] t_r43_c61_6;
  wire [7:0] t_r43_c61_7;
  wire [7:0] t_r43_c61_8;
  wire [7:0] t_r43_c61_9;
  wire [7:0] t_r43_c61_10;
  wire [7:0] t_r43_c61_11;
  wire [7:0] t_r43_c61_12;
  wire [7:0] t_r43_c62_0;
  wire [7:0] t_r43_c62_1;
  wire [7:0] t_r43_c62_2;
  wire [7:0] t_r43_c62_3;
  wire [7:0] t_r43_c62_4;
  wire [7:0] t_r43_c62_5;
  wire [7:0] t_r43_c62_6;
  wire [7:0] t_r43_c62_7;
  wire [7:0] t_r43_c62_8;
  wire [7:0] t_r43_c62_9;
  wire [7:0] t_r43_c62_10;
  wire [7:0] t_r43_c62_11;
  wire [7:0] t_r43_c62_12;
  wire [7:0] t_r43_c63_0;
  wire [7:0] t_r43_c63_1;
  wire [7:0] t_r43_c63_2;
  wire [7:0] t_r43_c63_3;
  wire [7:0] t_r43_c63_4;
  wire [7:0] t_r43_c63_5;
  wire [7:0] t_r43_c63_6;
  wire [7:0] t_r43_c63_7;
  wire [7:0] t_r43_c63_8;
  wire [7:0] t_r43_c63_9;
  wire [7:0] t_r43_c63_10;
  wire [7:0] t_r43_c63_11;
  wire [7:0] t_r43_c63_12;
  wire [7:0] t_r43_c64_0;
  wire [7:0] t_r43_c64_1;
  wire [7:0] t_r43_c64_2;
  wire [7:0] t_r43_c64_3;
  wire [7:0] t_r43_c64_4;
  wire [7:0] t_r43_c64_5;
  wire [7:0] t_r43_c64_6;
  wire [7:0] t_r43_c64_7;
  wire [7:0] t_r43_c64_8;
  wire [7:0] t_r43_c64_9;
  wire [7:0] t_r43_c64_10;
  wire [7:0] t_r43_c64_11;
  wire [7:0] t_r43_c64_12;
  wire [7:0] t_r43_c65_0;
  wire [7:0] t_r43_c65_1;
  wire [7:0] t_r43_c65_2;
  wire [7:0] t_r43_c65_3;
  wire [7:0] t_r43_c65_4;
  wire [7:0] t_r43_c65_5;
  wire [7:0] t_r43_c65_6;
  wire [7:0] t_r43_c65_7;
  wire [7:0] t_r43_c65_8;
  wire [7:0] t_r43_c65_9;
  wire [7:0] t_r43_c65_10;
  wire [7:0] t_r43_c65_11;
  wire [7:0] t_r43_c65_12;
  wire [7:0] t_r44_c0_0;
  wire [7:0] t_r44_c0_1;
  wire [7:0] t_r44_c0_2;
  wire [7:0] t_r44_c0_3;
  wire [7:0] t_r44_c0_4;
  wire [7:0] t_r44_c0_5;
  wire [7:0] t_r44_c0_6;
  wire [7:0] t_r44_c0_7;
  wire [7:0] t_r44_c0_8;
  wire [7:0] t_r44_c0_9;
  wire [7:0] t_r44_c0_10;
  wire [7:0] t_r44_c0_11;
  wire [7:0] t_r44_c0_12;
  wire [7:0] t_r44_c1_0;
  wire [7:0] t_r44_c1_1;
  wire [7:0] t_r44_c1_2;
  wire [7:0] t_r44_c1_3;
  wire [7:0] t_r44_c1_4;
  wire [7:0] t_r44_c1_5;
  wire [7:0] t_r44_c1_6;
  wire [7:0] t_r44_c1_7;
  wire [7:0] t_r44_c1_8;
  wire [7:0] t_r44_c1_9;
  wire [7:0] t_r44_c1_10;
  wire [7:0] t_r44_c1_11;
  wire [7:0] t_r44_c1_12;
  wire [7:0] t_r44_c2_0;
  wire [7:0] t_r44_c2_1;
  wire [7:0] t_r44_c2_2;
  wire [7:0] t_r44_c2_3;
  wire [7:0] t_r44_c2_4;
  wire [7:0] t_r44_c2_5;
  wire [7:0] t_r44_c2_6;
  wire [7:0] t_r44_c2_7;
  wire [7:0] t_r44_c2_8;
  wire [7:0] t_r44_c2_9;
  wire [7:0] t_r44_c2_10;
  wire [7:0] t_r44_c2_11;
  wire [7:0] t_r44_c2_12;
  wire [7:0] t_r44_c3_0;
  wire [7:0] t_r44_c3_1;
  wire [7:0] t_r44_c3_2;
  wire [7:0] t_r44_c3_3;
  wire [7:0] t_r44_c3_4;
  wire [7:0] t_r44_c3_5;
  wire [7:0] t_r44_c3_6;
  wire [7:0] t_r44_c3_7;
  wire [7:0] t_r44_c3_8;
  wire [7:0] t_r44_c3_9;
  wire [7:0] t_r44_c3_10;
  wire [7:0] t_r44_c3_11;
  wire [7:0] t_r44_c3_12;
  wire [7:0] t_r44_c4_0;
  wire [7:0] t_r44_c4_1;
  wire [7:0] t_r44_c4_2;
  wire [7:0] t_r44_c4_3;
  wire [7:0] t_r44_c4_4;
  wire [7:0] t_r44_c4_5;
  wire [7:0] t_r44_c4_6;
  wire [7:0] t_r44_c4_7;
  wire [7:0] t_r44_c4_8;
  wire [7:0] t_r44_c4_9;
  wire [7:0] t_r44_c4_10;
  wire [7:0] t_r44_c4_11;
  wire [7:0] t_r44_c4_12;
  wire [7:0] t_r44_c5_0;
  wire [7:0] t_r44_c5_1;
  wire [7:0] t_r44_c5_2;
  wire [7:0] t_r44_c5_3;
  wire [7:0] t_r44_c5_4;
  wire [7:0] t_r44_c5_5;
  wire [7:0] t_r44_c5_6;
  wire [7:0] t_r44_c5_7;
  wire [7:0] t_r44_c5_8;
  wire [7:0] t_r44_c5_9;
  wire [7:0] t_r44_c5_10;
  wire [7:0] t_r44_c5_11;
  wire [7:0] t_r44_c5_12;
  wire [7:0] t_r44_c6_0;
  wire [7:0] t_r44_c6_1;
  wire [7:0] t_r44_c6_2;
  wire [7:0] t_r44_c6_3;
  wire [7:0] t_r44_c6_4;
  wire [7:0] t_r44_c6_5;
  wire [7:0] t_r44_c6_6;
  wire [7:0] t_r44_c6_7;
  wire [7:0] t_r44_c6_8;
  wire [7:0] t_r44_c6_9;
  wire [7:0] t_r44_c6_10;
  wire [7:0] t_r44_c6_11;
  wire [7:0] t_r44_c6_12;
  wire [7:0] t_r44_c7_0;
  wire [7:0] t_r44_c7_1;
  wire [7:0] t_r44_c7_2;
  wire [7:0] t_r44_c7_3;
  wire [7:0] t_r44_c7_4;
  wire [7:0] t_r44_c7_5;
  wire [7:0] t_r44_c7_6;
  wire [7:0] t_r44_c7_7;
  wire [7:0] t_r44_c7_8;
  wire [7:0] t_r44_c7_9;
  wire [7:0] t_r44_c7_10;
  wire [7:0] t_r44_c7_11;
  wire [7:0] t_r44_c7_12;
  wire [7:0] t_r44_c8_0;
  wire [7:0] t_r44_c8_1;
  wire [7:0] t_r44_c8_2;
  wire [7:0] t_r44_c8_3;
  wire [7:0] t_r44_c8_4;
  wire [7:0] t_r44_c8_5;
  wire [7:0] t_r44_c8_6;
  wire [7:0] t_r44_c8_7;
  wire [7:0] t_r44_c8_8;
  wire [7:0] t_r44_c8_9;
  wire [7:0] t_r44_c8_10;
  wire [7:0] t_r44_c8_11;
  wire [7:0] t_r44_c8_12;
  wire [7:0] t_r44_c9_0;
  wire [7:0] t_r44_c9_1;
  wire [7:0] t_r44_c9_2;
  wire [7:0] t_r44_c9_3;
  wire [7:0] t_r44_c9_4;
  wire [7:0] t_r44_c9_5;
  wire [7:0] t_r44_c9_6;
  wire [7:0] t_r44_c9_7;
  wire [7:0] t_r44_c9_8;
  wire [7:0] t_r44_c9_9;
  wire [7:0] t_r44_c9_10;
  wire [7:0] t_r44_c9_11;
  wire [7:0] t_r44_c9_12;
  wire [7:0] t_r44_c10_0;
  wire [7:0] t_r44_c10_1;
  wire [7:0] t_r44_c10_2;
  wire [7:0] t_r44_c10_3;
  wire [7:0] t_r44_c10_4;
  wire [7:0] t_r44_c10_5;
  wire [7:0] t_r44_c10_6;
  wire [7:0] t_r44_c10_7;
  wire [7:0] t_r44_c10_8;
  wire [7:0] t_r44_c10_9;
  wire [7:0] t_r44_c10_10;
  wire [7:0] t_r44_c10_11;
  wire [7:0] t_r44_c10_12;
  wire [7:0] t_r44_c11_0;
  wire [7:0] t_r44_c11_1;
  wire [7:0] t_r44_c11_2;
  wire [7:0] t_r44_c11_3;
  wire [7:0] t_r44_c11_4;
  wire [7:0] t_r44_c11_5;
  wire [7:0] t_r44_c11_6;
  wire [7:0] t_r44_c11_7;
  wire [7:0] t_r44_c11_8;
  wire [7:0] t_r44_c11_9;
  wire [7:0] t_r44_c11_10;
  wire [7:0] t_r44_c11_11;
  wire [7:0] t_r44_c11_12;
  wire [7:0] t_r44_c12_0;
  wire [7:0] t_r44_c12_1;
  wire [7:0] t_r44_c12_2;
  wire [7:0] t_r44_c12_3;
  wire [7:0] t_r44_c12_4;
  wire [7:0] t_r44_c12_5;
  wire [7:0] t_r44_c12_6;
  wire [7:0] t_r44_c12_7;
  wire [7:0] t_r44_c12_8;
  wire [7:0] t_r44_c12_9;
  wire [7:0] t_r44_c12_10;
  wire [7:0] t_r44_c12_11;
  wire [7:0] t_r44_c12_12;
  wire [7:0] t_r44_c13_0;
  wire [7:0] t_r44_c13_1;
  wire [7:0] t_r44_c13_2;
  wire [7:0] t_r44_c13_3;
  wire [7:0] t_r44_c13_4;
  wire [7:0] t_r44_c13_5;
  wire [7:0] t_r44_c13_6;
  wire [7:0] t_r44_c13_7;
  wire [7:0] t_r44_c13_8;
  wire [7:0] t_r44_c13_9;
  wire [7:0] t_r44_c13_10;
  wire [7:0] t_r44_c13_11;
  wire [7:0] t_r44_c13_12;
  wire [7:0] t_r44_c14_0;
  wire [7:0] t_r44_c14_1;
  wire [7:0] t_r44_c14_2;
  wire [7:0] t_r44_c14_3;
  wire [7:0] t_r44_c14_4;
  wire [7:0] t_r44_c14_5;
  wire [7:0] t_r44_c14_6;
  wire [7:0] t_r44_c14_7;
  wire [7:0] t_r44_c14_8;
  wire [7:0] t_r44_c14_9;
  wire [7:0] t_r44_c14_10;
  wire [7:0] t_r44_c14_11;
  wire [7:0] t_r44_c14_12;
  wire [7:0] t_r44_c15_0;
  wire [7:0] t_r44_c15_1;
  wire [7:0] t_r44_c15_2;
  wire [7:0] t_r44_c15_3;
  wire [7:0] t_r44_c15_4;
  wire [7:0] t_r44_c15_5;
  wire [7:0] t_r44_c15_6;
  wire [7:0] t_r44_c15_7;
  wire [7:0] t_r44_c15_8;
  wire [7:0] t_r44_c15_9;
  wire [7:0] t_r44_c15_10;
  wire [7:0] t_r44_c15_11;
  wire [7:0] t_r44_c15_12;
  wire [7:0] t_r44_c16_0;
  wire [7:0] t_r44_c16_1;
  wire [7:0] t_r44_c16_2;
  wire [7:0] t_r44_c16_3;
  wire [7:0] t_r44_c16_4;
  wire [7:0] t_r44_c16_5;
  wire [7:0] t_r44_c16_6;
  wire [7:0] t_r44_c16_7;
  wire [7:0] t_r44_c16_8;
  wire [7:0] t_r44_c16_9;
  wire [7:0] t_r44_c16_10;
  wire [7:0] t_r44_c16_11;
  wire [7:0] t_r44_c16_12;
  wire [7:0] t_r44_c17_0;
  wire [7:0] t_r44_c17_1;
  wire [7:0] t_r44_c17_2;
  wire [7:0] t_r44_c17_3;
  wire [7:0] t_r44_c17_4;
  wire [7:0] t_r44_c17_5;
  wire [7:0] t_r44_c17_6;
  wire [7:0] t_r44_c17_7;
  wire [7:0] t_r44_c17_8;
  wire [7:0] t_r44_c17_9;
  wire [7:0] t_r44_c17_10;
  wire [7:0] t_r44_c17_11;
  wire [7:0] t_r44_c17_12;
  wire [7:0] t_r44_c18_0;
  wire [7:0] t_r44_c18_1;
  wire [7:0] t_r44_c18_2;
  wire [7:0] t_r44_c18_3;
  wire [7:0] t_r44_c18_4;
  wire [7:0] t_r44_c18_5;
  wire [7:0] t_r44_c18_6;
  wire [7:0] t_r44_c18_7;
  wire [7:0] t_r44_c18_8;
  wire [7:0] t_r44_c18_9;
  wire [7:0] t_r44_c18_10;
  wire [7:0] t_r44_c18_11;
  wire [7:0] t_r44_c18_12;
  wire [7:0] t_r44_c19_0;
  wire [7:0] t_r44_c19_1;
  wire [7:0] t_r44_c19_2;
  wire [7:0] t_r44_c19_3;
  wire [7:0] t_r44_c19_4;
  wire [7:0] t_r44_c19_5;
  wire [7:0] t_r44_c19_6;
  wire [7:0] t_r44_c19_7;
  wire [7:0] t_r44_c19_8;
  wire [7:0] t_r44_c19_9;
  wire [7:0] t_r44_c19_10;
  wire [7:0] t_r44_c19_11;
  wire [7:0] t_r44_c19_12;
  wire [7:0] t_r44_c20_0;
  wire [7:0] t_r44_c20_1;
  wire [7:0] t_r44_c20_2;
  wire [7:0] t_r44_c20_3;
  wire [7:0] t_r44_c20_4;
  wire [7:0] t_r44_c20_5;
  wire [7:0] t_r44_c20_6;
  wire [7:0] t_r44_c20_7;
  wire [7:0] t_r44_c20_8;
  wire [7:0] t_r44_c20_9;
  wire [7:0] t_r44_c20_10;
  wire [7:0] t_r44_c20_11;
  wire [7:0] t_r44_c20_12;
  wire [7:0] t_r44_c21_0;
  wire [7:0] t_r44_c21_1;
  wire [7:0] t_r44_c21_2;
  wire [7:0] t_r44_c21_3;
  wire [7:0] t_r44_c21_4;
  wire [7:0] t_r44_c21_5;
  wire [7:0] t_r44_c21_6;
  wire [7:0] t_r44_c21_7;
  wire [7:0] t_r44_c21_8;
  wire [7:0] t_r44_c21_9;
  wire [7:0] t_r44_c21_10;
  wire [7:0] t_r44_c21_11;
  wire [7:0] t_r44_c21_12;
  wire [7:0] t_r44_c22_0;
  wire [7:0] t_r44_c22_1;
  wire [7:0] t_r44_c22_2;
  wire [7:0] t_r44_c22_3;
  wire [7:0] t_r44_c22_4;
  wire [7:0] t_r44_c22_5;
  wire [7:0] t_r44_c22_6;
  wire [7:0] t_r44_c22_7;
  wire [7:0] t_r44_c22_8;
  wire [7:0] t_r44_c22_9;
  wire [7:0] t_r44_c22_10;
  wire [7:0] t_r44_c22_11;
  wire [7:0] t_r44_c22_12;
  wire [7:0] t_r44_c23_0;
  wire [7:0] t_r44_c23_1;
  wire [7:0] t_r44_c23_2;
  wire [7:0] t_r44_c23_3;
  wire [7:0] t_r44_c23_4;
  wire [7:0] t_r44_c23_5;
  wire [7:0] t_r44_c23_6;
  wire [7:0] t_r44_c23_7;
  wire [7:0] t_r44_c23_8;
  wire [7:0] t_r44_c23_9;
  wire [7:0] t_r44_c23_10;
  wire [7:0] t_r44_c23_11;
  wire [7:0] t_r44_c23_12;
  wire [7:0] t_r44_c24_0;
  wire [7:0] t_r44_c24_1;
  wire [7:0] t_r44_c24_2;
  wire [7:0] t_r44_c24_3;
  wire [7:0] t_r44_c24_4;
  wire [7:0] t_r44_c24_5;
  wire [7:0] t_r44_c24_6;
  wire [7:0] t_r44_c24_7;
  wire [7:0] t_r44_c24_8;
  wire [7:0] t_r44_c24_9;
  wire [7:0] t_r44_c24_10;
  wire [7:0] t_r44_c24_11;
  wire [7:0] t_r44_c24_12;
  wire [7:0] t_r44_c25_0;
  wire [7:0] t_r44_c25_1;
  wire [7:0] t_r44_c25_2;
  wire [7:0] t_r44_c25_3;
  wire [7:0] t_r44_c25_4;
  wire [7:0] t_r44_c25_5;
  wire [7:0] t_r44_c25_6;
  wire [7:0] t_r44_c25_7;
  wire [7:0] t_r44_c25_8;
  wire [7:0] t_r44_c25_9;
  wire [7:0] t_r44_c25_10;
  wire [7:0] t_r44_c25_11;
  wire [7:0] t_r44_c25_12;
  wire [7:0] t_r44_c26_0;
  wire [7:0] t_r44_c26_1;
  wire [7:0] t_r44_c26_2;
  wire [7:0] t_r44_c26_3;
  wire [7:0] t_r44_c26_4;
  wire [7:0] t_r44_c26_5;
  wire [7:0] t_r44_c26_6;
  wire [7:0] t_r44_c26_7;
  wire [7:0] t_r44_c26_8;
  wire [7:0] t_r44_c26_9;
  wire [7:0] t_r44_c26_10;
  wire [7:0] t_r44_c26_11;
  wire [7:0] t_r44_c26_12;
  wire [7:0] t_r44_c27_0;
  wire [7:0] t_r44_c27_1;
  wire [7:0] t_r44_c27_2;
  wire [7:0] t_r44_c27_3;
  wire [7:0] t_r44_c27_4;
  wire [7:0] t_r44_c27_5;
  wire [7:0] t_r44_c27_6;
  wire [7:0] t_r44_c27_7;
  wire [7:0] t_r44_c27_8;
  wire [7:0] t_r44_c27_9;
  wire [7:0] t_r44_c27_10;
  wire [7:0] t_r44_c27_11;
  wire [7:0] t_r44_c27_12;
  wire [7:0] t_r44_c28_0;
  wire [7:0] t_r44_c28_1;
  wire [7:0] t_r44_c28_2;
  wire [7:0] t_r44_c28_3;
  wire [7:0] t_r44_c28_4;
  wire [7:0] t_r44_c28_5;
  wire [7:0] t_r44_c28_6;
  wire [7:0] t_r44_c28_7;
  wire [7:0] t_r44_c28_8;
  wire [7:0] t_r44_c28_9;
  wire [7:0] t_r44_c28_10;
  wire [7:0] t_r44_c28_11;
  wire [7:0] t_r44_c28_12;
  wire [7:0] t_r44_c29_0;
  wire [7:0] t_r44_c29_1;
  wire [7:0] t_r44_c29_2;
  wire [7:0] t_r44_c29_3;
  wire [7:0] t_r44_c29_4;
  wire [7:0] t_r44_c29_5;
  wire [7:0] t_r44_c29_6;
  wire [7:0] t_r44_c29_7;
  wire [7:0] t_r44_c29_8;
  wire [7:0] t_r44_c29_9;
  wire [7:0] t_r44_c29_10;
  wire [7:0] t_r44_c29_11;
  wire [7:0] t_r44_c29_12;
  wire [7:0] t_r44_c30_0;
  wire [7:0] t_r44_c30_1;
  wire [7:0] t_r44_c30_2;
  wire [7:0] t_r44_c30_3;
  wire [7:0] t_r44_c30_4;
  wire [7:0] t_r44_c30_5;
  wire [7:0] t_r44_c30_6;
  wire [7:0] t_r44_c30_7;
  wire [7:0] t_r44_c30_8;
  wire [7:0] t_r44_c30_9;
  wire [7:0] t_r44_c30_10;
  wire [7:0] t_r44_c30_11;
  wire [7:0] t_r44_c30_12;
  wire [7:0] t_r44_c31_0;
  wire [7:0] t_r44_c31_1;
  wire [7:0] t_r44_c31_2;
  wire [7:0] t_r44_c31_3;
  wire [7:0] t_r44_c31_4;
  wire [7:0] t_r44_c31_5;
  wire [7:0] t_r44_c31_6;
  wire [7:0] t_r44_c31_7;
  wire [7:0] t_r44_c31_8;
  wire [7:0] t_r44_c31_9;
  wire [7:0] t_r44_c31_10;
  wire [7:0] t_r44_c31_11;
  wire [7:0] t_r44_c31_12;
  wire [7:0] t_r44_c32_0;
  wire [7:0] t_r44_c32_1;
  wire [7:0] t_r44_c32_2;
  wire [7:0] t_r44_c32_3;
  wire [7:0] t_r44_c32_4;
  wire [7:0] t_r44_c32_5;
  wire [7:0] t_r44_c32_6;
  wire [7:0] t_r44_c32_7;
  wire [7:0] t_r44_c32_8;
  wire [7:0] t_r44_c32_9;
  wire [7:0] t_r44_c32_10;
  wire [7:0] t_r44_c32_11;
  wire [7:0] t_r44_c32_12;
  wire [7:0] t_r44_c33_0;
  wire [7:0] t_r44_c33_1;
  wire [7:0] t_r44_c33_2;
  wire [7:0] t_r44_c33_3;
  wire [7:0] t_r44_c33_4;
  wire [7:0] t_r44_c33_5;
  wire [7:0] t_r44_c33_6;
  wire [7:0] t_r44_c33_7;
  wire [7:0] t_r44_c33_8;
  wire [7:0] t_r44_c33_9;
  wire [7:0] t_r44_c33_10;
  wire [7:0] t_r44_c33_11;
  wire [7:0] t_r44_c33_12;
  wire [7:0] t_r44_c34_0;
  wire [7:0] t_r44_c34_1;
  wire [7:0] t_r44_c34_2;
  wire [7:0] t_r44_c34_3;
  wire [7:0] t_r44_c34_4;
  wire [7:0] t_r44_c34_5;
  wire [7:0] t_r44_c34_6;
  wire [7:0] t_r44_c34_7;
  wire [7:0] t_r44_c34_8;
  wire [7:0] t_r44_c34_9;
  wire [7:0] t_r44_c34_10;
  wire [7:0] t_r44_c34_11;
  wire [7:0] t_r44_c34_12;
  wire [7:0] t_r44_c35_0;
  wire [7:0] t_r44_c35_1;
  wire [7:0] t_r44_c35_2;
  wire [7:0] t_r44_c35_3;
  wire [7:0] t_r44_c35_4;
  wire [7:0] t_r44_c35_5;
  wire [7:0] t_r44_c35_6;
  wire [7:0] t_r44_c35_7;
  wire [7:0] t_r44_c35_8;
  wire [7:0] t_r44_c35_9;
  wire [7:0] t_r44_c35_10;
  wire [7:0] t_r44_c35_11;
  wire [7:0] t_r44_c35_12;
  wire [7:0] t_r44_c36_0;
  wire [7:0] t_r44_c36_1;
  wire [7:0] t_r44_c36_2;
  wire [7:0] t_r44_c36_3;
  wire [7:0] t_r44_c36_4;
  wire [7:0] t_r44_c36_5;
  wire [7:0] t_r44_c36_6;
  wire [7:0] t_r44_c36_7;
  wire [7:0] t_r44_c36_8;
  wire [7:0] t_r44_c36_9;
  wire [7:0] t_r44_c36_10;
  wire [7:0] t_r44_c36_11;
  wire [7:0] t_r44_c36_12;
  wire [7:0] t_r44_c37_0;
  wire [7:0] t_r44_c37_1;
  wire [7:0] t_r44_c37_2;
  wire [7:0] t_r44_c37_3;
  wire [7:0] t_r44_c37_4;
  wire [7:0] t_r44_c37_5;
  wire [7:0] t_r44_c37_6;
  wire [7:0] t_r44_c37_7;
  wire [7:0] t_r44_c37_8;
  wire [7:0] t_r44_c37_9;
  wire [7:0] t_r44_c37_10;
  wire [7:0] t_r44_c37_11;
  wire [7:0] t_r44_c37_12;
  wire [7:0] t_r44_c38_0;
  wire [7:0] t_r44_c38_1;
  wire [7:0] t_r44_c38_2;
  wire [7:0] t_r44_c38_3;
  wire [7:0] t_r44_c38_4;
  wire [7:0] t_r44_c38_5;
  wire [7:0] t_r44_c38_6;
  wire [7:0] t_r44_c38_7;
  wire [7:0] t_r44_c38_8;
  wire [7:0] t_r44_c38_9;
  wire [7:0] t_r44_c38_10;
  wire [7:0] t_r44_c38_11;
  wire [7:0] t_r44_c38_12;
  wire [7:0] t_r44_c39_0;
  wire [7:0] t_r44_c39_1;
  wire [7:0] t_r44_c39_2;
  wire [7:0] t_r44_c39_3;
  wire [7:0] t_r44_c39_4;
  wire [7:0] t_r44_c39_5;
  wire [7:0] t_r44_c39_6;
  wire [7:0] t_r44_c39_7;
  wire [7:0] t_r44_c39_8;
  wire [7:0] t_r44_c39_9;
  wire [7:0] t_r44_c39_10;
  wire [7:0] t_r44_c39_11;
  wire [7:0] t_r44_c39_12;
  wire [7:0] t_r44_c40_0;
  wire [7:0] t_r44_c40_1;
  wire [7:0] t_r44_c40_2;
  wire [7:0] t_r44_c40_3;
  wire [7:0] t_r44_c40_4;
  wire [7:0] t_r44_c40_5;
  wire [7:0] t_r44_c40_6;
  wire [7:0] t_r44_c40_7;
  wire [7:0] t_r44_c40_8;
  wire [7:0] t_r44_c40_9;
  wire [7:0] t_r44_c40_10;
  wire [7:0] t_r44_c40_11;
  wire [7:0] t_r44_c40_12;
  wire [7:0] t_r44_c41_0;
  wire [7:0] t_r44_c41_1;
  wire [7:0] t_r44_c41_2;
  wire [7:0] t_r44_c41_3;
  wire [7:0] t_r44_c41_4;
  wire [7:0] t_r44_c41_5;
  wire [7:0] t_r44_c41_6;
  wire [7:0] t_r44_c41_7;
  wire [7:0] t_r44_c41_8;
  wire [7:0] t_r44_c41_9;
  wire [7:0] t_r44_c41_10;
  wire [7:0] t_r44_c41_11;
  wire [7:0] t_r44_c41_12;
  wire [7:0] t_r44_c42_0;
  wire [7:0] t_r44_c42_1;
  wire [7:0] t_r44_c42_2;
  wire [7:0] t_r44_c42_3;
  wire [7:0] t_r44_c42_4;
  wire [7:0] t_r44_c42_5;
  wire [7:0] t_r44_c42_6;
  wire [7:0] t_r44_c42_7;
  wire [7:0] t_r44_c42_8;
  wire [7:0] t_r44_c42_9;
  wire [7:0] t_r44_c42_10;
  wire [7:0] t_r44_c42_11;
  wire [7:0] t_r44_c42_12;
  wire [7:0] t_r44_c43_0;
  wire [7:0] t_r44_c43_1;
  wire [7:0] t_r44_c43_2;
  wire [7:0] t_r44_c43_3;
  wire [7:0] t_r44_c43_4;
  wire [7:0] t_r44_c43_5;
  wire [7:0] t_r44_c43_6;
  wire [7:0] t_r44_c43_7;
  wire [7:0] t_r44_c43_8;
  wire [7:0] t_r44_c43_9;
  wire [7:0] t_r44_c43_10;
  wire [7:0] t_r44_c43_11;
  wire [7:0] t_r44_c43_12;
  wire [7:0] t_r44_c44_0;
  wire [7:0] t_r44_c44_1;
  wire [7:0] t_r44_c44_2;
  wire [7:0] t_r44_c44_3;
  wire [7:0] t_r44_c44_4;
  wire [7:0] t_r44_c44_5;
  wire [7:0] t_r44_c44_6;
  wire [7:0] t_r44_c44_7;
  wire [7:0] t_r44_c44_8;
  wire [7:0] t_r44_c44_9;
  wire [7:0] t_r44_c44_10;
  wire [7:0] t_r44_c44_11;
  wire [7:0] t_r44_c44_12;
  wire [7:0] t_r44_c45_0;
  wire [7:0] t_r44_c45_1;
  wire [7:0] t_r44_c45_2;
  wire [7:0] t_r44_c45_3;
  wire [7:0] t_r44_c45_4;
  wire [7:0] t_r44_c45_5;
  wire [7:0] t_r44_c45_6;
  wire [7:0] t_r44_c45_7;
  wire [7:0] t_r44_c45_8;
  wire [7:0] t_r44_c45_9;
  wire [7:0] t_r44_c45_10;
  wire [7:0] t_r44_c45_11;
  wire [7:0] t_r44_c45_12;
  wire [7:0] t_r44_c46_0;
  wire [7:0] t_r44_c46_1;
  wire [7:0] t_r44_c46_2;
  wire [7:0] t_r44_c46_3;
  wire [7:0] t_r44_c46_4;
  wire [7:0] t_r44_c46_5;
  wire [7:0] t_r44_c46_6;
  wire [7:0] t_r44_c46_7;
  wire [7:0] t_r44_c46_8;
  wire [7:0] t_r44_c46_9;
  wire [7:0] t_r44_c46_10;
  wire [7:0] t_r44_c46_11;
  wire [7:0] t_r44_c46_12;
  wire [7:0] t_r44_c47_0;
  wire [7:0] t_r44_c47_1;
  wire [7:0] t_r44_c47_2;
  wire [7:0] t_r44_c47_3;
  wire [7:0] t_r44_c47_4;
  wire [7:0] t_r44_c47_5;
  wire [7:0] t_r44_c47_6;
  wire [7:0] t_r44_c47_7;
  wire [7:0] t_r44_c47_8;
  wire [7:0] t_r44_c47_9;
  wire [7:0] t_r44_c47_10;
  wire [7:0] t_r44_c47_11;
  wire [7:0] t_r44_c47_12;
  wire [7:0] t_r44_c48_0;
  wire [7:0] t_r44_c48_1;
  wire [7:0] t_r44_c48_2;
  wire [7:0] t_r44_c48_3;
  wire [7:0] t_r44_c48_4;
  wire [7:0] t_r44_c48_5;
  wire [7:0] t_r44_c48_6;
  wire [7:0] t_r44_c48_7;
  wire [7:0] t_r44_c48_8;
  wire [7:0] t_r44_c48_9;
  wire [7:0] t_r44_c48_10;
  wire [7:0] t_r44_c48_11;
  wire [7:0] t_r44_c48_12;
  wire [7:0] t_r44_c49_0;
  wire [7:0] t_r44_c49_1;
  wire [7:0] t_r44_c49_2;
  wire [7:0] t_r44_c49_3;
  wire [7:0] t_r44_c49_4;
  wire [7:0] t_r44_c49_5;
  wire [7:0] t_r44_c49_6;
  wire [7:0] t_r44_c49_7;
  wire [7:0] t_r44_c49_8;
  wire [7:0] t_r44_c49_9;
  wire [7:0] t_r44_c49_10;
  wire [7:0] t_r44_c49_11;
  wire [7:0] t_r44_c49_12;
  wire [7:0] t_r44_c50_0;
  wire [7:0] t_r44_c50_1;
  wire [7:0] t_r44_c50_2;
  wire [7:0] t_r44_c50_3;
  wire [7:0] t_r44_c50_4;
  wire [7:0] t_r44_c50_5;
  wire [7:0] t_r44_c50_6;
  wire [7:0] t_r44_c50_7;
  wire [7:0] t_r44_c50_8;
  wire [7:0] t_r44_c50_9;
  wire [7:0] t_r44_c50_10;
  wire [7:0] t_r44_c50_11;
  wire [7:0] t_r44_c50_12;
  wire [7:0] t_r44_c51_0;
  wire [7:0] t_r44_c51_1;
  wire [7:0] t_r44_c51_2;
  wire [7:0] t_r44_c51_3;
  wire [7:0] t_r44_c51_4;
  wire [7:0] t_r44_c51_5;
  wire [7:0] t_r44_c51_6;
  wire [7:0] t_r44_c51_7;
  wire [7:0] t_r44_c51_8;
  wire [7:0] t_r44_c51_9;
  wire [7:0] t_r44_c51_10;
  wire [7:0] t_r44_c51_11;
  wire [7:0] t_r44_c51_12;
  wire [7:0] t_r44_c52_0;
  wire [7:0] t_r44_c52_1;
  wire [7:0] t_r44_c52_2;
  wire [7:0] t_r44_c52_3;
  wire [7:0] t_r44_c52_4;
  wire [7:0] t_r44_c52_5;
  wire [7:0] t_r44_c52_6;
  wire [7:0] t_r44_c52_7;
  wire [7:0] t_r44_c52_8;
  wire [7:0] t_r44_c52_9;
  wire [7:0] t_r44_c52_10;
  wire [7:0] t_r44_c52_11;
  wire [7:0] t_r44_c52_12;
  wire [7:0] t_r44_c53_0;
  wire [7:0] t_r44_c53_1;
  wire [7:0] t_r44_c53_2;
  wire [7:0] t_r44_c53_3;
  wire [7:0] t_r44_c53_4;
  wire [7:0] t_r44_c53_5;
  wire [7:0] t_r44_c53_6;
  wire [7:0] t_r44_c53_7;
  wire [7:0] t_r44_c53_8;
  wire [7:0] t_r44_c53_9;
  wire [7:0] t_r44_c53_10;
  wire [7:0] t_r44_c53_11;
  wire [7:0] t_r44_c53_12;
  wire [7:0] t_r44_c54_0;
  wire [7:0] t_r44_c54_1;
  wire [7:0] t_r44_c54_2;
  wire [7:0] t_r44_c54_3;
  wire [7:0] t_r44_c54_4;
  wire [7:0] t_r44_c54_5;
  wire [7:0] t_r44_c54_6;
  wire [7:0] t_r44_c54_7;
  wire [7:0] t_r44_c54_8;
  wire [7:0] t_r44_c54_9;
  wire [7:0] t_r44_c54_10;
  wire [7:0] t_r44_c54_11;
  wire [7:0] t_r44_c54_12;
  wire [7:0] t_r44_c55_0;
  wire [7:0] t_r44_c55_1;
  wire [7:0] t_r44_c55_2;
  wire [7:0] t_r44_c55_3;
  wire [7:0] t_r44_c55_4;
  wire [7:0] t_r44_c55_5;
  wire [7:0] t_r44_c55_6;
  wire [7:0] t_r44_c55_7;
  wire [7:0] t_r44_c55_8;
  wire [7:0] t_r44_c55_9;
  wire [7:0] t_r44_c55_10;
  wire [7:0] t_r44_c55_11;
  wire [7:0] t_r44_c55_12;
  wire [7:0] t_r44_c56_0;
  wire [7:0] t_r44_c56_1;
  wire [7:0] t_r44_c56_2;
  wire [7:0] t_r44_c56_3;
  wire [7:0] t_r44_c56_4;
  wire [7:0] t_r44_c56_5;
  wire [7:0] t_r44_c56_6;
  wire [7:0] t_r44_c56_7;
  wire [7:0] t_r44_c56_8;
  wire [7:0] t_r44_c56_9;
  wire [7:0] t_r44_c56_10;
  wire [7:0] t_r44_c56_11;
  wire [7:0] t_r44_c56_12;
  wire [7:0] t_r44_c57_0;
  wire [7:0] t_r44_c57_1;
  wire [7:0] t_r44_c57_2;
  wire [7:0] t_r44_c57_3;
  wire [7:0] t_r44_c57_4;
  wire [7:0] t_r44_c57_5;
  wire [7:0] t_r44_c57_6;
  wire [7:0] t_r44_c57_7;
  wire [7:0] t_r44_c57_8;
  wire [7:0] t_r44_c57_9;
  wire [7:0] t_r44_c57_10;
  wire [7:0] t_r44_c57_11;
  wire [7:0] t_r44_c57_12;
  wire [7:0] t_r44_c58_0;
  wire [7:0] t_r44_c58_1;
  wire [7:0] t_r44_c58_2;
  wire [7:0] t_r44_c58_3;
  wire [7:0] t_r44_c58_4;
  wire [7:0] t_r44_c58_5;
  wire [7:0] t_r44_c58_6;
  wire [7:0] t_r44_c58_7;
  wire [7:0] t_r44_c58_8;
  wire [7:0] t_r44_c58_9;
  wire [7:0] t_r44_c58_10;
  wire [7:0] t_r44_c58_11;
  wire [7:0] t_r44_c58_12;
  wire [7:0] t_r44_c59_0;
  wire [7:0] t_r44_c59_1;
  wire [7:0] t_r44_c59_2;
  wire [7:0] t_r44_c59_3;
  wire [7:0] t_r44_c59_4;
  wire [7:0] t_r44_c59_5;
  wire [7:0] t_r44_c59_6;
  wire [7:0] t_r44_c59_7;
  wire [7:0] t_r44_c59_8;
  wire [7:0] t_r44_c59_9;
  wire [7:0] t_r44_c59_10;
  wire [7:0] t_r44_c59_11;
  wire [7:0] t_r44_c59_12;
  wire [7:0] t_r44_c60_0;
  wire [7:0] t_r44_c60_1;
  wire [7:0] t_r44_c60_2;
  wire [7:0] t_r44_c60_3;
  wire [7:0] t_r44_c60_4;
  wire [7:0] t_r44_c60_5;
  wire [7:0] t_r44_c60_6;
  wire [7:0] t_r44_c60_7;
  wire [7:0] t_r44_c60_8;
  wire [7:0] t_r44_c60_9;
  wire [7:0] t_r44_c60_10;
  wire [7:0] t_r44_c60_11;
  wire [7:0] t_r44_c60_12;
  wire [7:0] t_r44_c61_0;
  wire [7:0] t_r44_c61_1;
  wire [7:0] t_r44_c61_2;
  wire [7:0] t_r44_c61_3;
  wire [7:0] t_r44_c61_4;
  wire [7:0] t_r44_c61_5;
  wire [7:0] t_r44_c61_6;
  wire [7:0] t_r44_c61_7;
  wire [7:0] t_r44_c61_8;
  wire [7:0] t_r44_c61_9;
  wire [7:0] t_r44_c61_10;
  wire [7:0] t_r44_c61_11;
  wire [7:0] t_r44_c61_12;
  wire [7:0] t_r44_c62_0;
  wire [7:0] t_r44_c62_1;
  wire [7:0] t_r44_c62_2;
  wire [7:0] t_r44_c62_3;
  wire [7:0] t_r44_c62_4;
  wire [7:0] t_r44_c62_5;
  wire [7:0] t_r44_c62_6;
  wire [7:0] t_r44_c62_7;
  wire [7:0] t_r44_c62_8;
  wire [7:0] t_r44_c62_9;
  wire [7:0] t_r44_c62_10;
  wire [7:0] t_r44_c62_11;
  wire [7:0] t_r44_c62_12;
  wire [7:0] t_r44_c63_0;
  wire [7:0] t_r44_c63_1;
  wire [7:0] t_r44_c63_2;
  wire [7:0] t_r44_c63_3;
  wire [7:0] t_r44_c63_4;
  wire [7:0] t_r44_c63_5;
  wire [7:0] t_r44_c63_6;
  wire [7:0] t_r44_c63_7;
  wire [7:0] t_r44_c63_8;
  wire [7:0] t_r44_c63_9;
  wire [7:0] t_r44_c63_10;
  wire [7:0] t_r44_c63_11;
  wire [7:0] t_r44_c63_12;
  wire [7:0] t_r44_c64_0;
  wire [7:0] t_r44_c64_1;
  wire [7:0] t_r44_c64_2;
  wire [7:0] t_r44_c64_3;
  wire [7:0] t_r44_c64_4;
  wire [7:0] t_r44_c64_5;
  wire [7:0] t_r44_c64_6;
  wire [7:0] t_r44_c64_7;
  wire [7:0] t_r44_c64_8;
  wire [7:0] t_r44_c64_9;
  wire [7:0] t_r44_c64_10;
  wire [7:0] t_r44_c64_11;
  wire [7:0] t_r44_c64_12;
  wire [7:0] t_r44_c65_0;
  wire [7:0] t_r44_c65_1;
  wire [7:0] t_r44_c65_2;
  wire [7:0] t_r44_c65_3;
  wire [7:0] t_r44_c65_4;
  wire [7:0] t_r44_c65_5;
  wire [7:0] t_r44_c65_6;
  wire [7:0] t_r44_c65_7;
  wire [7:0] t_r44_c65_8;
  wire [7:0] t_r44_c65_9;
  wire [7:0] t_r44_c65_10;
  wire [7:0] t_r44_c65_11;
  wire [7:0] t_r44_c65_12;

  assign t_r1_c1_0 = p_0_1 << 1;
  assign t_r1_c1_1 = p_1_0 << 1;
  assign t_r1_c1_2 = p_1_1 << 2;
  assign t_r1_c1_3 = p_1_2 << 1;
  assign t_r1_c1_4 = p_2_1 << 1;
  assign t_r1_c1_5 = t_r1_c1_0 + p_0_0;
  assign t_r1_c1_6 = t_r1_c1_1 + p_0_2;
  assign t_r1_c1_7 = t_r1_c1_2 + t_r1_c1_3;
  assign t_r1_c1_8 = t_r1_c1_4 + p_2_0;
  assign t_r1_c1_9 = t_r1_c1_5 + t_r1_c1_6;
  assign t_r1_c1_10 = t_r1_c1_7 + t_r1_c1_8;
  assign t_r1_c1_11 = t_r1_c1_9 + t_r1_c1_10;
  assign t_r1_c1_12 = t_r1_c1_11 + p_2_2;
  assign out_1_1 = t_r1_c1_12 >> 4;

  assign t_r1_c2_0 = p_0_2 << 1;
  assign t_r1_c2_1 = p_1_1 << 1;
  assign t_r1_c2_2 = p_1_2 << 2;
  assign t_r1_c2_3 = p_1_3 << 1;
  assign t_r1_c2_4 = p_2_2 << 1;
  assign t_r1_c2_5 = t_r1_c2_0 + p_0_1;
  assign t_r1_c2_6 = t_r1_c2_1 + p_0_3;
  assign t_r1_c2_7 = t_r1_c2_2 + t_r1_c2_3;
  assign t_r1_c2_8 = t_r1_c2_4 + p_2_1;
  assign t_r1_c2_9 = t_r1_c2_5 + t_r1_c2_6;
  assign t_r1_c2_10 = t_r1_c2_7 + t_r1_c2_8;
  assign t_r1_c2_11 = t_r1_c2_9 + t_r1_c2_10;
  assign t_r1_c2_12 = t_r1_c2_11 + p_2_3;
  assign out_1_2 = t_r1_c2_12 >> 4;

  assign t_r1_c3_0 = p_0_3 << 1;
  assign t_r1_c3_1 = p_1_2 << 1;
  assign t_r1_c3_2 = p_1_3 << 2;
  assign t_r1_c3_3 = p_1_4 << 1;
  assign t_r1_c3_4 = p_2_3 << 1;
  assign t_r1_c3_5 = t_r1_c3_0 + p_0_2;
  assign t_r1_c3_6 = t_r1_c3_1 + p_0_4;
  assign t_r1_c3_7 = t_r1_c3_2 + t_r1_c3_3;
  assign t_r1_c3_8 = t_r1_c3_4 + p_2_2;
  assign t_r1_c3_9 = t_r1_c3_5 + t_r1_c3_6;
  assign t_r1_c3_10 = t_r1_c3_7 + t_r1_c3_8;
  assign t_r1_c3_11 = t_r1_c3_9 + t_r1_c3_10;
  assign t_r1_c3_12 = t_r1_c3_11 + p_2_4;
  assign out_1_3 = t_r1_c3_12 >> 4;

  assign t_r1_c4_0 = p_0_4 << 1;
  assign t_r1_c4_1 = p_1_3 << 1;
  assign t_r1_c4_2 = p_1_4 << 2;
  assign t_r1_c4_3 = p_1_5 << 1;
  assign t_r1_c4_4 = p_2_4 << 1;
  assign t_r1_c4_5 = t_r1_c4_0 + p_0_3;
  assign t_r1_c4_6 = t_r1_c4_1 + p_0_5;
  assign t_r1_c4_7 = t_r1_c4_2 + t_r1_c4_3;
  assign t_r1_c4_8 = t_r1_c4_4 + p_2_3;
  assign t_r1_c4_9 = t_r1_c4_5 + t_r1_c4_6;
  assign t_r1_c4_10 = t_r1_c4_7 + t_r1_c4_8;
  assign t_r1_c4_11 = t_r1_c4_9 + t_r1_c4_10;
  assign t_r1_c4_12 = t_r1_c4_11 + p_2_5;
  assign out_1_4 = t_r1_c4_12 >> 4;

  assign t_r1_c5_0 = p_0_5 << 1;
  assign t_r1_c5_1 = p_1_4 << 1;
  assign t_r1_c5_2 = p_1_5 << 2;
  assign t_r1_c5_3 = p_1_6 << 1;
  assign t_r1_c5_4 = p_2_5 << 1;
  assign t_r1_c5_5 = t_r1_c5_0 + p_0_4;
  assign t_r1_c5_6 = t_r1_c5_1 + p_0_6;
  assign t_r1_c5_7 = t_r1_c5_2 + t_r1_c5_3;
  assign t_r1_c5_8 = t_r1_c5_4 + p_2_4;
  assign t_r1_c5_9 = t_r1_c5_5 + t_r1_c5_6;
  assign t_r1_c5_10 = t_r1_c5_7 + t_r1_c5_8;
  assign t_r1_c5_11 = t_r1_c5_9 + t_r1_c5_10;
  assign t_r1_c5_12 = t_r1_c5_11 + p_2_6;
  assign out_1_5 = t_r1_c5_12 >> 4;

  assign t_r1_c6_0 = p_0_6 << 1;
  assign t_r1_c6_1 = p_1_5 << 1;
  assign t_r1_c6_2 = p_1_6 << 2;
  assign t_r1_c6_3 = p_1_7 << 1;
  assign t_r1_c6_4 = p_2_6 << 1;
  assign t_r1_c6_5 = t_r1_c6_0 + p_0_5;
  assign t_r1_c6_6 = t_r1_c6_1 + p_0_7;
  assign t_r1_c6_7 = t_r1_c6_2 + t_r1_c6_3;
  assign t_r1_c6_8 = t_r1_c6_4 + p_2_5;
  assign t_r1_c6_9 = t_r1_c6_5 + t_r1_c6_6;
  assign t_r1_c6_10 = t_r1_c6_7 + t_r1_c6_8;
  assign t_r1_c6_11 = t_r1_c6_9 + t_r1_c6_10;
  assign t_r1_c6_12 = t_r1_c6_11 + p_2_7;
  assign out_1_6 = t_r1_c6_12 >> 4;

  assign t_r1_c7_0 = p_0_7 << 1;
  assign t_r1_c7_1 = p_1_6 << 1;
  assign t_r1_c7_2 = p_1_7 << 2;
  assign t_r1_c7_3 = p_1_8 << 1;
  assign t_r1_c7_4 = p_2_7 << 1;
  assign t_r1_c7_5 = t_r1_c7_0 + p_0_6;
  assign t_r1_c7_6 = t_r1_c7_1 + p_0_8;
  assign t_r1_c7_7 = t_r1_c7_2 + t_r1_c7_3;
  assign t_r1_c7_8 = t_r1_c7_4 + p_2_6;
  assign t_r1_c7_9 = t_r1_c7_5 + t_r1_c7_6;
  assign t_r1_c7_10 = t_r1_c7_7 + t_r1_c7_8;
  assign t_r1_c7_11 = t_r1_c7_9 + t_r1_c7_10;
  assign t_r1_c7_12 = t_r1_c7_11 + p_2_8;
  assign out_1_7 = t_r1_c7_12 >> 4;

  assign t_r1_c8_0 = p_0_8 << 1;
  assign t_r1_c8_1 = p_1_7 << 1;
  assign t_r1_c8_2 = p_1_8 << 2;
  assign t_r1_c8_3 = p_1_9 << 1;
  assign t_r1_c8_4 = p_2_8 << 1;
  assign t_r1_c8_5 = t_r1_c8_0 + p_0_7;
  assign t_r1_c8_6 = t_r1_c8_1 + p_0_9;
  assign t_r1_c8_7 = t_r1_c8_2 + t_r1_c8_3;
  assign t_r1_c8_8 = t_r1_c8_4 + p_2_7;
  assign t_r1_c8_9 = t_r1_c8_5 + t_r1_c8_6;
  assign t_r1_c8_10 = t_r1_c8_7 + t_r1_c8_8;
  assign t_r1_c8_11 = t_r1_c8_9 + t_r1_c8_10;
  assign t_r1_c8_12 = t_r1_c8_11 + p_2_9;
  assign out_1_8 = t_r1_c8_12 >> 4;

  assign t_r1_c9_0 = p_0_9 << 1;
  assign t_r1_c9_1 = p_1_8 << 1;
  assign t_r1_c9_2 = p_1_9 << 2;
  assign t_r1_c9_3 = p_1_10 << 1;
  assign t_r1_c9_4 = p_2_9 << 1;
  assign t_r1_c9_5 = t_r1_c9_0 + p_0_8;
  assign t_r1_c9_6 = t_r1_c9_1 + p_0_10;
  assign t_r1_c9_7 = t_r1_c9_2 + t_r1_c9_3;
  assign t_r1_c9_8 = t_r1_c9_4 + p_2_8;
  assign t_r1_c9_9 = t_r1_c9_5 + t_r1_c9_6;
  assign t_r1_c9_10 = t_r1_c9_7 + t_r1_c9_8;
  assign t_r1_c9_11 = t_r1_c9_9 + t_r1_c9_10;
  assign t_r1_c9_12 = t_r1_c9_11 + p_2_10;
  assign out_1_9 = t_r1_c9_12 >> 4;

  assign t_r1_c10_0 = p_0_10 << 1;
  assign t_r1_c10_1 = p_1_9 << 1;
  assign t_r1_c10_2 = p_1_10 << 2;
  assign t_r1_c10_3 = p_1_11 << 1;
  assign t_r1_c10_4 = p_2_10 << 1;
  assign t_r1_c10_5 = t_r1_c10_0 + p_0_9;
  assign t_r1_c10_6 = t_r1_c10_1 + p_0_11;
  assign t_r1_c10_7 = t_r1_c10_2 + t_r1_c10_3;
  assign t_r1_c10_8 = t_r1_c10_4 + p_2_9;
  assign t_r1_c10_9 = t_r1_c10_5 + t_r1_c10_6;
  assign t_r1_c10_10 = t_r1_c10_7 + t_r1_c10_8;
  assign t_r1_c10_11 = t_r1_c10_9 + t_r1_c10_10;
  assign t_r1_c10_12 = t_r1_c10_11 + p_2_11;
  assign out_1_10 = t_r1_c10_12 >> 4;

  assign t_r1_c11_0 = p_0_11 << 1;
  assign t_r1_c11_1 = p_1_10 << 1;
  assign t_r1_c11_2 = p_1_11 << 2;
  assign t_r1_c11_3 = p_1_12 << 1;
  assign t_r1_c11_4 = p_2_11 << 1;
  assign t_r1_c11_5 = t_r1_c11_0 + p_0_10;
  assign t_r1_c11_6 = t_r1_c11_1 + p_0_12;
  assign t_r1_c11_7 = t_r1_c11_2 + t_r1_c11_3;
  assign t_r1_c11_8 = t_r1_c11_4 + p_2_10;
  assign t_r1_c11_9 = t_r1_c11_5 + t_r1_c11_6;
  assign t_r1_c11_10 = t_r1_c11_7 + t_r1_c11_8;
  assign t_r1_c11_11 = t_r1_c11_9 + t_r1_c11_10;
  assign t_r1_c11_12 = t_r1_c11_11 + p_2_12;
  assign out_1_11 = t_r1_c11_12 >> 4;

  assign t_r1_c12_0 = p_0_12 << 1;
  assign t_r1_c12_1 = p_1_11 << 1;
  assign t_r1_c12_2 = p_1_12 << 2;
  assign t_r1_c12_3 = p_1_13 << 1;
  assign t_r1_c12_4 = p_2_12 << 1;
  assign t_r1_c12_5 = t_r1_c12_0 + p_0_11;
  assign t_r1_c12_6 = t_r1_c12_1 + p_0_13;
  assign t_r1_c12_7 = t_r1_c12_2 + t_r1_c12_3;
  assign t_r1_c12_8 = t_r1_c12_4 + p_2_11;
  assign t_r1_c12_9 = t_r1_c12_5 + t_r1_c12_6;
  assign t_r1_c12_10 = t_r1_c12_7 + t_r1_c12_8;
  assign t_r1_c12_11 = t_r1_c12_9 + t_r1_c12_10;
  assign t_r1_c12_12 = t_r1_c12_11 + p_2_13;
  assign out_1_12 = t_r1_c12_12 >> 4;

  assign t_r1_c13_0 = p_0_13 << 1;
  assign t_r1_c13_1 = p_1_12 << 1;
  assign t_r1_c13_2 = p_1_13 << 2;
  assign t_r1_c13_3 = p_1_14 << 1;
  assign t_r1_c13_4 = p_2_13 << 1;
  assign t_r1_c13_5 = t_r1_c13_0 + p_0_12;
  assign t_r1_c13_6 = t_r1_c13_1 + p_0_14;
  assign t_r1_c13_7 = t_r1_c13_2 + t_r1_c13_3;
  assign t_r1_c13_8 = t_r1_c13_4 + p_2_12;
  assign t_r1_c13_9 = t_r1_c13_5 + t_r1_c13_6;
  assign t_r1_c13_10 = t_r1_c13_7 + t_r1_c13_8;
  assign t_r1_c13_11 = t_r1_c13_9 + t_r1_c13_10;
  assign t_r1_c13_12 = t_r1_c13_11 + p_2_14;
  assign out_1_13 = t_r1_c13_12 >> 4;

  assign t_r1_c14_0 = p_0_14 << 1;
  assign t_r1_c14_1 = p_1_13 << 1;
  assign t_r1_c14_2 = p_1_14 << 2;
  assign t_r1_c14_3 = p_1_15 << 1;
  assign t_r1_c14_4 = p_2_14 << 1;
  assign t_r1_c14_5 = t_r1_c14_0 + p_0_13;
  assign t_r1_c14_6 = t_r1_c14_1 + p_0_15;
  assign t_r1_c14_7 = t_r1_c14_2 + t_r1_c14_3;
  assign t_r1_c14_8 = t_r1_c14_4 + p_2_13;
  assign t_r1_c14_9 = t_r1_c14_5 + t_r1_c14_6;
  assign t_r1_c14_10 = t_r1_c14_7 + t_r1_c14_8;
  assign t_r1_c14_11 = t_r1_c14_9 + t_r1_c14_10;
  assign t_r1_c14_12 = t_r1_c14_11 + p_2_15;
  assign out_1_14 = t_r1_c14_12 >> 4;

  assign t_r1_c15_0 = p_0_15 << 1;
  assign t_r1_c15_1 = p_1_14 << 1;
  assign t_r1_c15_2 = p_1_15 << 2;
  assign t_r1_c15_3 = p_1_16 << 1;
  assign t_r1_c15_4 = p_2_15 << 1;
  assign t_r1_c15_5 = t_r1_c15_0 + p_0_14;
  assign t_r1_c15_6 = t_r1_c15_1 + p_0_16;
  assign t_r1_c15_7 = t_r1_c15_2 + t_r1_c15_3;
  assign t_r1_c15_8 = t_r1_c15_4 + p_2_14;
  assign t_r1_c15_9 = t_r1_c15_5 + t_r1_c15_6;
  assign t_r1_c15_10 = t_r1_c15_7 + t_r1_c15_8;
  assign t_r1_c15_11 = t_r1_c15_9 + t_r1_c15_10;
  assign t_r1_c15_12 = t_r1_c15_11 + p_2_16;
  assign out_1_15 = t_r1_c15_12 >> 4;

  assign t_r1_c16_0 = p_0_16 << 1;
  assign t_r1_c16_1 = p_1_15 << 1;
  assign t_r1_c16_2 = p_1_16 << 2;
  assign t_r1_c16_3 = p_1_17 << 1;
  assign t_r1_c16_4 = p_2_16 << 1;
  assign t_r1_c16_5 = t_r1_c16_0 + p_0_15;
  assign t_r1_c16_6 = t_r1_c16_1 + p_0_17;
  assign t_r1_c16_7 = t_r1_c16_2 + t_r1_c16_3;
  assign t_r1_c16_8 = t_r1_c16_4 + p_2_15;
  assign t_r1_c16_9 = t_r1_c16_5 + t_r1_c16_6;
  assign t_r1_c16_10 = t_r1_c16_7 + t_r1_c16_8;
  assign t_r1_c16_11 = t_r1_c16_9 + t_r1_c16_10;
  assign t_r1_c16_12 = t_r1_c16_11 + p_2_17;
  assign out_1_16 = t_r1_c16_12 >> 4;

  assign t_r1_c17_0 = p_0_17 << 1;
  assign t_r1_c17_1 = p_1_16 << 1;
  assign t_r1_c17_2 = p_1_17 << 2;
  assign t_r1_c17_3 = p_1_18 << 1;
  assign t_r1_c17_4 = p_2_17 << 1;
  assign t_r1_c17_5 = t_r1_c17_0 + p_0_16;
  assign t_r1_c17_6 = t_r1_c17_1 + p_0_18;
  assign t_r1_c17_7 = t_r1_c17_2 + t_r1_c17_3;
  assign t_r1_c17_8 = t_r1_c17_4 + p_2_16;
  assign t_r1_c17_9 = t_r1_c17_5 + t_r1_c17_6;
  assign t_r1_c17_10 = t_r1_c17_7 + t_r1_c17_8;
  assign t_r1_c17_11 = t_r1_c17_9 + t_r1_c17_10;
  assign t_r1_c17_12 = t_r1_c17_11 + p_2_18;
  assign out_1_17 = t_r1_c17_12 >> 4;

  assign t_r1_c18_0 = p_0_18 << 1;
  assign t_r1_c18_1 = p_1_17 << 1;
  assign t_r1_c18_2 = p_1_18 << 2;
  assign t_r1_c18_3 = p_1_19 << 1;
  assign t_r1_c18_4 = p_2_18 << 1;
  assign t_r1_c18_5 = t_r1_c18_0 + p_0_17;
  assign t_r1_c18_6 = t_r1_c18_1 + p_0_19;
  assign t_r1_c18_7 = t_r1_c18_2 + t_r1_c18_3;
  assign t_r1_c18_8 = t_r1_c18_4 + p_2_17;
  assign t_r1_c18_9 = t_r1_c18_5 + t_r1_c18_6;
  assign t_r1_c18_10 = t_r1_c18_7 + t_r1_c18_8;
  assign t_r1_c18_11 = t_r1_c18_9 + t_r1_c18_10;
  assign t_r1_c18_12 = t_r1_c18_11 + p_2_19;
  assign out_1_18 = t_r1_c18_12 >> 4;

  assign t_r1_c19_0 = p_0_19 << 1;
  assign t_r1_c19_1 = p_1_18 << 1;
  assign t_r1_c19_2 = p_1_19 << 2;
  assign t_r1_c19_3 = p_1_20 << 1;
  assign t_r1_c19_4 = p_2_19 << 1;
  assign t_r1_c19_5 = t_r1_c19_0 + p_0_18;
  assign t_r1_c19_6 = t_r1_c19_1 + p_0_20;
  assign t_r1_c19_7 = t_r1_c19_2 + t_r1_c19_3;
  assign t_r1_c19_8 = t_r1_c19_4 + p_2_18;
  assign t_r1_c19_9 = t_r1_c19_5 + t_r1_c19_6;
  assign t_r1_c19_10 = t_r1_c19_7 + t_r1_c19_8;
  assign t_r1_c19_11 = t_r1_c19_9 + t_r1_c19_10;
  assign t_r1_c19_12 = t_r1_c19_11 + p_2_20;
  assign out_1_19 = t_r1_c19_12 >> 4;

  assign t_r1_c20_0 = p_0_20 << 1;
  assign t_r1_c20_1 = p_1_19 << 1;
  assign t_r1_c20_2 = p_1_20 << 2;
  assign t_r1_c20_3 = p_1_21 << 1;
  assign t_r1_c20_4 = p_2_20 << 1;
  assign t_r1_c20_5 = t_r1_c20_0 + p_0_19;
  assign t_r1_c20_6 = t_r1_c20_1 + p_0_21;
  assign t_r1_c20_7 = t_r1_c20_2 + t_r1_c20_3;
  assign t_r1_c20_8 = t_r1_c20_4 + p_2_19;
  assign t_r1_c20_9 = t_r1_c20_5 + t_r1_c20_6;
  assign t_r1_c20_10 = t_r1_c20_7 + t_r1_c20_8;
  assign t_r1_c20_11 = t_r1_c20_9 + t_r1_c20_10;
  assign t_r1_c20_12 = t_r1_c20_11 + p_2_21;
  assign out_1_20 = t_r1_c20_12 >> 4;

  assign t_r1_c21_0 = p_0_21 << 1;
  assign t_r1_c21_1 = p_1_20 << 1;
  assign t_r1_c21_2 = p_1_21 << 2;
  assign t_r1_c21_3 = p_1_22 << 1;
  assign t_r1_c21_4 = p_2_21 << 1;
  assign t_r1_c21_5 = t_r1_c21_0 + p_0_20;
  assign t_r1_c21_6 = t_r1_c21_1 + p_0_22;
  assign t_r1_c21_7 = t_r1_c21_2 + t_r1_c21_3;
  assign t_r1_c21_8 = t_r1_c21_4 + p_2_20;
  assign t_r1_c21_9 = t_r1_c21_5 + t_r1_c21_6;
  assign t_r1_c21_10 = t_r1_c21_7 + t_r1_c21_8;
  assign t_r1_c21_11 = t_r1_c21_9 + t_r1_c21_10;
  assign t_r1_c21_12 = t_r1_c21_11 + p_2_22;
  assign out_1_21 = t_r1_c21_12 >> 4;

  assign t_r1_c22_0 = p_0_22 << 1;
  assign t_r1_c22_1 = p_1_21 << 1;
  assign t_r1_c22_2 = p_1_22 << 2;
  assign t_r1_c22_3 = p_1_23 << 1;
  assign t_r1_c22_4 = p_2_22 << 1;
  assign t_r1_c22_5 = t_r1_c22_0 + p_0_21;
  assign t_r1_c22_6 = t_r1_c22_1 + p_0_23;
  assign t_r1_c22_7 = t_r1_c22_2 + t_r1_c22_3;
  assign t_r1_c22_8 = t_r1_c22_4 + p_2_21;
  assign t_r1_c22_9 = t_r1_c22_5 + t_r1_c22_6;
  assign t_r1_c22_10 = t_r1_c22_7 + t_r1_c22_8;
  assign t_r1_c22_11 = t_r1_c22_9 + t_r1_c22_10;
  assign t_r1_c22_12 = t_r1_c22_11 + p_2_23;
  assign out_1_22 = t_r1_c22_12 >> 4;

  assign t_r1_c23_0 = p_0_23 << 1;
  assign t_r1_c23_1 = p_1_22 << 1;
  assign t_r1_c23_2 = p_1_23 << 2;
  assign t_r1_c23_3 = p_1_24 << 1;
  assign t_r1_c23_4 = p_2_23 << 1;
  assign t_r1_c23_5 = t_r1_c23_0 + p_0_22;
  assign t_r1_c23_6 = t_r1_c23_1 + p_0_24;
  assign t_r1_c23_7 = t_r1_c23_2 + t_r1_c23_3;
  assign t_r1_c23_8 = t_r1_c23_4 + p_2_22;
  assign t_r1_c23_9 = t_r1_c23_5 + t_r1_c23_6;
  assign t_r1_c23_10 = t_r1_c23_7 + t_r1_c23_8;
  assign t_r1_c23_11 = t_r1_c23_9 + t_r1_c23_10;
  assign t_r1_c23_12 = t_r1_c23_11 + p_2_24;
  assign out_1_23 = t_r1_c23_12 >> 4;

  assign t_r1_c24_0 = p_0_24 << 1;
  assign t_r1_c24_1 = p_1_23 << 1;
  assign t_r1_c24_2 = p_1_24 << 2;
  assign t_r1_c24_3 = p_1_25 << 1;
  assign t_r1_c24_4 = p_2_24 << 1;
  assign t_r1_c24_5 = t_r1_c24_0 + p_0_23;
  assign t_r1_c24_6 = t_r1_c24_1 + p_0_25;
  assign t_r1_c24_7 = t_r1_c24_2 + t_r1_c24_3;
  assign t_r1_c24_8 = t_r1_c24_4 + p_2_23;
  assign t_r1_c24_9 = t_r1_c24_5 + t_r1_c24_6;
  assign t_r1_c24_10 = t_r1_c24_7 + t_r1_c24_8;
  assign t_r1_c24_11 = t_r1_c24_9 + t_r1_c24_10;
  assign t_r1_c24_12 = t_r1_c24_11 + p_2_25;
  assign out_1_24 = t_r1_c24_12 >> 4;

  assign t_r1_c25_0 = p_0_25 << 1;
  assign t_r1_c25_1 = p_1_24 << 1;
  assign t_r1_c25_2 = p_1_25 << 2;
  assign t_r1_c25_3 = p_1_26 << 1;
  assign t_r1_c25_4 = p_2_25 << 1;
  assign t_r1_c25_5 = t_r1_c25_0 + p_0_24;
  assign t_r1_c25_6 = t_r1_c25_1 + p_0_26;
  assign t_r1_c25_7 = t_r1_c25_2 + t_r1_c25_3;
  assign t_r1_c25_8 = t_r1_c25_4 + p_2_24;
  assign t_r1_c25_9 = t_r1_c25_5 + t_r1_c25_6;
  assign t_r1_c25_10 = t_r1_c25_7 + t_r1_c25_8;
  assign t_r1_c25_11 = t_r1_c25_9 + t_r1_c25_10;
  assign t_r1_c25_12 = t_r1_c25_11 + p_2_26;
  assign out_1_25 = t_r1_c25_12 >> 4;

  assign t_r1_c26_0 = p_0_26 << 1;
  assign t_r1_c26_1 = p_1_25 << 1;
  assign t_r1_c26_2 = p_1_26 << 2;
  assign t_r1_c26_3 = p_1_27 << 1;
  assign t_r1_c26_4 = p_2_26 << 1;
  assign t_r1_c26_5 = t_r1_c26_0 + p_0_25;
  assign t_r1_c26_6 = t_r1_c26_1 + p_0_27;
  assign t_r1_c26_7 = t_r1_c26_2 + t_r1_c26_3;
  assign t_r1_c26_8 = t_r1_c26_4 + p_2_25;
  assign t_r1_c26_9 = t_r1_c26_5 + t_r1_c26_6;
  assign t_r1_c26_10 = t_r1_c26_7 + t_r1_c26_8;
  assign t_r1_c26_11 = t_r1_c26_9 + t_r1_c26_10;
  assign t_r1_c26_12 = t_r1_c26_11 + p_2_27;
  assign out_1_26 = t_r1_c26_12 >> 4;

  assign t_r1_c27_0 = p_0_27 << 1;
  assign t_r1_c27_1 = p_1_26 << 1;
  assign t_r1_c27_2 = p_1_27 << 2;
  assign t_r1_c27_3 = p_1_28 << 1;
  assign t_r1_c27_4 = p_2_27 << 1;
  assign t_r1_c27_5 = t_r1_c27_0 + p_0_26;
  assign t_r1_c27_6 = t_r1_c27_1 + p_0_28;
  assign t_r1_c27_7 = t_r1_c27_2 + t_r1_c27_3;
  assign t_r1_c27_8 = t_r1_c27_4 + p_2_26;
  assign t_r1_c27_9 = t_r1_c27_5 + t_r1_c27_6;
  assign t_r1_c27_10 = t_r1_c27_7 + t_r1_c27_8;
  assign t_r1_c27_11 = t_r1_c27_9 + t_r1_c27_10;
  assign t_r1_c27_12 = t_r1_c27_11 + p_2_28;
  assign out_1_27 = t_r1_c27_12 >> 4;

  assign t_r1_c28_0 = p_0_28 << 1;
  assign t_r1_c28_1 = p_1_27 << 1;
  assign t_r1_c28_2 = p_1_28 << 2;
  assign t_r1_c28_3 = p_1_29 << 1;
  assign t_r1_c28_4 = p_2_28 << 1;
  assign t_r1_c28_5 = t_r1_c28_0 + p_0_27;
  assign t_r1_c28_6 = t_r1_c28_1 + p_0_29;
  assign t_r1_c28_7 = t_r1_c28_2 + t_r1_c28_3;
  assign t_r1_c28_8 = t_r1_c28_4 + p_2_27;
  assign t_r1_c28_9 = t_r1_c28_5 + t_r1_c28_6;
  assign t_r1_c28_10 = t_r1_c28_7 + t_r1_c28_8;
  assign t_r1_c28_11 = t_r1_c28_9 + t_r1_c28_10;
  assign t_r1_c28_12 = t_r1_c28_11 + p_2_29;
  assign out_1_28 = t_r1_c28_12 >> 4;

  assign t_r1_c29_0 = p_0_29 << 1;
  assign t_r1_c29_1 = p_1_28 << 1;
  assign t_r1_c29_2 = p_1_29 << 2;
  assign t_r1_c29_3 = p_1_30 << 1;
  assign t_r1_c29_4 = p_2_29 << 1;
  assign t_r1_c29_5 = t_r1_c29_0 + p_0_28;
  assign t_r1_c29_6 = t_r1_c29_1 + p_0_30;
  assign t_r1_c29_7 = t_r1_c29_2 + t_r1_c29_3;
  assign t_r1_c29_8 = t_r1_c29_4 + p_2_28;
  assign t_r1_c29_9 = t_r1_c29_5 + t_r1_c29_6;
  assign t_r1_c29_10 = t_r1_c29_7 + t_r1_c29_8;
  assign t_r1_c29_11 = t_r1_c29_9 + t_r1_c29_10;
  assign t_r1_c29_12 = t_r1_c29_11 + p_2_30;
  assign out_1_29 = t_r1_c29_12 >> 4;

  assign t_r1_c30_0 = p_0_30 << 1;
  assign t_r1_c30_1 = p_1_29 << 1;
  assign t_r1_c30_2 = p_1_30 << 2;
  assign t_r1_c30_3 = p_1_31 << 1;
  assign t_r1_c30_4 = p_2_30 << 1;
  assign t_r1_c30_5 = t_r1_c30_0 + p_0_29;
  assign t_r1_c30_6 = t_r1_c30_1 + p_0_31;
  assign t_r1_c30_7 = t_r1_c30_2 + t_r1_c30_3;
  assign t_r1_c30_8 = t_r1_c30_4 + p_2_29;
  assign t_r1_c30_9 = t_r1_c30_5 + t_r1_c30_6;
  assign t_r1_c30_10 = t_r1_c30_7 + t_r1_c30_8;
  assign t_r1_c30_11 = t_r1_c30_9 + t_r1_c30_10;
  assign t_r1_c30_12 = t_r1_c30_11 + p_2_31;
  assign out_1_30 = t_r1_c30_12 >> 4;

  assign t_r1_c31_0 = p_0_31 << 1;
  assign t_r1_c31_1 = p_1_30 << 1;
  assign t_r1_c31_2 = p_1_31 << 2;
  assign t_r1_c31_3 = p_1_32 << 1;
  assign t_r1_c31_4 = p_2_31 << 1;
  assign t_r1_c31_5 = t_r1_c31_0 + p_0_30;
  assign t_r1_c31_6 = t_r1_c31_1 + p_0_32;
  assign t_r1_c31_7 = t_r1_c31_2 + t_r1_c31_3;
  assign t_r1_c31_8 = t_r1_c31_4 + p_2_30;
  assign t_r1_c31_9 = t_r1_c31_5 + t_r1_c31_6;
  assign t_r1_c31_10 = t_r1_c31_7 + t_r1_c31_8;
  assign t_r1_c31_11 = t_r1_c31_9 + t_r1_c31_10;
  assign t_r1_c31_12 = t_r1_c31_11 + p_2_32;
  assign out_1_31 = t_r1_c31_12 >> 4;

  assign t_r1_c32_0 = p_0_32 << 1;
  assign t_r1_c32_1 = p_1_31 << 1;
  assign t_r1_c32_2 = p_1_32 << 2;
  assign t_r1_c32_3 = p_1_33 << 1;
  assign t_r1_c32_4 = p_2_32 << 1;
  assign t_r1_c32_5 = t_r1_c32_0 + p_0_31;
  assign t_r1_c32_6 = t_r1_c32_1 + p_0_33;
  assign t_r1_c32_7 = t_r1_c32_2 + t_r1_c32_3;
  assign t_r1_c32_8 = t_r1_c32_4 + p_2_31;
  assign t_r1_c32_9 = t_r1_c32_5 + t_r1_c32_6;
  assign t_r1_c32_10 = t_r1_c32_7 + t_r1_c32_8;
  assign t_r1_c32_11 = t_r1_c32_9 + t_r1_c32_10;
  assign t_r1_c32_12 = t_r1_c32_11 + p_2_33;
  assign out_1_32 = t_r1_c32_12 >> 4;

  assign t_r1_c33_0 = p_0_33 << 1;
  assign t_r1_c33_1 = p_1_32 << 1;
  assign t_r1_c33_2 = p_1_33 << 2;
  assign t_r1_c33_3 = p_1_34 << 1;
  assign t_r1_c33_4 = p_2_33 << 1;
  assign t_r1_c33_5 = t_r1_c33_0 + p_0_32;
  assign t_r1_c33_6 = t_r1_c33_1 + p_0_34;
  assign t_r1_c33_7 = t_r1_c33_2 + t_r1_c33_3;
  assign t_r1_c33_8 = t_r1_c33_4 + p_2_32;
  assign t_r1_c33_9 = t_r1_c33_5 + t_r1_c33_6;
  assign t_r1_c33_10 = t_r1_c33_7 + t_r1_c33_8;
  assign t_r1_c33_11 = t_r1_c33_9 + t_r1_c33_10;
  assign t_r1_c33_12 = t_r1_c33_11 + p_2_34;
  assign out_1_33 = t_r1_c33_12 >> 4;

  assign t_r1_c34_0 = p_0_34 << 1;
  assign t_r1_c34_1 = p_1_33 << 1;
  assign t_r1_c34_2 = p_1_34 << 2;
  assign t_r1_c34_3 = p_1_35 << 1;
  assign t_r1_c34_4 = p_2_34 << 1;
  assign t_r1_c34_5 = t_r1_c34_0 + p_0_33;
  assign t_r1_c34_6 = t_r1_c34_1 + p_0_35;
  assign t_r1_c34_7 = t_r1_c34_2 + t_r1_c34_3;
  assign t_r1_c34_8 = t_r1_c34_4 + p_2_33;
  assign t_r1_c34_9 = t_r1_c34_5 + t_r1_c34_6;
  assign t_r1_c34_10 = t_r1_c34_7 + t_r1_c34_8;
  assign t_r1_c34_11 = t_r1_c34_9 + t_r1_c34_10;
  assign t_r1_c34_12 = t_r1_c34_11 + p_2_35;
  assign out_1_34 = t_r1_c34_12 >> 4;

  assign t_r1_c35_0 = p_0_35 << 1;
  assign t_r1_c35_1 = p_1_34 << 1;
  assign t_r1_c35_2 = p_1_35 << 2;
  assign t_r1_c35_3 = p_1_36 << 1;
  assign t_r1_c35_4 = p_2_35 << 1;
  assign t_r1_c35_5 = t_r1_c35_0 + p_0_34;
  assign t_r1_c35_6 = t_r1_c35_1 + p_0_36;
  assign t_r1_c35_7 = t_r1_c35_2 + t_r1_c35_3;
  assign t_r1_c35_8 = t_r1_c35_4 + p_2_34;
  assign t_r1_c35_9 = t_r1_c35_5 + t_r1_c35_6;
  assign t_r1_c35_10 = t_r1_c35_7 + t_r1_c35_8;
  assign t_r1_c35_11 = t_r1_c35_9 + t_r1_c35_10;
  assign t_r1_c35_12 = t_r1_c35_11 + p_2_36;
  assign out_1_35 = t_r1_c35_12 >> 4;

  assign t_r1_c36_0 = p_0_36 << 1;
  assign t_r1_c36_1 = p_1_35 << 1;
  assign t_r1_c36_2 = p_1_36 << 2;
  assign t_r1_c36_3 = p_1_37 << 1;
  assign t_r1_c36_4 = p_2_36 << 1;
  assign t_r1_c36_5 = t_r1_c36_0 + p_0_35;
  assign t_r1_c36_6 = t_r1_c36_1 + p_0_37;
  assign t_r1_c36_7 = t_r1_c36_2 + t_r1_c36_3;
  assign t_r1_c36_8 = t_r1_c36_4 + p_2_35;
  assign t_r1_c36_9 = t_r1_c36_5 + t_r1_c36_6;
  assign t_r1_c36_10 = t_r1_c36_7 + t_r1_c36_8;
  assign t_r1_c36_11 = t_r1_c36_9 + t_r1_c36_10;
  assign t_r1_c36_12 = t_r1_c36_11 + p_2_37;
  assign out_1_36 = t_r1_c36_12 >> 4;

  assign t_r1_c37_0 = p_0_37 << 1;
  assign t_r1_c37_1 = p_1_36 << 1;
  assign t_r1_c37_2 = p_1_37 << 2;
  assign t_r1_c37_3 = p_1_38 << 1;
  assign t_r1_c37_4 = p_2_37 << 1;
  assign t_r1_c37_5 = t_r1_c37_0 + p_0_36;
  assign t_r1_c37_6 = t_r1_c37_1 + p_0_38;
  assign t_r1_c37_7 = t_r1_c37_2 + t_r1_c37_3;
  assign t_r1_c37_8 = t_r1_c37_4 + p_2_36;
  assign t_r1_c37_9 = t_r1_c37_5 + t_r1_c37_6;
  assign t_r1_c37_10 = t_r1_c37_7 + t_r1_c37_8;
  assign t_r1_c37_11 = t_r1_c37_9 + t_r1_c37_10;
  assign t_r1_c37_12 = t_r1_c37_11 + p_2_38;
  assign out_1_37 = t_r1_c37_12 >> 4;

  assign t_r1_c38_0 = p_0_38 << 1;
  assign t_r1_c38_1 = p_1_37 << 1;
  assign t_r1_c38_2 = p_1_38 << 2;
  assign t_r1_c38_3 = p_1_39 << 1;
  assign t_r1_c38_4 = p_2_38 << 1;
  assign t_r1_c38_5 = t_r1_c38_0 + p_0_37;
  assign t_r1_c38_6 = t_r1_c38_1 + p_0_39;
  assign t_r1_c38_7 = t_r1_c38_2 + t_r1_c38_3;
  assign t_r1_c38_8 = t_r1_c38_4 + p_2_37;
  assign t_r1_c38_9 = t_r1_c38_5 + t_r1_c38_6;
  assign t_r1_c38_10 = t_r1_c38_7 + t_r1_c38_8;
  assign t_r1_c38_11 = t_r1_c38_9 + t_r1_c38_10;
  assign t_r1_c38_12 = t_r1_c38_11 + p_2_39;
  assign out_1_38 = t_r1_c38_12 >> 4;

  assign t_r1_c39_0 = p_0_39 << 1;
  assign t_r1_c39_1 = p_1_38 << 1;
  assign t_r1_c39_2 = p_1_39 << 2;
  assign t_r1_c39_3 = p_1_40 << 1;
  assign t_r1_c39_4 = p_2_39 << 1;
  assign t_r1_c39_5 = t_r1_c39_0 + p_0_38;
  assign t_r1_c39_6 = t_r1_c39_1 + p_0_40;
  assign t_r1_c39_7 = t_r1_c39_2 + t_r1_c39_3;
  assign t_r1_c39_8 = t_r1_c39_4 + p_2_38;
  assign t_r1_c39_9 = t_r1_c39_5 + t_r1_c39_6;
  assign t_r1_c39_10 = t_r1_c39_7 + t_r1_c39_8;
  assign t_r1_c39_11 = t_r1_c39_9 + t_r1_c39_10;
  assign t_r1_c39_12 = t_r1_c39_11 + p_2_40;
  assign out_1_39 = t_r1_c39_12 >> 4;

  assign t_r1_c40_0 = p_0_40 << 1;
  assign t_r1_c40_1 = p_1_39 << 1;
  assign t_r1_c40_2 = p_1_40 << 2;
  assign t_r1_c40_3 = p_1_41 << 1;
  assign t_r1_c40_4 = p_2_40 << 1;
  assign t_r1_c40_5 = t_r1_c40_0 + p_0_39;
  assign t_r1_c40_6 = t_r1_c40_1 + p_0_41;
  assign t_r1_c40_7 = t_r1_c40_2 + t_r1_c40_3;
  assign t_r1_c40_8 = t_r1_c40_4 + p_2_39;
  assign t_r1_c40_9 = t_r1_c40_5 + t_r1_c40_6;
  assign t_r1_c40_10 = t_r1_c40_7 + t_r1_c40_8;
  assign t_r1_c40_11 = t_r1_c40_9 + t_r1_c40_10;
  assign t_r1_c40_12 = t_r1_c40_11 + p_2_41;
  assign out_1_40 = t_r1_c40_12 >> 4;

  assign t_r1_c41_0 = p_0_41 << 1;
  assign t_r1_c41_1 = p_1_40 << 1;
  assign t_r1_c41_2 = p_1_41 << 2;
  assign t_r1_c41_3 = p_1_42 << 1;
  assign t_r1_c41_4 = p_2_41 << 1;
  assign t_r1_c41_5 = t_r1_c41_0 + p_0_40;
  assign t_r1_c41_6 = t_r1_c41_1 + p_0_42;
  assign t_r1_c41_7 = t_r1_c41_2 + t_r1_c41_3;
  assign t_r1_c41_8 = t_r1_c41_4 + p_2_40;
  assign t_r1_c41_9 = t_r1_c41_5 + t_r1_c41_6;
  assign t_r1_c41_10 = t_r1_c41_7 + t_r1_c41_8;
  assign t_r1_c41_11 = t_r1_c41_9 + t_r1_c41_10;
  assign t_r1_c41_12 = t_r1_c41_11 + p_2_42;
  assign out_1_41 = t_r1_c41_12 >> 4;

  assign t_r1_c42_0 = p_0_42 << 1;
  assign t_r1_c42_1 = p_1_41 << 1;
  assign t_r1_c42_2 = p_1_42 << 2;
  assign t_r1_c42_3 = p_1_43 << 1;
  assign t_r1_c42_4 = p_2_42 << 1;
  assign t_r1_c42_5 = t_r1_c42_0 + p_0_41;
  assign t_r1_c42_6 = t_r1_c42_1 + p_0_43;
  assign t_r1_c42_7 = t_r1_c42_2 + t_r1_c42_3;
  assign t_r1_c42_8 = t_r1_c42_4 + p_2_41;
  assign t_r1_c42_9 = t_r1_c42_5 + t_r1_c42_6;
  assign t_r1_c42_10 = t_r1_c42_7 + t_r1_c42_8;
  assign t_r1_c42_11 = t_r1_c42_9 + t_r1_c42_10;
  assign t_r1_c42_12 = t_r1_c42_11 + p_2_43;
  assign out_1_42 = t_r1_c42_12 >> 4;

  assign t_r1_c43_0 = p_0_43 << 1;
  assign t_r1_c43_1 = p_1_42 << 1;
  assign t_r1_c43_2 = p_1_43 << 2;
  assign t_r1_c43_3 = p_1_44 << 1;
  assign t_r1_c43_4 = p_2_43 << 1;
  assign t_r1_c43_5 = t_r1_c43_0 + p_0_42;
  assign t_r1_c43_6 = t_r1_c43_1 + p_0_44;
  assign t_r1_c43_7 = t_r1_c43_2 + t_r1_c43_3;
  assign t_r1_c43_8 = t_r1_c43_4 + p_2_42;
  assign t_r1_c43_9 = t_r1_c43_5 + t_r1_c43_6;
  assign t_r1_c43_10 = t_r1_c43_7 + t_r1_c43_8;
  assign t_r1_c43_11 = t_r1_c43_9 + t_r1_c43_10;
  assign t_r1_c43_12 = t_r1_c43_11 + p_2_44;
  assign out_1_43 = t_r1_c43_12 >> 4;

  assign t_r1_c44_0 = p_0_44 << 1;
  assign t_r1_c44_1 = p_1_43 << 1;
  assign t_r1_c44_2 = p_1_44 << 2;
  assign t_r1_c44_3 = p_1_45 << 1;
  assign t_r1_c44_4 = p_2_44 << 1;
  assign t_r1_c44_5 = t_r1_c44_0 + p_0_43;
  assign t_r1_c44_6 = t_r1_c44_1 + p_0_45;
  assign t_r1_c44_7 = t_r1_c44_2 + t_r1_c44_3;
  assign t_r1_c44_8 = t_r1_c44_4 + p_2_43;
  assign t_r1_c44_9 = t_r1_c44_5 + t_r1_c44_6;
  assign t_r1_c44_10 = t_r1_c44_7 + t_r1_c44_8;
  assign t_r1_c44_11 = t_r1_c44_9 + t_r1_c44_10;
  assign t_r1_c44_12 = t_r1_c44_11 + p_2_45;
  assign out_1_44 = t_r1_c44_12 >> 4;

  assign t_r1_c45_0 = p_0_45 << 1;
  assign t_r1_c45_1 = p_1_44 << 1;
  assign t_r1_c45_2 = p_1_45 << 2;
  assign t_r1_c45_3 = p_1_46 << 1;
  assign t_r1_c45_4 = p_2_45 << 1;
  assign t_r1_c45_5 = t_r1_c45_0 + p_0_44;
  assign t_r1_c45_6 = t_r1_c45_1 + p_0_46;
  assign t_r1_c45_7 = t_r1_c45_2 + t_r1_c45_3;
  assign t_r1_c45_8 = t_r1_c45_4 + p_2_44;
  assign t_r1_c45_9 = t_r1_c45_5 + t_r1_c45_6;
  assign t_r1_c45_10 = t_r1_c45_7 + t_r1_c45_8;
  assign t_r1_c45_11 = t_r1_c45_9 + t_r1_c45_10;
  assign t_r1_c45_12 = t_r1_c45_11 + p_2_46;
  assign out_1_45 = t_r1_c45_12 >> 4;

  assign t_r1_c46_0 = p_0_46 << 1;
  assign t_r1_c46_1 = p_1_45 << 1;
  assign t_r1_c46_2 = p_1_46 << 2;
  assign t_r1_c46_3 = p_1_47 << 1;
  assign t_r1_c46_4 = p_2_46 << 1;
  assign t_r1_c46_5 = t_r1_c46_0 + p_0_45;
  assign t_r1_c46_6 = t_r1_c46_1 + p_0_47;
  assign t_r1_c46_7 = t_r1_c46_2 + t_r1_c46_3;
  assign t_r1_c46_8 = t_r1_c46_4 + p_2_45;
  assign t_r1_c46_9 = t_r1_c46_5 + t_r1_c46_6;
  assign t_r1_c46_10 = t_r1_c46_7 + t_r1_c46_8;
  assign t_r1_c46_11 = t_r1_c46_9 + t_r1_c46_10;
  assign t_r1_c46_12 = t_r1_c46_11 + p_2_47;
  assign out_1_46 = t_r1_c46_12 >> 4;

  assign t_r1_c47_0 = p_0_47 << 1;
  assign t_r1_c47_1 = p_1_46 << 1;
  assign t_r1_c47_2 = p_1_47 << 2;
  assign t_r1_c47_3 = p_1_48 << 1;
  assign t_r1_c47_4 = p_2_47 << 1;
  assign t_r1_c47_5 = t_r1_c47_0 + p_0_46;
  assign t_r1_c47_6 = t_r1_c47_1 + p_0_48;
  assign t_r1_c47_7 = t_r1_c47_2 + t_r1_c47_3;
  assign t_r1_c47_8 = t_r1_c47_4 + p_2_46;
  assign t_r1_c47_9 = t_r1_c47_5 + t_r1_c47_6;
  assign t_r1_c47_10 = t_r1_c47_7 + t_r1_c47_8;
  assign t_r1_c47_11 = t_r1_c47_9 + t_r1_c47_10;
  assign t_r1_c47_12 = t_r1_c47_11 + p_2_48;
  assign out_1_47 = t_r1_c47_12 >> 4;

  assign t_r1_c48_0 = p_0_48 << 1;
  assign t_r1_c48_1 = p_1_47 << 1;
  assign t_r1_c48_2 = p_1_48 << 2;
  assign t_r1_c48_3 = p_1_49 << 1;
  assign t_r1_c48_4 = p_2_48 << 1;
  assign t_r1_c48_5 = t_r1_c48_0 + p_0_47;
  assign t_r1_c48_6 = t_r1_c48_1 + p_0_49;
  assign t_r1_c48_7 = t_r1_c48_2 + t_r1_c48_3;
  assign t_r1_c48_8 = t_r1_c48_4 + p_2_47;
  assign t_r1_c48_9 = t_r1_c48_5 + t_r1_c48_6;
  assign t_r1_c48_10 = t_r1_c48_7 + t_r1_c48_8;
  assign t_r1_c48_11 = t_r1_c48_9 + t_r1_c48_10;
  assign t_r1_c48_12 = t_r1_c48_11 + p_2_49;
  assign out_1_48 = t_r1_c48_12 >> 4;

  assign t_r1_c49_0 = p_0_49 << 1;
  assign t_r1_c49_1 = p_1_48 << 1;
  assign t_r1_c49_2 = p_1_49 << 2;
  assign t_r1_c49_3 = p_1_50 << 1;
  assign t_r1_c49_4 = p_2_49 << 1;
  assign t_r1_c49_5 = t_r1_c49_0 + p_0_48;
  assign t_r1_c49_6 = t_r1_c49_1 + p_0_50;
  assign t_r1_c49_7 = t_r1_c49_2 + t_r1_c49_3;
  assign t_r1_c49_8 = t_r1_c49_4 + p_2_48;
  assign t_r1_c49_9 = t_r1_c49_5 + t_r1_c49_6;
  assign t_r1_c49_10 = t_r1_c49_7 + t_r1_c49_8;
  assign t_r1_c49_11 = t_r1_c49_9 + t_r1_c49_10;
  assign t_r1_c49_12 = t_r1_c49_11 + p_2_50;
  assign out_1_49 = t_r1_c49_12 >> 4;

  assign t_r1_c50_0 = p_0_50 << 1;
  assign t_r1_c50_1 = p_1_49 << 1;
  assign t_r1_c50_2 = p_1_50 << 2;
  assign t_r1_c50_3 = p_1_51 << 1;
  assign t_r1_c50_4 = p_2_50 << 1;
  assign t_r1_c50_5 = t_r1_c50_0 + p_0_49;
  assign t_r1_c50_6 = t_r1_c50_1 + p_0_51;
  assign t_r1_c50_7 = t_r1_c50_2 + t_r1_c50_3;
  assign t_r1_c50_8 = t_r1_c50_4 + p_2_49;
  assign t_r1_c50_9 = t_r1_c50_5 + t_r1_c50_6;
  assign t_r1_c50_10 = t_r1_c50_7 + t_r1_c50_8;
  assign t_r1_c50_11 = t_r1_c50_9 + t_r1_c50_10;
  assign t_r1_c50_12 = t_r1_c50_11 + p_2_51;
  assign out_1_50 = t_r1_c50_12 >> 4;

  assign t_r1_c51_0 = p_0_51 << 1;
  assign t_r1_c51_1 = p_1_50 << 1;
  assign t_r1_c51_2 = p_1_51 << 2;
  assign t_r1_c51_3 = p_1_52 << 1;
  assign t_r1_c51_4 = p_2_51 << 1;
  assign t_r1_c51_5 = t_r1_c51_0 + p_0_50;
  assign t_r1_c51_6 = t_r1_c51_1 + p_0_52;
  assign t_r1_c51_7 = t_r1_c51_2 + t_r1_c51_3;
  assign t_r1_c51_8 = t_r1_c51_4 + p_2_50;
  assign t_r1_c51_9 = t_r1_c51_5 + t_r1_c51_6;
  assign t_r1_c51_10 = t_r1_c51_7 + t_r1_c51_8;
  assign t_r1_c51_11 = t_r1_c51_9 + t_r1_c51_10;
  assign t_r1_c51_12 = t_r1_c51_11 + p_2_52;
  assign out_1_51 = t_r1_c51_12 >> 4;

  assign t_r1_c52_0 = p_0_52 << 1;
  assign t_r1_c52_1 = p_1_51 << 1;
  assign t_r1_c52_2 = p_1_52 << 2;
  assign t_r1_c52_3 = p_1_53 << 1;
  assign t_r1_c52_4 = p_2_52 << 1;
  assign t_r1_c52_5 = t_r1_c52_0 + p_0_51;
  assign t_r1_c52_6 = t_r1_c52_1 + p_0_53;
  assign t_r1_c52_7 = t_r1_c52_2 + t_r1_c52_3;
  assign t_r1_c52_8 = t_r1_c52_4 + p_2_51;
  assign t_r1_c52_9 = t_r1_c52_5 + t_r1_c52_6;
  assign t_r1_c52_10 = t_r1_c52_7 + t_r1_c52_8;
  assign t_r1_c52_11 = t_r1_c52_9 + t_r1_c52_10;
  assign t_r1_c52_12 = t_r1_c52_11 + p_2_53;
  assign out_1_52 = t_r1_c52_12 >> 4;

  assign t_r1_c53_0 = p_0_53 << 1;
  assign t_r1_c53_1 = p_1_52 << 1;
  assign t_r1_c53_2 = p_1_53 << 2;
  assign t_r1_c53_3 = p_1_54 << 1;
  assign t_r1_c53_4 = p_2_53 << 1;
  assign t_r1_c53_5 = t_r1_c53_0 + p_0_52;
  assign t_r1_c53_6 = t_r1_c53_1 + p_0_54;
  assign t_r1_c53_7 = t_r1_c53_2 + t_r1_c53_3;
  assign t_r1_c53_8 = t_r1_c53_4 + p_2_52;
  assign t_r1_c53_9 = t_r1_c53_5 + t_r1_c53_6;
  assign t_r1_c53_10 = t_r1_c53_7 + t_r1_c53_8;
  assign t_r1_c53_11 = t_r1_c53_9 + t_r1_c53_10;
  assign t_r1_c53_12 = t_r1_c53_11 + p_2_54;
  assign out_1_53 = t_r1_c53_12 >> 4;

  assign t_r1_c54_0 = p_0_54 << 1;
  assign t_r1_c54_1 = p_1_53 << 1;
  assign t_r1_c54_2 = p_1_54 << 2;
  assign t_r1_c54_3 = p_1_55 << 1;
  assign t_r1_c54_4 = p_2_54 << 1;
  assign t_r1_c54_5 = t_r1_c54_0 + p_0_53;
  assign t_r1_c54_6 = t_r1_c54_1 + p_0_55;
  assign t_r1_c54_7 = t_r1_c54_2 + t_r1_c54_3;
  assign t_r1_c54_8 = t_r1_c54_4 + p_2_53;
  assign t_r1_c54_9 = t_r1_c54_5 + t_r1_c54_6;
  assign t_r1_c54_10 = t_r1_c54_7 + t_r1_c54_8;
  assign t_r1_c54_11 = t_r1_c54_9 + t_r1_c54_10;
  assign t_r1_c54_12 = t_r1_c54_11 + p_2_55;
  assign out_1_54 = t_r1_c54_12 >> 4;

  assign t_r1_c55_0 = p_0_55 << 1;
  assign t_r1_c55_1 = p_1_54 << 1;
  assign t_r1_c55_2 = p_1_55 << 2;
  assign t_r1_c55_3 = p_1_56 << 1;
  assign t_r1_c55_4 = p_2_55 << 1;
  assign t_r1_c55_5 = t_r1_c55_0 + p_0_54;
  assign t_r1_c55_6 = t_r1_c55_1 + p_0_56;
  assign t_r1_c55_7 = t_r1_c55_2 + t_r1_c55_3;
  assign t_r1_c55_8 = t_r1_c55_4 + p_2_54;
  assign t_r1_c55_9 = t_r1_c55_5 + t_r1_c55_6;
  assign t_r1_c55_10 = t_r1_c55_7 + t_r1_c55_8;
  assign t_r1_c55_11 = t_r1_c55_9 + t_r1_c55_10;
  assign t_r1_c55_12 = t_r1_c55_11 + p_2_56;
  assign out_1_55 = t_r1_c55_12 >> 4;

  assign t_r1_c56_0 = p_0_56 << 1;
  assign t_r1_c56_1 = p_1_55 << 1;
  assign t_r1_c56_2 = p_1_56 << 2;
  assign t_r1_c56_3 = p_1_57 << 1;
  assign t_r1_c56_4 = p_2_56 << 1;
  assign t_r1_c56_5 = t_r1_c56_0 + p_0_55;
  assign t_r1_c56_6 = t_r1_c56_1 + p_0_57;
  assign t_r1_c56_7 = t_r1_c56_2 + t_r1_c56_3;
  assign t_r1_c56_8 = t_r1_c56_4 + p_2_55;
  assign t_r1_c56_9 = t_r1_c56_5 + t_r1_c56_6;
  assign t_r1_c56_10 = t_r1_c56_7 + t_r1_c56_8;
  assign t_r1_c56_11 = t_r1_c56_9 + t_r1_c56_10;
  assign t_r1_c56_12 = t_r1_c56_11 + p_2_57;
  assign out_1_56 = t_r1_c56_12 >> 4;

  assign t_r1_c57_0 = p_0_57 << 1;
  assign t_r1_c57_1 = p_1_56 << 1;
  assign t_r1_c57_2 = p_1_57 << 2;
  assign t_r1_c57_3 = p_1_58 << 1;
  assign t_r1_c57_4 = p_2_57 << 1;
  assign t_r1_c57_5 = t_r1_c57_0 + p_0_56;
  assign t_r1_c57_6 = t_r1_c57_1 + p_0_58;
  assign t_r1_c57_7 = t_r1_c57_2 + t_r1_c57_3;
  assign t_r1_c57_8 = t_r1_c57_4 + p_2_56;
  assign t_r1_c57_9 = t_r1_c57_5 + t_r1_c57_6;
  assign t_r1_c57_10 = t_r1_c57_7 + t_r1_c57_8;
  assign t_r1_c57_11 = t_r1_c57_9 + t_r1_c57_10;
  assign t_r1_c57_12 = t_r1_c57_11 + p_2_58;
  assign out_1_57 = t_r1_c57_12 >> 4;

  assign t_r1_c58_0 = p_0_58 << 1;
  assign t_r1_c58_1 = p_1_57 << 1;
  assign t_r1_c58_2 = p_1_58 << 2;
  assign t_r1_c58_3 = p_1_59 << 1;
  assign t_r1_c58_4 = p_2_58 << 1;
  assign t_r1_c58_5 = t_r1_c58_0 + p_0_57;
  assign t_r1_c58_6 = t_r1_c58_1 + p_0_59;
  assign t_r1_c58_7 = t_r1_c58_2 + t_r1_c58_3;
  assign t_r1_c58_8 = t_r1_c58_4 + p_2_57;
  assign t_r1_c58_9 = t_r1_c58_5 + t_r1_c58_6;
  assign t_r1_c58_10 = t_r1_c58_7 + t_r1_c58_8;
  assign t_r1_c58_11 = t_r1_c58_9 + t_r1_c58_10;
  assign t_r1_c58_12 = t_r1_c58_11 + p_2_59;
  assign out_1_58 = t_r1_c58_12 >> 4;

  assign t_r1_c59_0 = p_0_59 << 1;
  assign t_r1_c59_1 = p_1_58 << 1;
  assign t_r1_c59_2 = p_1_59 << 2;
  assign t_r1_c59_3 = p_1_60 << 1;
  assign t_r1_c59_4 = p_2_59 << 1;
  assign t_r1_c59_5 = t_r1_c59_0 + p_0_58;
  assign t_r1_c59_6 = t_r1_c59_1 + p_0_60;
  assign t_r1_c59_7 = t_r1_c59_2 + t_r1_c59_3;
  assign t_r1_c59_8 = t_r1_c59_4 + p_2_58;
  assign t_r1_c59_9 = t_r1_c59_5 + t_r1_c59_6;
  assign t_r1_c59_10 = t_r1_c59_7 + t_r1_c59_8;
  assign t_r1_c59_11 = t_r1_c59_9 + t_r1_c59_10;
  assign t_r1_c59_12 = t_r1_c59_11 + p_2_60;
  assign out_1_59 = t_r1_c59_12 >> 4;

  assign t_r1_c60_0 = p_0_60 << 1;
  assign t_r1_c60_1 = p_1_59 << 1;
  assign t_r1_c60_2 = p_1_60 << 2;
  assign t_r1_c60_3 = p_1_61 << 1;
  assign t_r1_c60_4 = p_2_60 << 1;
  assign t_r1_c60_5 = t_r1_c60_0 + p_0_59;
  assign t_r1_c60_6 = t_r1_c60_1 + p_0_61;
  assign t_r1_c60_7 = t_r1_c60_2 + t_r1_c60_3;
  assign t_r1_c60_8 = t_r1_c60_4 + p_2_59;
  assign t_r1_c60_9 = t_r1_c60_5 + t_r1_c60_6;
  assign t_r1_c60_10 = t_r1_c60_7 + t_r1_c60_8;
  assign t_r1_c60_11 = t_r1_c60_9 + t_r1_c60_10;
  assign t_r1_c60_12 = t_r1_c60_11 + p_2_61;
  assign out_1_60 = t_r1_c60_12 >> 4;

  assign t_r1_c61_0 = p_0_61 << 1;
  assign t_r1_c61_1 = p_1_60 << 1;
  assign t_r1_c61_2 = p_1_61 << 2;
  assign t_r1_c61_3 = p_1_62 << 1;
  assign t_r1_c61_4 = p_2_61 << 1;
  assign t_r1_c61_5 = t_r1_c61_0 + p_0_60;
  assign t_r1_c61_6 = t_r1_c61_1 + p_0_62;
  assign t_r1_c61_7 = t_r1_c61_2 + t_r1_c61_3;
  assign t_r1_c61_8 = t_r1_c61_4 + p_2_60;
  assign t_r1_c61_9 = t_r1_c61_5 + t_r1_c61_6;
  assign t_r1_c61_10 = t_r1_c61_7 + t_r1_c61_8;
  assign t_r1_c61_11 = t_r1_c61_9 + t_r1_c61_10;
  assign t_r1_c61_12 = t_r1_c61_11 + p_2_62;
  assign out_1_61 = t_r1_c61_12 >> 4;

  assign t_r1_c62_0 = p_0_62 << 1;
  assign t_r1_c62_1 = p_1_61 << 1;
  assign t_r1_c62_2 = p_1_62 << 2;
  assign t_r1_c62_3 = p_1_63 << 1;
  assign t_r1_c62_4 = p_2_62 << 1;
  assign t_r1_c62_5 = t_r1_c62_0 + p_0_61;
  assign t_r1_c62_6 = t_r1_c62_1 + p_0_63;
  assign t_r1_c62_7 = t_r1_c62_2 + t_r1_c62_3;
  assign t_r1_c62_8 = t_r1_c62_4 + p_2_61;
  assign t_r1_c62_9 = t_r1_c62_5 + t_r1_c62_6;
  assign t_r1_c62_10 = t_r1_c62_7 + t_r1_c62_8;
  assign t_r1_c62_11 = t_r1_c62_9 + t_r1_c62_10;
  assign t_r1_c62_12 = t_r1_c62_11 + p_2_63;
  assign out_1_62 = t_r1_c62_12 >> 4;

  assign t_r1_c63_0 = p_0_63 << 1;
  assign t_r1_c63_1 = p_1_62 << 1;
  assign t_r1_c63_2 = p_1_63 << 2;
  assign t_r1_c63_3 = p_1_64 << 1;
  assign t_r1_c63_4 = p_2_63 << 1;
  assign t_r1_c63_5 = t_r1_c63_0 + p_0_62;
  assign t_r1_c63_6 = t_r1_c63_1 + p_0_64;
  assign t_r1_c63_7 = t_r1_c63_2 + t_r1_c63_3;
  assign t_r1_c63_8 = t_r1_c63_4 + p_2_62;
  assign t_r1_c63_9 = t_r1_c63_5 + t_r1_c63_6;
  assign t_r1_c63_10 = t_r1_c63_7 + t_r1_c63_8;
  assign t_r1_c63_11 = t_r1_c63_9 + t_r1_c63_10;
  assign t_r1_c63_12 = t_r1_c63_11 + p_2_64;
  assign out_1_63 = t_r1_c63_12 >> 4;

  assign t_r1_c64_0 = p_0_64 << 1;
  assign t_r1_c64_1 = p_1_63 << 1;
  assign t_r1_c64_2 = p_1_64 << 2;
  assign t_r1_c64_3 = p_1_65 << 1;
  assign t_r1_c64_4 = p_2_64 << 1;
  assign t_r1_c64_5 = t_r1_c64_0 + p_0_63;
  assign t_r1_c64_6 = t_r1_c64_1 + p_0_65;
  assign t_r1_c64_7 = t_r1_c64_2 + t_r1_c64_3;
  assign t_r1_c64_8 = t_r1_c64_4 + p_2_63;
  assign t_r1_c64_9 = t_r1_c64_5 + t_r1_c64_6;
  assign t_r1_c64_10 = t_r1_c64_7 + t_r1_c64_8;
  assign t_r1_c64_11 = t_r1_c64_9 + t_r1_c64_10;
  assign t_r1_c64_12 = t_r1_c64_11 + p_2_65;
  assign out_1_64 = t_r1_c64_12 >> 4;

  assign t_r2_c1_0 = p_1_1 << 1;
  assign t_r2_c1_1 = p_2_0 << 1;
  assign t_r2_c1_2 = p_2_1 << 2;
  assign t_r2_c1_3 = p_2_2 << 1;
  assign t_r2_c1_4 = p_3_1 << 1;
  assign t_r2_c1_5 = t_r2_c1_0 + p_1_0;
  assign t_r2_c1_6 = t_r2_c1_1 + p_1_2;
  assign t_r2_c1_7 = t_r2_c1_2 + t_r2_c1_3;
  assign t_r2_c1_8 = t_r2_c1_4 + p_3_0;
  assign t_r2_c1_9 = t_r2_c1_5 + t_r2_c1_6;
  assign t_r2_c1_10 = t_r2_c1_7 + t_r2_c1_8;
  assign t_r2_c1_11 = t_r2_c1_9 + t_r2_c1_10;
  assign t_r2_c1_12 = t_r2_c1_11 + p_3_2;
  assign out_2_1 = t_r2_c1_12 >> 4;

  assign t_r2_c2_0 = p_1_2 << 1;
  assign t_r2_c2_1 = p_2_1 << 1;
  assign t_r2_c2_2 = p_2_2 << 2;
  assign t_r2_c2_3 = p_2_3 << 1;
  assign t_r2_c2_4 = p_3_2 << 1;
  assign t_r2_c2_5 = t_r2_c2_0 + p_1_1;
  assign t_r2_c2_6 = t_r2_c2_1 + p_1_3;
  assign t_r2_c2_7 = t_r2_c2_2 + t_r2_c2_3;
  assign t_r2_c2_8 = t_r2_c2_4 + p_3_1;
  assign t_r2_c2_9 = t_r2_c2_5 + t_r2_c2_6;
  assign t_r2_c2_10 = t_r2_c2_7 + t_r2_c2_8;
  assign t_r2_c2_11 = t_r2_c2_9 + t_r2_c2_10;
  assign t_r2_c2_12 = t_r2_c2_11 + p_3_3;
  assign out_2_2 = t_r2_c2_12 >> 4;

  assign t_r2_c3_0 = p_1_3 << 1;
  assign t_r2_c3_1 = p_2_2 << 1;
  assign t_r2_c3_2 = p_2_3 << 2;
  assign t_r2_c3_3 = p_2_4 << 1;
  assign t_r2_c3_4 = p_3_3 << 1;
  assign t_r2_c3_5 = t_r2_c3_0 + p_1_2;
  assign t_r2_c3_6 = t_r2_c3_1 + p_1_4;
  assign t_r2_c3_7 = t_r2_c3_2 + t_r2_c3_3;
  assign t_r2_c3_8 = t_r2_c3_4 + p_3_2;
  assign t_r2_c3_9 = t_r2_c3_5 + t_r2_c3_6;
  assign t_r2_c3_10 = t_r2_c3_7 + t_r2_c3_8;
  assign t_r2_c3_11 = t_r2_c3_9 + t_r2_c3_10;
  assign t_r2_c3_12 = t_r2_c3_11 + p_3_4;
  assign out_2_3 = t_r2_c3_12 >> 4;

  assign t_r2_c4_0 = p_1_4 << 1;
  assign t_r2_c4_1 = p_2_3 << 1;
  assign t_r2_c4_2 = p_2_4 << 2;
  assign t_r2_c4_3 = p_2_5 << 1;
  assign t_r2_c4_4 = p_3_4 << 1;
  assign t_r2_c4_5 = t_r2_c4_0 + p_1_3;
  assign t_r2_c4_6 = t_r2_c4_1 + p_1_5;
  assign t_r2_c4_7 = t_r2_c4_2 + t_r2_c4_3;
  assign t_r2_c4_8 = t_r2_c4_4 + p_3_3;
  assign t_r2_c4_9 = t_r2_c4_5 + t_r2_c4_6;
  assign t_r2_c4_10 = t_r2_c4_7 + t_r2_c4_8;
  assign t_r2_c4_11 = t_r2_c4_9 + t_r2_c4_10;
  assign t_r2_c4_12 = t_r2_c4_11 + p_3_5;
  assign out_2_4 = t_r2_c4_12 >> 4;

  assign t_r2_c5_0 = p_1_5 << 1;
  assign t_r2_c5_1 = p_2_4 << 1;
  assign t_r2_c5_2 = p_2_5 << 2;
  assign t_r2_c5_3 = p_2_6 << 1;
  assign t_r2_c5_4 = p_3_5 << 1;
  assign t_r2_c5_5 = t_r2_c5_0 + p_1_4;
  assign t_r2_c5_6 = t_r2_c5_1 + p_1_6;
  assign t_r2_c5_7 = t_r2_c5_2 + t_r2_c5_3;
  assign t_r2_c5_8 = t_r2_c5_4 + p_3_4;
  assign t_r2_c5_9 = t_r2_c5_5 + t_r2_c5_6;
  assign t_r2_c5_10 = t_r2_c5_7 + t_r2_c5_8;
  assign t_r2_c5_11 = t_r2_c5_9 + t_r2_c5_10;
  assign t_r2_c5_12 = t_r2_c5_11 + p_3_6;
  assign out_2_5 = t_r2_c5_12 >> 4;

  assign t_r2_c6_0 = p_1_6 << 1;
  assign t_r2_c6_1 = p_2_5 << 1;
  assign t_r2_c6_2 = p_2_6 << 2;
  assign t_r2_c6_3 = p_2_7 << 1;
  assign t_r2_c6_4 = p_3_6 << 1;
  assign t_r2_c6_5 = t_r2_c6_0 + p_1_5;
  assign t_r2_c6_6 = t_r2_c6_1 + p_1_7;
  assign t_r2_c6_7 = t_r2_c6_2 + t_r2_c6_3;
  assign t_r2_c6_8 = t_r2_c6_4 + p_3_5;
  assign t_r2_c6_9 = t_r2_c6_5 + t_r2_c6_6;
  assign t_r2_c6_10 = t_r2_c6_7 + t_r2_c6_8;
  assign t_r2_c6_11 = t_r2_c6_9 + t_r2_c6_10;
  assign t_r2_c6_12 = t_r2_c6_11 + p_3_7;
  assign out_2_6 = t_r2_c6_12 >> 4;

  assign t_r2_c7_0 = p_1_7 << 1;
  assign t_r2_c7_1 = p_2_6 << 1;
  assign t_r2_c7_2 = p_2_7 << 2;
  assign t_r2_c7_3 = p_2_8 << 1;
  assign t_r2_c7_4 = p_3_7 << 1;
  assign t_r2_c7_5 = t_r2_c7_0 + p_1_6;
  assign t_r2_c7_6 = t_r2_c7_1 + p_1_8;
  assign t_r2_c7_7 = t_r2_c7_2 + t_r2_c7_3;
  assign t_r2_c7_8 = t_r2_c7_4 + p_3_6;
  assign t_r2_c7_9 = t_r2_c7_5 + t_r2_c7_6;
  assign t_r2_c7_10 = t_r2_c7_7 + t_r2_c7_8;
  assign t_r2_c7_11 = t_r2_c7_9 + t_r2_c7_10;
  assign t_r2_c7_12 = t_r2_c7_11 + p_3_8;
  assign out_2_7 = t_r2_c7_12 >> 4;

  assign t_r2_c8_0 = p_1_8 << 1;
  assign t_r2_c8_1 = p_2_7 << 1;
  assign t_r2_c8_2 = p_2_8 << 2;
  assign t_r2_c8_3 = p_2_9 << 1;
  assign t_r2_c8_4 = p_3_8 << 1;
  assign t_r2_c8_5 = t_r2_c8_0 + p_1_7;
  assign t_r2_c8_6 = t_r2_c8_1 + p_1_9;
  assign t_r2_c8_7 = t_r2_c8_2 + t_r2_c8_3;
  assign t_r2_c8_8 = t_r2_c8_4 + p_3_7;
  assign t_r2_c8_9 = t_r2_c8_5 + t_r2_c8_6;
  assign t_r2_c8_10 = t_r2_c8_7 + t_r2_c8_8;
  assign t_r2_c8_11 = t_r2_c8_9 + t_r2_c8_10;
  assign t_r2_c8_12 = t_r2_c8_11 + p_3_9;
  assign out_2_8 = t_r2_c8_12 >> 4;

  assign t_r2_c9_0 = p_1_9 << 1;
  assign t_r2_c9_1 = p_2_8 << 1;
  assign t_r2_c9_2 = p_2_9 << 2;
  assign t_r2_c9_3 = p_2_10 << 1;
  assign t_r2_c9_4 = p_3_9 << 1;
  assign t_r2_c9_5 = t_r2_c9_0 + p_1_8;
  assign t_r2_c9_6 = t_r2_c9_1 + p_1_10;
  assign t_r2_c9_7 = t_r2_c9_2 + t_r2_c9_3;
  assign t_r2_c9_8 = t_r2_c9_4 + p_3_8;
  assign t_r2_c9_9 = t_r2_c9_5 + t_r2_c9_6;
  assign t_r2_c9_10 = t_r2_c9_7 + t_r2_c9_8;
  assign t_r2_c9_11 = t_r2_c9_9 + t_r2_c9_10;
  assign t_r2_c9_12 = t_r2_c9_11 + p_3_10;
  assign out_2_9 = t_r2_c9_12 >> 4;

  assign t_r2_c10_0 = p_1_10 << 1;
  assign t_r2_c10_1 = p_2_9 << 1;
  assign t_r2_c10_2 = p_2_10 << 2;
  assign t_r2_c10_3 = p_2_11 << 1;
  assign t_r2_c10_4 = p_3_10 << 1;
  assign t_r2_c10_5 = t_r2_c10_0 + p_1_9;
  assign t_r2_c10_6 = t_r2_c10_1 + p_1_11;
  assign t_r2_c10_7 = t_r2_c10_2 + t_r2_c10_3;
  assign t_r2_c10_8 = t_r2_c10_4 + p_3_9;
  assign t_r2_c10_9 = t_r2_c10_5 + t_r2_c10_6;
  assign t_r2_c10_10 = t_r2_c10_7 + t_r2_c10_8;
  assign t_r2_c10_11 = t_r2_c10_9 + t_r2_c10_10;
  assign t_r2_c10_12 = t_r2_c10_11 + p_3_11;
  assign out_2_10 = t_r2_c10_12 >> 4;

  assign t_r2_c11_0 = p_1_11 << 1;
  assign t_r2_c11_1 = p_2_10 << 1;
  assign t_r2_c11_2 = p_2_11 << 2;
  assign t_r2_c11_3 = p_2_12 << 1;
  assign t_r2_c11_4 = p_3_11 << 1;
  assign t_r2_c11_5 = t_r2_c11_0 + p_1_10;
  assign t_r2_c11_6 = t_r2_c11_1 + p_1_12;
  assign t_r2_c11_7 = t_r2_c11_2 + t_r2_c11_3;
  assign t_r2_c11_8 = t_r2_c11_4 + p_3_10;
  assign t_r2_c11_9 = t_r2_c11_5 + t_r2_c11_6;
  assign t_r2_c11_10 = t_r2_c11_7 + t_r2_c11_8;
  assign t_r2_c11_11 = t_r2_c11_9 + t_r2_c11_10;
  assign t_r2_c11_12 = t_r2_c11_11 + p_3_12;
  assign out_2_11 = t_r2_c11_12 >> 4;

  assign t_r2_c12_0 = p_1_12 << 1;
  assign t_r2_c12_1 = p_2_11 << 1;
  assign t_r2_c12_2 = p_2_12 << 2;
  assign t_r2_c12_3 = p_2_13 << 1;
  assign t_r2_c12_4 = p_3_12 << 1;
  assign t_r2_c12_5 = t_r2_c12_0 + p_1_11;
  assign t_r2_c12_6 = t_r2_c12_1 + p_1_13;
  assign t_r2_c12_7 = t_r2_c12_2 + t_r2_c12_3;
  assign t_r2_c12_8 = t_r2_c12_4 + p_3_11;
  assign t_r2_c12_9 = t_r2_c12_5 + t_r2_c12_6;
  assign t_r2_c12_10 = t_r2_c12_7 + t_r2_c12_8;
  assign t_r2_c12_11 = t_r2_c12_9 + t_r2_c12_10;
  assign t_r2_c12_12 = t_r2_c12_11 + p_3_13;
  assign out_2_12 = t_r2_c12_12 >> 4;

  assign t_r2_c13_0 = p_1_13 << 1;
  assign t_r2_c13_1 = p_2_12 << 1;
  assign t_r2_c13_2 = p_2_13 << 2;
  assign t_r2_c13_3 = p_2_14 << 1;
  assign t_r2_c13_4 = p_3_13 << 1;
  assign t_r2_c13_5 = t_r2_c13_0 + p_1_12;
  assign t_r2_c13_6 = t_r2_c13_1 + p_1_14;
  assign t_r2_c13_7 = t_r2_c13_2 + t_r2_c13_3;
  assign t_r2_c13_8 = t_r2_c13_4 + p_3_12;
  assign t_r2_c13_9 = t_r2_c13_5 + t_r2_c13_6;
  assign t_r2_c13_10 = t_r2_c13_7 + t_r2_c13_8;
  assign t_r2_c13_11 = t_r2_c13_9 + t_r2_c13_10;
  assign t_r2_c13_12 = t_r2_c13_11 + p_3_14;
  assign out_2_13 = t_r2_c13_12 >> 4;

  assign t_r2_c14_0 = p_1_14 << 1;
  assign t_r2_c14_1 = p_2_13 << 1;
  assign t_r2_c14_2 = p_2_14 << 2;
  assign t_r2_c14_3 = p_2_15 << 1;
  assign t_r2_c14_4 = p_3_14 << 1;
  assign t_r2_c14_5 = t_r2_c14_0 + p_1_13;
  assign t_r2_c14_6 = t_r2_c14_1 + p_1_15;
  assign t_r2_c14_7 = t_r2_c14_2 + t_r2_c14_3;
  assign t_r2_c14_8 = t_r2_c14_4 + p_3_13;
  assign t_r2_c14_9 = t_r2_c14_5 + t_r2_c14_6;
  assign t_r2_c14_10 = t_r2_c14_7 + t_r2_c14_8;
  assign t_r2_c14_11 = t_r2_c14_9 + t_r2_c14_10;
  assign t_r2_c14_12 = t_r2_c14_11 + p_3_15;
  assign out_2_14 = t_r2_c14_12 >> 4;

  assign t_r2_c15_0 = p_1_15 << 1;
  assign t_r2_c15_1 = p_2_14 << 1;
  assign t_r2_c15_2 = p_2_15 << 2;
  assign t_r2_c15_3 = p_2_16 << 1;
  assign t_r2_c15_4 = p_3_15 << 1;
  assign t_r2_c15_5 = t_r2_c15_0 + p_1_14;
  assign t_r2_c15_6 = t_r2_c15_1 + p_1_16;
  assign t_r2_c15_7 = t_r2_c15_2 + t_r2_c15_3;
  assign t_r2_c15_8 = t_r2_c15_4 + p_3_14;
  assign t_r2_c15_9 = t_r2_c15_5 + t_r2_c15_6;
  assign t_r2_c15_10 = t_r2_c15_7 + t_r2_c15_8;
  assign t_r2_c15_11 = t_r2_c15_9 + t_r2_c15_10;
  assign t_r2_c15_12 = t_r2_c15_11 + p_3_16;
  assign out_2_15 = t_r2_c15_12 >> 4;

  assign t_r2_c16_0 = p_1_16 << 1;
  assign t_r2_c16_1 = p_2_15 << 1;
  assign t_r2_c16_2 = p_2_16 << 2;
  assign t_r2_c16_3 = p_2_17 << 1;
  assign t_r2_c16_4 = p_3_16 << 1;
  assign t_r2_c16_5 = t_r2_c16_0 + p_1_15;
  assign t_r2_c16_6 = t_r2_c16_1 + p_1_17;
  assign t_r2_c16_7 = t_r2_c16_2 + t_r2_c16_3;
  assign t_r2_c16_8 = t_r2_c16_4 + p_3_15;
  assign t_r2_c16_9 = t_r2_c16_5 + t_r2_c16_6;
  assign t_r2_c16_10 = t_r2_c16_7 + t_r2_c16_8;
  assign t_r2_c16_11 = t_r2_c16_9 + t_r2_c16_10;
  assign t_r2_c16_12 = t_r2_c16_11 + p_3_17;
  assign out_2_16 = t_r2_c16_12 >> 4;

  assign t_r2_c17_0 = p_1_17 << 1;
  assign t_r2_c17_1 = p_2_16 << 1;
  assign t_r2_c17_2 = p_2_17 << 2;
  assign t_r2_c17_3 = p_2_18 << 1;
  assign t_r2_c17_4 = p_3_17 << 1;
  assign t_r2_c17_5 = t_r2_c17_0 + p_1_16;
  assign t_r2_c17_6 = t_r2_c17_1 + p_1_18;
  assign t_r2_c17_7 = t_r2_c17_2 + t_r2_c17_3;
  assign t_r2_c17_8 = t_r2_c17_4 + p_3_16;
  assign t_r2_c17_9 = t_r2_c17_5 + t_r2_c17_6;
  assign t_r2_c17_10 = t_r2_c17_7 + t_r2_c17_8;
  assign t_r2_c17_11 = t_r2_c17_9 + t_r2_c17_10;
  assign t_r2_c17_12 = t_r2_c17_11 + p_3_18;
  assign out_2_17 = t_r2_c17_12 >> 4;

  assign t_r2_c18_0 = p_1_18 << 1;
  assign t_r2_c18_1 = p_2_17 << 1;
  assign t_r2_c18_2 = p_2_18 << 2;
  assign t_r2_c18_3 = p_2_19 << 1;
  assign t_r2_c18_4 = p_3_18 << 1;
  assign t_r2_c18_5 = t_r2_c18_0 + p_1_17;
  assign t_r2_c18_6 = t_r2_c18_1 + p_1_19;
  assign t_r2_c18_7 = t_r2_c18_2 + t_r2_c18_3;
  assign t_r2_c18_8 = t_r2_c18_4 + p_3_17;
  assign t_r2_c18_9 = t_r2_c18_5 + t_r2_c18_6;
  assign t_r2_c18_10 = t_r2_c18_7 + t_r2_c18_8;
  assign t_r2_c18_11 = t_r2_c18_9 + t_r2_c18_10;
  assign t_r2_c18_12 = t_r2_c18_11 + p_3_19;
  assign out_2_18 = t_r2_c18_12 >> 4;

  assign t_r2_c19_0 = p_1_19 << 1;
  assign t_r2_c19_1 = p_2_18 << 1;
  assign t_r2_c19_2 = p_2_19 << 2;
  assign t_r2_c19_3 = p_2_20 << 1;
  assign t_r2_c19_4 = p_3_19 << 1;
  assign t_r2_c19_5 = t_r2_c19_0 + p_1_18;
  assign t_r2_c19_6 = t_r2_c19_1 + p_1_20;
  assign t_r2_c19_7 = t_r2_c19_2 + t_r2_c19_3;
  assign t_r2_c19_8 = t_r2_c19_4 + p_3_18;
  assign t_r2_c19_9 = t_r2_c19_5 + t_r2_c19_6;
  assign t_r2_c19_10 = t_r2_c19_7 + t_r2_c19_8;
  assign t_r2_c19_11 = t_r2_c19_9 + t_r2_c19_10;
  assign t_r2_c19_12 = t_r2_c19_11 + p_3_20;
  assign out_2_19 = t_r2_c19_12 >> 4;

  assign t_r2_c20_0 = p_1_20 << 1;
  assign t_r2_c20_1 = p_2_19 << 1;
  assign t_r2_c20_2 = p_2_20 << 2;
  assign t_r2_c20_3 = p_2_21 << 1;
  assign t_r2_c20_4 = p_3_20 << 1;
  assign t_r2_c20_5 = t_r2_c20_0 + p_1_19;
  assign t_r2_c20_6 = t_r2_c20_1 + p_1_21;
  assign t_r2_c20_7 = t_r2_c20_2 + t_r2_c20_3;
  assign t_r2_c20_8 = t_r2_c20_4 + p_3_19;
  assign t_r2_c20_9 = t_r2_c20_5 + t_r2_c20_6;
  assign t_r2_c20_10 = t_r2_c20_7 + t_r2_c20_8;
  assign t_r2_c20_11 = t_r2_c20_9 + t_r2_c20_10;
  assign t_r2_c20_12 = t_r2_c20_11 + p_3_21;
  assign out_2_20 = t_r2_c20_12 >> 4;

  assign t_r2_c21_0 = p_1_21 << 1;
  assign t_r2_c21_1 = p_2_20 << 1;
  assign t_r2_c21_2 = p_2_21 << 2;
  assign t_r2_c21_3 = p_2_22 << 1;
  assign t_r2_c21_4 = p_3_21 << 1;
  assign t_r2_c21_5 = t_r2_c21_0 + p_1_20;
  assign t_r2_c21_6 = t_r2_c21_1 + p_1_22;
  assign t_r2_c21_7 = t_r2_c21_2 + t_r2_c21_3;
  assign t_r2_c21_8 = t_r2_c21_4 + p_3_20;
  assign t_r2_c21_9 = t_r2_c21_5 + t_r2_c21_6;
  assign t_r2_c21_10 = t_r2_c21_7 + t_r2_c21_8;
  assign t_r2_c21_11 = t_r2_c21_9 + t_r2_c21_10;
  assign t_r2_c21_12 = t_r2_c21_11 + p_3_22;
  assign out_2_21 = t_r2_c21_12 >> 4;

  assign t_r2_c22_0 = p_1_22 << 1;
  assign t_r2_c22_1 = p_2_21 << 1;
  assign t_r2_c22_2 = p_2_22 << 2;
  assign t_r2_c22_3 = p_2_23 << 1;
  assign t_r2_c22_4 = p_3_22 << 1;
  assign t_r2_c22_5 = t_r2_c22_0 + p_1_21;
  assign t_r2_c22_6 = t_r2_c22_1 + p_1_23;
  assign t_r2_c22_7 = t_r2_c22_2 + t_r2_c22_3;
  assign t_r2_c22_8 = t_r2_c22_4 + p_3_21;
  assign t_r2_c22_9 = t_r2_c22_5 + t_r2_c22_6;
  assign t_r2_c22_10 = t_r2_c22_7 + t_r2_c22_8;
  assign t_r2_c22_11 = t_r2_c22_9 + t_r2_c22_10;
  assign t_r2_c22_12 = t_r2_c22_11 + p_3_23;
  assign out_2_22 = t_r2_c22_12 >> 4;

  assign t_r2_c23_0 = p_1_23 << 1;
  assign t_r2_c23_1 = p_2_22 << 1;
  assign t_r2_c23_2 = p_2_23 << 2;
  assign t_r2_c23_3 = p_2_24 << 1;
  assign t_r2_c23_4 = p_3_23 << 1;
  assign t_r2_c23_5 = t_r2_c23_0 + p_1_22;
  assign t_r2_c23_6 = t_r2_c23_1 + p_1_24;
  assign t_r2_c23_7 = t_r2_c23_2 + t_r2_c23_3;
  assign t_r2_c23_8 = t_r2_c23_4 + p_3_22;
  assign t_r2_c23_9 = t_r2_c23_5 + t_r2_c23_6;
  assign t_r2_c23_10 = t_r2_c23_7 + t_r2_c23_8;
  assign t_r2_c23_11 = t_r2_c23_9 + t_r2_c23_10;
  assign t_r2_c23_12 = t_r2_c23_11 + p_3_24;
  assign out_2_23 = t_r2_c23_12 >> 4;

  assign t_r2_c24_0 = p_1_24 << 1;
  assign t_r2_c24_1 = p_2_23 << 1;
  assign t_r2_c24_2 = p_2_24 << 2;
  assign t_r2_c24_3 = p_2_25 << 1;
  assign t_r2_c24_4 = p_3_24 << 1;
  assign t_r2_c24_5 = t_r2_c24_0 + p_1_23;
  assign t_r2_c24_6 = t_r2_c24_1 + p_1_25;
  assign t_r2_c24_7 = t_r2_c24_2 + t_r2_c24_3;
  assign t_r2_c24_8 = t_r2_c24_4 + p_3_23;
  assign t_r2_c24_9 = t_r2_c24_5 + t_r2_c24_6;
  assign t_r2_c24_10 = t_r2_c24_7 + t_r2_c24_8;
  assign t_r2_c24_11 = t_r2_c24_9 + t_r2_c24_10;
  assign t_r2_c24_12 = t_r2_c24_11 + p_3_25;
  assign out_2_24 = t_r2_c24_12 >> 4;

  assign t_r2_c25_0 = p_1_25 << 1;
  assign t_r2_c25_1 = p_2_24 << 1;
  assign t_r2_c25_2 = p_2_25 << 2;
  assign t_r2_c25_3 = p_2_26 << 1;
  assign t_r2_c25_4 = p_3_25 << 1;
  assign t_r2_c25_5 = t_r2_c25_0 + p_1_24;
  assign t_r2_c25_6 = t_r2_c25_1 + p_1_26;
  assign t_r2_c25_7 = t_r2_c25_2 + t_r2_c25_3;
  assign t_r2_c25_8 = t_r2_c25_4 + p_3_24;
  assign t_r2_c25_9 = t_r2_c25_5 + t_r2_c25_6;
  assign t_r2_c25_10 = t_r2_c25_7 + t_r2_c25_8;
  assign t_r2_c25_11 = t_r2_c25_9 + t_r2_c25_10;
  assign t_r2_c25_12 = t_r2_c25_11 + p_3_26;
  assign out_2_25 = t_r2_c25_12 >> 4;

  assign t_r2_c26_0 = p_1_26 << 1;
  assign t_r2_c26_1 = p_2_25 << 1;
  assign t_r2_c26_2 = p_2_26 << 2;
  assign t_r2_c26_3 = p_2_27 << 1;
  assign t_r2_c26_4 = p_3_26 << 1;
  assign t_r2_c26_5 = t_r2_c26_0 + p_1_25;
  assign t_r2_c26_6 = t_r2_c26_1 + p_1_27;
  assign t_r2_c26_7 = t_r2_c26_2 + t_r2_c26_3;
  assign t_r2_c26_8 = t_r2_c26_4 + p_3_25;
  assign t_r2_c26_9 = t_r2_c26_5 + t_r2_c26_6;
  assign t_r2_c26_10 = t_r2_c26_7 + t_r2_c26_8;
  assign t_r2_c26_11 = t_r2_c26_9 + t_r2_c26_10;
  assign t_r2_c26_12 = t_r2_c26_11 + p_3_27;
  assign out_2_26 = t_r2_c26_12 >> 4;

  assign t_r2_c27_0 = p_1_27 << 1;
  assign t_r2_c27_1 = p_2_26 << 1;
  assign t_r2_c27_2 = p_2_27 << 2;
  assign t_r2_c27_3 = p_2_28 << 1;
  assign t_r2_c27_4 = p_3_27 << 1;
  assign t_r2_c27_5 = t_r2_c27_0 + p_1_26;
  assign t_r2_c27_6 = t_r2_c27_1 + p_1_28;
  assign t_r2_c27_7 = t_r2_c27_2 + t_r2_c27_3;
  assign t_r2_c27_8 = t_r2_c27_4 + p_3_26;
  assign t_r2_c27_9 = t_r2_c27_5 + t_r2_c27_6;
  assign t_r2_c27_10 = t_r2_c27_7 + t_r2_c27_8;
  assign t_r2_c27_11 = t_r2_c27_9 + t_r2_c27_10;
  assign t_r2_c27_12 = t_r2_c27_11 + p_3_28;
  assign out_2_27 = t_r2_c27_12 >> 4;

  assign t_r2_c28_0 = p_1_28 << 1;
  assign t_r2_c28_1 = p_2_27 << 1;
  assign t_r2_c28_2 = p_2_28 << 2;
  assign t_r2_c28_3 = p_2_29 << 1;
  assign t_r2_c28_4 = p_3_28 << 1;
  assign t_r2_c28_5 = t_r2_c28_0 + p_1_27;
  assign t_r2_c28_6 = t_r2_c28_1 + p_1_29;
  assign t_r2_c28_7 = t_r2_c28_2 + t_r2_c28_3;
  assign t_r2_c28_8 = t_r2_c28_4 + p_3_27;
  assign t_r2_c28_9 = t_r2_c28_5 + t_r2_c28_6;
  assign t_r2_c28_10 = t_r2_c28_7 + t_r2_c28_8;
  assign t_r2_c28_11 = t_r2_c28_9 + t_r2_c28_10;
  assign t_r2_c28_12 = t_r2_c28_11 + p_3_29;
  assign out_2_28 = t_r2_c28_12 >> 4;

  assign t_r2_c29_0 = p_1_29 << 1;
  assign t_r2_c29_1 = p_2_28 << 1;
  assign t_r2_c29_2 = p_2_29 << 2;
  assign t_r2_c29_3 = p_2_30 << 1;
  assign t_r2_c29_4 = p_3_29 << 1;
  assign t_r2_c29_5 = t_r2_c29_0 + p_1_28;
  assign t_r2_c29_6 = t_r2_c29_1 + p_1_30;
  assign t_r2_c29_7 = t_r2_c29_2 + t_r2_c29_3;
  assign t_r2_c29_8 = t_r2_c29_4 + p_3_28;
  assign t_r2_c29_9 = t_r2_c29_5 + t_r2_c29_6;
  assign t_r2_c29_10 = t_r2_c29_7 + t_r2_c29_8;
  assign t_r2_c29_11 = t_r2_c29_9 + t_r2_c29_10;
  assign t_r2_c29_12 = t_r2_c29_11 + p_3_30;
  assign out_2_29 = t_r2_c29_12 >> 4;

  assign t_r2_c30_0 = p_1_30 << 1;
  assign t_r2_c30_1 = p_2_29 << 1;
  assign t_r2_c30_2 = p_2_30 << 2;
  assign t_r2_c30_3 = p_2_31 << 1;
  assign t_r2_c30_4 = p_3_30 << 1;
  assign t_r2_c30_5 = t_r2_c30_0 + p_1_29;
  assign t_r2_c30_6 = t_r2_c30_1 + p_1_31;
  assign t_r2_c30_7 = t_r2_c30_2 + t_r2_c30_3;
  assign t_r2_c30_8 = t_r2_c30_4 + p_3_29;
  assign t_r2_c30_9 = t_r2_c30_5 + t_r2_c30_6;
  assign t_r2_c30_10 = t_r2_c30_7 + t_r2_c30_8;
  assign t_r2_c30_11 = t_r2_c30_9 + t_r2_c30_10;
  assign t_r2_c30_12 = t_r2_c30_11 + p_3_31;
  assign out_2_30 = t_r2_c30_12 >> 4;

  assign t_r2_c31_0 = p_1_31 << 1;
  assign t_r2_c31_1 = p_2_30 << 1;
  assign t_r2_c31_2 = p_2_31 << 2;
  assign t_r2_c31_3 = p_2_32 << 1;
  assign t_r2_c31_4 = p_3_31 << 1;
  assign t_r2_c31_5 = t_r2_c31_0 + p_1_30;
  assign t_r2_c31_6 = t_r2_c31_1 + p_1_32;
  assign t_r2_c31_7 = t_r2_c31_2 + t_r2_c31_3;
  assign t_r2_c31_8 = t_r2_c31_4 + p_3_30;
  assign t_r2_c31_9 = t_r2_c31_5 + t_r2_c31_6;
  assign t_r2_c31_10 = t_r2_c31_7 + t_r2_c31_8;
  assign t_r2_c31_11 = t_r2_c31_9 + t_r2_c31_10;
  assign t_r2_c31_12 = t_r2_c31_11 + p_3_32;
  assign out_2_31 = t_r2_c31_12 >> 4;

  assign t_r2_c32_0 = p_1_32 << 1;
  assign t_r2_c32_1 = p_2_31 << 1;
  assign t_r2_c32_2 = p_2_32 << 2;
  assign t_r2_c32_3 = p_2_33 << 1;
  assign t_r2_c32_4 = p_3_32 << 1;
  assign t_r2_c32_5 = t_r2_c32_0 + p_1_31;
  assign t_r2_c32_6 = t_r2_c32_1 + p_1_33;
  assign t_r2_c32_7 = t_r2_c32_2 + t_r2_c32_3;
  assign t_r2_c32_8 = t_r2_c32_4 + p_3_31;
  assign t_r2_c32_9 = t_r2_c32_5 + t_r2_c32_6;
  assign t_r2_c32_10 = t_r2_c32_7 + t_r2_c32_8;
  assign t_r2_c32_11 = t_r2_c32_9 + t_r2_c32_10;
  assign t_r2_c32_12 = t_r2_c32_11 + p_3_33;
  assign out_2_32 = t_r2_c32_12 >> 4;

  assign t_r2_c33_0 = p_1_33 << 1;
  assign t_r2_c33_1 = p_2_32 << 1;
  assign t_r2_c33_2 = p_2_33 << 2;
  assign t_r2_c33_3 = p_2_34 << 1;
  assign t_r2_c33_4 = p_3_33 << 1;
  assign t_r2_c33_5 = t_r2_c33_0 + p_1_32;
  assign t_r2_c33_6 = t_r2_c33_1 + p_1_34;
  assign t_r2_c33_7 = t_r2_c33_2 + t_r2_c33_3;
  assign t_r2_c33_8 = t_r2_c33_4 + p_3_32;
  assign t_r2_c33_9 = t_r2_c33_5 + t_r2_c33_6;
  assign t_r2_c33_10 = t_r2_c33_7 + t_r2_c33_8;
  assign t_r2_c33_11 = t_r2_c33_9 + t_r2_c33_10;
  assign t_r2_c33_12 = t_r2_c33_11 + p_3_34;
  assign out_2_33 = t_r2_c33_12 >> 4;

  assign t_r2_c34_0 = p_1_34 << 1;
  assign t_r2_c34_1 = p_2_33 << 1;
  assign t_r2_c34_2 = p_2_34 << 2;
  assign t_r2_c34_3 = p_2_35 << 1;
  assign t_r2_c34_4 = p_3_34 << 1;
  assign t_r2_c34_5 = t_r2_c34_0 + p_1_33;
  assign t_r2_c34_6 = t_r2_c34_1 + p_1_35;
  assign t_r2_c34_7 = t_r2_c34_2 + t_r2_c34_3;
  assign t_r2_c34_8 = t_r2_c34_4 + p_3_33;
  assign t_r2_c34_9 = t_r2_c34_5 + t_r2_c34_6;
  assign t_r2_c34_10 = t_r2_c34_7 + t_r2_c34_8;
  assign t_r2_c34_11 = t_r2_c34_9 + t_r2_c34_10;
  assign t_r2_c34_12 = t_r2_c34_11 + p_3_35;
  assign out_2_34 = t_r2_c34_12 >> 4;

  assign t_r2_c35_0 = p_1_35 << 1;
  assign t_r2_c35_1 = p_2_34 << 1;
  assign t_r2_c35_2 = p_2_35 << 2;
  assign t_r2_c35_3 = p_2_36 << 1;
  assign t_r2_c35_4 = p_3_35 << 1;
  assign t_r2_c35_5 = t_r2_c35_0 + p_1_34;
  assign t_r2_c35_6 = t_r2_c35_1 + p_1_36;
  assign t_r2_c35_7 = t_r2_c35_2 + t_r2_c35_3;
  assign t_r2_c35_8 = t_r2_c35_4 + p_3_34;
  assign t_r2_c35_9 = t_r2_c35_5 + t_r2_c35_6;
  assign t_r2_c35_10 = t_r2_c35_7 + t_r2_c35_8;
  assign t_r2_c35_11 = t_r2_c35_9 + t_r2_c35_10;
  assign t_r2_c35_12 = t_r2_c35_11 + p_3_36;
  assign out_2_35 = t_r2_c35_12 >> 4;

  assign t_r2_c36_0 = p_1_36 << 1;
  assign t_r2_c36_1 = p_2_35 << 1;
  assign t_r2_c36_2 = p_2_36 << 2;
  assign t_r2_c36_3 = p_2_37 << 1;
  assign t_r2_c36_4 = p_3_36 << 1;
  assign t_r2_c36_5 = t_r2_c36_0 + p_1_35;
  assign t_r2_c36_6 = t_r2_c36_1 + p_1_37;
  assign t_r2_c36_7 = t_r2_c36_2 + t_r2_c36_3;
  assign t_r2_c36_8 = t_r2_c36_4 + p_3_35;
  assign t_r2_c36_9 = t_r2_c36_5 + t_r2_c36_6;
  assign t_r2_c36_10 = t_r2_c36_7 + t_r2_c36_8;
  assign t_r2_c36_11 = t_r2_c36_9 + t_r2_c36_10;
  assign t_r2_c36_12 = t_r2_c36_11 + p_3_37;
  assign out_2_36 = t_r2_c36_12 >> 4;

  assign t_r2_c37_0 = p_1_37 << 1;
  assign t_r2_c37_1 = p_2_36 << 1;
  assign t_r2_c37_2 = p_2_37 << 2;
  assign t_r2_c37_3 = p_2_38 << 1;
  assign t_r2_c37_4 = p_3_37 << 1;
  assign t_r2_c37_5 = t_r2_c37_0 + p_1_36;
  assign t_r2_c37_6 = t_r2_c37_1 + p_1_38;
  assign t_r2_c37_7 = t_r2_c37_2 + t_r2_c37_3;
  assign t_r2_c37_8 = t_r2_c37_4 + p_3_36;
  assign t_r2_c37_9 = t_r2_c37_5 + t_r2_c37_6;
  assign t_r2_c37_10 = t_r2_c37_7 + t_r2_c37_8;
  assign t_r2_c37_11 = t_r2_c37_9 + t_r2_c37_10;
  assign t_r2_c37_12 = t_r2_c37_11 + p_3_38;
  assign out_2_37 = t_r2_c37_12 >> 4;

  assign t_r2_c38_0 = p_1_38 << 1;
  assign t_r2_c38_1 = p_2_37 << 1;
  assign t_r2_c38_2 = p_2_38 << 2;
  assign t_r2_c38_3 = p_2_39 << 1;
  assign t_r2_c38_4 = p_3_38 << 1;
  assign t_r2_c38_5 = t_r2_c38_0 + p_1_37;
  assign t_r2_c38_6 = t_r2_c38_1 + p_1_39;
  assign t_r2_c38_7 = t_r2_c38_2 + t_r2_c38_3;
  assign t_r2_c38_8 = t_r2_c38_4 + p_3_37;
  assign t_r2_c38_9 = t_r2_c38_5 + t_r2_c38_6;
  assign t_r2_c38_10 = t_r2_c38_7 + t_r2_c38_8;
  assign t_r2_c38_11 = t_r2_c38_9 + t_r2_c38_10;
  assign t_r2_c38_12 = t_r2_c38_11 + p_3_39;
  assign out_2_38 = t_r2_c38_12 >> 4;

  assign t_r2_c39_0 = p_1_39 << 1;
  assign t_r2_c39_1 = p_2_38 << 1;
  assign t_r2_c39_2 = p_2_39 << 2;
  assign t_r2_c39_3 = p_2_40 << 1;
  assign t_r2_c39_4 = p_3_39 << 1;
  assign t_r2_c39_5 = t_r2_c39_0 + p_1_38;
  assign t_r2_c39_6 = t_r2_c39_1 + p_1_40;
  assign t_r2_c39_7 = t_r2_c39_2 + t_r2_c39_3;
  assign t_r2_c39_8 = t_r2_c39_4 + p_3_38;
  assign t_r2_c39_9 = t_r2_c39_5 + t_r2_c39_6;
  assign t_r2_c39_10 = t_r2_c39_7 + t_r2_c39_8;
  assign t_r2_c39_11 = t_r2_c39_9 + t_r2_c39_10;
  assign t_r2_c39_12 = t_r2_c39_11 + p_3_40;
  assign out_2_39 = t_r2_c39_12 >> 4;

  assign t_r2_c40_0 = p_1_40 << 1;
  assign t_r2_c40_1 = p_2_39 << 1;
  assign t_r2_c40_2 = p_2_40 << 2;
  assign t_r2_c40_3 = p_2_41 << 1;
  assign t_r2_c40_4 = p_3_40 << 1;
  assign t_r2_c40_5 = t_r2_c40_0 + p_1_39;
  assign t_r2_c40_6 = t_r2_c40_1 + p_1_41;
  assign t_r2_c40_7 = t_r2_c40_2 + t_r2_c40_3;
  assign t_r2_c40_8 = t_r2_c40_4 + p_3_39;
  assign t_r2_c40_9 = t_r2_c40_5 + t_r2_c40_6;
  assign t_r2_c40_10 = t_r2_c40_7 + t_r2_c40_8;
  assign t_r2_c40_11 = t_r2_c40_9 + t_r2_c40_10;
  assign t_r2_c40_12 = t_r2_c40_11 + p_3_41;
  assign out_2_40 = t_r2_c40_12 >> 4;

  assign t_r2_c41_0 = p_1_41 << 1;
  assign t_r2_c41_1 = p_2_40 << 1;
  assign t_r2_c41_2 = p_2_41 << 2;
  assign t_r2_c41_3 = p_2_42 << 1;
  assign t_r2_c41_4 = p_3_41 << 1;
  assign t_r2_c41_5 = t_r2_c41_0 + p_1_40;
  assign t_r2_c41_6 = t_r2_c41_1 + p_1_42;
  assign t_r2_c41_7 = t_r2_c41_2 + t_r2_c41_3;
  assign t_r2_c41_8 = t_r2_c41_4 + p_3_40;
  assign t_r2_c41_9 = t_r2_c41_5 + t_r2_c41_6;
  assign t_r2_c41_10 = t_r2_c41_7 + t_r2_c41_8;
  assign t_r2_c41_11 = t_r2_c41_9 + t_r2_c41_10;
  assign t_r2_c41_12 = t_r2_c41_11 + p_3_42;
  assign out_2_41 = t_r2_c41_12 >> 4;

  assign t_r2_c42_0 = p_1_42 << 1;
  assign t_r2_c42_1 = p_2_41 << 1;
  assign t_r2_c42_2 = p_2_42 << 2;
  assign t_r2_c42_3 = p_2_43 << 1;
  assign t_r2_c42_4 = p_3_42 << 1;
  assign t_r2_c42_5 = t_r2_c42_0 + p_1_41;
  assign t_r2_c42_6 = t_r2_c42_1 + p_1_43;
  assign t_r2_c42_7 = t_r2_c42_2 + t_r2_c42_3;
  assign t_r2_c42_8 = t_r2_c42_4 + p_3_41;
  assign t_r2_c42_9 = t_r2_c42_5 + t_r2_c42_6;
  assign t_r2_c42_10 = t_r2_c42_7 + t_r2_c42_8;
  assign t_r2_c42_11 = t_r2_c42_9 + t_r2_c42_10;
  assign t_r2_c42_12 = t_r2_c42_11 + p_3_43;
  assign out_2_42 = t_r2_c42_12 >> 4;

  assign t_r2_c43_0 = p_1_43 << 1;
  assign t_r2_c43_1 = p_2_42 << 1;
  assign t_r2_c43_2 = p_2_43 << 2;
  assign t_r2_c43_3 = p_2_44 << 1;
  assign t_r2_c43_4 = p_3_43 << 1;
  assign t_r2_c43_5 = t_r2_c43_0 + p_1_42;
  assign t_r2_c43_6 = t_r2_c43_1 + p_1_44;
  assign t_r2_c43_7 = t_r2_c43_2 + t_r2_c43_3;
  assign t_r2_c43_8 = t_r2_c43_4 + p_3_42;
  assign t_r2_c43_9 = t_r2_c43_5 + t_r2_c43_6;
  assign t_r2_c43_10 = t_r2_c43_7 + t_r2_c43_8;
  assign t_r2_c43_11 = t_r2_c43_9 + t_r2_c43_10;
  assign t_r2_c43_12 = t_r2_c43_11 + p_3_44;
  assign out_2_43 = t_r2_c43_12 >> 4;

  assign t_r2_c44_0 = p_1_44 << 1;
  assign t_r2_c44_1 = p_2_43 << 1;
  assign t_r2_c44_2 = p_2_44 << 2;
  assign t_r2_c44_3 = p_2_45 << 1;
  assign t_r2_c44_4 = p_3_44 << 1;
  assign t_r2_c44_5 = t_r2_c44_0 + p_1_43;
  assign t_r2_c44_6 = t_r2_c44_1 + p_1_45;
  assign t_r2_c44_7 = t_r2_c44_2 + t_r2_c44_3;
  assign t_r2_c44_8 = t_r2_c44_4 + p_3_43;
  assign t_r2_c44_9 = t_r2_c44_5 + t_r2_c44_6;
  assign t_r2_c44_10 = t_r2_c44_7 + t_r2_c44_8;
  assign t_r2_c44_11 = t_r2_c44_9 + t_r2_c44_10;
  assign t_r2_c44_12 = t_r2_c44_11 + p_3_45;
  assign out_2_44 = t_r2_c44_12 >> 4;

  assign t_r2_c45_0 = p_1_45 << 1;
  assign t_r2_c45_1 = p_2_44 << 1;
  assign t_r2_c45_2 = p_2_45 << 2;
  assign t_r2_c45_3 = p_2_46 << 1;
  assign t_r2_c45_4 = p_3_45 << 1;
  assign t_r2_c45_5 = t_r2_c45_0 + p_1_44;
  assign t_r2_c45_6 = t_r2_c45_1 + p_1_46;
  assign t_r2_c45_7 = t_r2_c45_2 + t_r2_c45_3;
  assign t_r2_c45_8 = t_r2_c45_4 + p_3_44;
  assign t_r2_c45_9 = t_r2_c45_5 + t_r2_c45_6;
  assign t_r2_c45_10 = t_r2_c45_7 + t_r2_c45_8;
  assign t_r2_c45_11 = t_r2_c45_9 + t_r2_c45_10;
  assign t_r2_c45_12 = t_r2_c45_11 + p_3_46;
  assign out_2_45 = t_r2_c45_12 >> 4;

  assign t_r2_c46_0 = p_1_46 << 1;
  assign t_r2_c46_1 = p_2_45 << 1;
  assign t_r2_c46_2 = p_2_46 << 2;
  assign t_r2_c46_3 = p_2_47 << 1;
  assign t_r2_c46_4 = p_3_46 << 1;
  assign t_r2_c46_5 = t_r2_c46_0 + p_1_45;
  assign t_r2_c46_6 = t_r2_c46_1 + p_1_47;
  assign t_r2_c46_7 = t_r2_c46_2 + t_r2_c46_3;
  assign t_r2_c46_8 = t_r2_c46_4 + p_3_45;
  assign t_r2_c46_9 = t_r2_c46_5 + t_r2_c46_6;
  assign t_r2_c46_10 = t_r2_c46_7 + t_r2_c46_8;
  assign t_r2_c46_11 = t_r2_c46_9 + t_r2_c46_10;
  assign t_r2_c46_12 = t_r2_c46_11 + p_3_47;
  assign out_2_46 = t_r2_c46_12 >> 4;

  assign t_r2_c47_0 = p_1_47 << 1;
  assign t_r2_c47_1 = p_2_46 << 1;
  assign t_r2_c47_2 = p_2_47 << 2;
  assign t_r2_c47_3 = p_2_48 << 1;
  assign t_r2_c47_4 = p_3_47 << 1;
  assign t_r2_c47_5 = t_r2_c47_0 + p_1_46;
  assign t_r2_c47_6 = t_r2_c47_1 + p_1_48;
  assign t_r2_c47_7 = t_r2_c47_2 + t_r2_c47_3;
  assign t_r2_c47_8 = t_r2_c47_4 + p_3_46;
  assign t_r2_c47_9 = t_r2_c47_5 + t_r2_c47_6;
  assign t_r2_c47_10 = t_r2_c47_7 + t_r2_c47_8;
  assign t_r2_c47_11 = t_r2_c47_9 + t_r2_c47_10;
  assign t_r2_c47_12 = t_r2_c47_11 + p_3_48;
  assign out_2_47 = t_r2_c47_12 >> 4;

  assign t_r2_c48_0 = p_1_48 << 1;
  assign t_r2_c48_1 = p_2_47 << 1;
  assign t_r2_c48_2 = p_2_48 << 2;
  assign t_r2_c48_3 = p_2_49 << 1;
  assign t_r2_c48_4 = p_3_48 << 1;
  assign t_r2_c48_5 = t_r2_c48_0 + p_1_47;
  assign t_r2_c48_6 = t_r2_c48_1 + p_1_49;
  assign t_r2_c48_7 = t_r2_c48_2 + t_r2_c48_3;
  assign t_r2_c48_8 = t_r2_c48_4 + p_3_47;
  assign t_r2_c48_9 = t_r2_c48_5 + t_r2_c48_6;
  assign t_r2_c48_10 = t_r2_c48_7 + t_r2_c48_8;
  assign t_r2_c48_11 = t_r2_c48_9 + t_r2_c48_10;
  assign t_r2_c48_12 = t_r2_c48_11 + p_3_49;
  assign out_2_48 = t_r2_c48_12 >> 4;

  assign t_r2_c49_0 = p_1_49 << 1;
  assign t_r2_c49_1 = p_2_48 << 1;
  assign t_r2_c49_2 = p_2_49 << 2;
  assign t_r2_c49_3 = p_2_50 << 1;
  assign t_r2_c49_4 = p_3_49 << 1;
  assign t_r2_c49_5 = t_r2_c49_0 + p_1_48;
  assign t_r2_c49_6 = t_r2_c49_1 + p_1_50;
  assign t_r2_c49_7 = t_r2_c49_2 + t_r2_c49_3;
  assign t_r2_c49_8 = t_r2_c49_4 + p_3_48;
  assign t_r2_c49_9 = t_r2_c49_5 + t_r2_c49_6;
  assign t_r2_c49_10 = t_r2_c49_7 + t_r2_c49_8;
  assign t_r2_c49_11 = t_r2_c49_9 + t_r2_c49_10;
  assign t_r2_c49_12 = t_r2_c49_11 + p_3_50;
  assign out_2_49 = t_r2_c49_12 >> 4;

  assign t_r2_c50_0 = p_1_50 << 1;
  assign t_r2_c50_1 = p_2_49 << 1;
  assign t_r2_c50_2 = p_2_50 << 2;
  assign t_r2_c50_3 = p_2_51 << 1;
  assign t_r2_c50_4 = p_3_50 << 1;
  assign t_r2_c50_5 = t_r2_c50_0 + p_1_49;
  assign t_r2_c50_6 = t_r2_c50_1 + p_1_51;
  assign t_r2_c50_7 = t_r2_c50_2 + t_r2_c50_3;
  assign t_r2_c50_8 = t_r2_c50_4 + p_3_49;
  assign t_r2_c50_9 = t_r2_c50_5 + t_r2_c50_6;
  assign t_r2_c50_10 = t_r2_c50_7 + t_r2_c50_8;
  assign t_r2_c50_11 = t_r2_c50_9 + t_r2_c50_10;
  assign t_r2_c50_12 = t_r2_c50_11 + p_3_51;
  assign out_2_50 = t_r2_c50_12 >> 4;

  assign t_r2_c51_0 = p_1_51 << 1;
  assign t_r2_c51_1 = p_2_50 << 1;
  assign t_r2_c51_2 = p_2_51 << 2;
  assign t_r2_c51_3 = p_2_52 << 1;
  assign t_r2_c51_4 = p_3_51 << 1;
  assign t_r2_c51_5 = t_r2_c51_0 + p_1_50;
  assign t_r2_c51_6 = t_r2_c51_1 + p_1_52;
  assign t_r2_c51_7 = t_r2_c51_2 + t_r2_c51_3;
  assign t_r2_c51_8 = t_r2_c51_4 + p_3_50;
  assign t_r2_c51_9 = t_r2_c51_5 + t_r2_c51_6;
  assign t_r2_c51_10 = t_r2_c51_7 + t_r2_c51_8;
  assign t_r2_c51_11 = t_r2_c51_9 + t_r2_c51_10;
  assign t_r2_c51_12 = t_r2_c51_11 + p_3_52;
  assign out_2_51 = t_r2_c51_12 >> 4;

  assign t_r2_c52_0 = p_1_52 << 1;
  assign t_r2_c52_1 = p_2_51 << 1;
  assign t_r2_c52_2 = p_2_52 << 2;
  assign t_r2_c52_3 = p_2_53 << 1;
  assign t_r2_c52_4 = p_3_52 << 1;
  assign t_r2_c52_5 = t_r2_c52_0 + p_1_51;
  assign t_r2_c52_6 = t_r2_c52_1 + p_1_53;
  assign t_r2_c52_7 = t_r2_c52_2 + t_r2_c52_3;
  assign t_r2_c52_8 = t_r2_c52_4 + p_3_51;
  assign t_r2_c52_9 = t_r2_c52_5 + t_r2_c52_6;
  assign t_r2_c52_10 = t_r2_c52_7 + t_r2_c52_8;
  assign t_r2_c52_11 = t_r2_c52_9 + t_r2_c52_10;
  assign t_r2_c52_12 = t_r2_c52_11 + p_3_53;
  assign out_2_52 = t_r2_c52_12 >> 4;

  assign t_r2_c53_0 = p_1_53 << 1;
  assign t_r2_c53_1 = p_2_52 << 1;
  assign t_r2_c53_2 = p_2_53 << 2;
  assign t_r2_c53_3 = p_2_54 << 1;
  assign t_r2_c53_4 = p_3_53 << 1;
  assign t_r2_c53_5 = t_r2_c53_0 + p_1_52;
  assign t_r2_c53_6 = t_r2_c53_1 + p_1_54;
  assign t_r2_c53_7 = t_r2_c53_2 + t_r2_c53_3;
  assign t_r2_c53_8 = t_r2_c53_4 + p_3_52;
  assign t_r2_c53_9 = t_r2_c53_5 + t_r2_c53_6;
  assign t_r2_c53_10 = t_r2_c53_7 + t_r2_c53_8;
  assign t_r2_c53_11 = t_r2_c53_9 + t_r2_c53_10;
  assign t_r2_c53_12 = t_r2_c53_11 + p_3_54;
  assign out_2_53 = t_r2_c53_12 >> 4;

  assign t_r2_c54_0 = p_1_54 << 1;
  assign t_r2_c54_1 = p_2_53 << 1;
  assign t_r2_c54_2 = p_2_54 << 2;
  assign t_r2_c54_3 = p_2_55 << 1;
  assign t_r2_c54_4 = p_3_54 << 1;
  assign t_r2_c54_5 = t_r2_c54_0 + p_1_53;
  assign t_r2_c54_6 = t_r2_c54_1 + p_1_55;
  assign t_r2_c54_7 = t_r2_c54_2 + t_r2_c54_3;
  assign t_r2_c54_8 = t_r2_c54_4 + p_3_53;
  assign t_r2_c54_9 = t_r2_c54_5 + t_r2_c54_6;
  assign t_r2_c54_10 = t_r2_c54_7 + t_r2_c54_8;
  assign t_r2_c54_11 = t_r2_c54_9 + t_r2_c54_10;
  assign t_r2_c54_12 = t_r2_c54_11 + p_3_55;
  assign out_2_54 = t_r2_c54_12 >> 4;

  assign t_r2_c55_0 = p_1_55 << 1;
  assign t_r2_c55_1 = p_2_54 << 1;
  assign t_r2_c55_2 = p_2_55 << 2;
  assign t_r2_c55_3 = p_2_56 << 1;
  assign t_r2_c55_4 = p_3_55 << 1;
  assign t_r2_c55_5 = t_r2_c55_0 + p_1_54;
  assign t_r2_c55_6 = t_r2_c55_1 + p_1_56;
  assign t_r2_c55_7 = t_r2_c55_2 + t_r2_c55_3;
  assign t_r2_c55_8 = t_r2_c55_4 + p_3_54;
  assign t_r2_c55_9 = t_r2_c55_5 + t_r2_c55_6;
  assign t_r2_c55_10 = t_r2_c55_7 + t_r2_c55_8;
  assign t_r2_c55_11 = t_r2_c55_9 + t_r2_c55_10;
  assign t_r2_c55_12 = t_r2_c55_11 + p_3_56;
  assign out_2_55 = t_r2_c55_12 >> 4;

  assign t_r2_c56_0 = p_1_56 << 1;
  assign t_r2_c56_1 = p_2_55 << 1;
  assign t_r2_c56_2 = p_2_56 << 2;
  assign t_r2_c56_3 = p_2_57 << 1;
  assign t_r2_c56_4 = p_3_56 << 1;
  assign t_r2_c56_5 = t_r2_c56_0 + p_1_55;
  assign t_r2_c56_6 = t_r2_c56_1 + p_1_57;
  assign t_r2_c56_7 = t_r2_c56_2 + t_r2_c56_3;
  assign t_r2_c56_8 = t_r2_c56_4 + p_3_55;
  assign t_r2_c56_9 = t_r2_c56_5 + t_r2_c56_6;
  assign t_r2_c56_10 = t_r2_c56_7 + t_r2_c56_8;
  assign t_r2_c56_11 = t_r2_c56_9 + t_r2_c56_10;
  assign t_r2_c56_12 = t_r2_c56_11 + p_3_57;
  assign out_2_56 = t_r2_c56_12 >> 4;

  assign t_r2_c57_0 = p_1_57 << 1;
  assign t_r2_c57_1 = p_2_56 << 1;
  assign t_r2_c57_2 = p_2_57 << 2;
  assign t_r2_c57_3 = p_2_58 << 1;
  assign t_r2_c57_4 = p_3_57 << 1;
  assign t_r2_c57_5 = t_r2_c57_0 + p_1_56;
  assign t_r2_c57_6 = t_r2_c57_1 + p_1_58;
  assign t_r2_c57_7 = t_r2_c57_2 + t_r2_c57_3;
  assign t_r2_c57_8 = t_r2_c57_4 + p_3_56;
  assign t_r2_c57_9 = t_r2_c57_5 + t_r2_c57_6;
  assign t_r2_c57_10 = t_r2_c57_7 + t_r2_c57_8;
  assign t_r2_c57_11 = t_r2_c57_9 + t_r2_c57_10;
  assign t_r2_c57_12 = t_r2_c57_11 + p_3_58;
  assign out_2_57 = t_r2_c57_12 >> 4;

  assign t_r2_c58_0 = p_1_58 << 1;
  assign t_r2_c58_1 = p_2_57 << 1;
  assign t_r2_c58_2 = p_2_58 << 2;
  assign t_r2_c58_3 = p_2_59 << 1;
  assign t_r2_c58_4 = p_3_58 << 1;
  assign t_r2_c58_5 = t_r2_c58_0 + p_1_57;
  assign t_r2_c58_6 = t_r2_c58_1 + p_1_59;
  assign t_r2_c58_7 = t_r2_c58_2 + t_r2_c58_3;
  assign t_r2_c58_8 = t_r2_c58_4 + p_3_57;
  assign t_r2_c58_9 = t_r2_c58_5 + t_r2_c58_6;
  assign t_r2_c58_10 = t_r2_c58_7 + t_r2_c58_8;
  assign t_r2_c58_11 = t_r2_c58_9 + t_r2_c58_10;
  assign t_r2_c58_12 = t_r2_c58_11 + p_3_59;
  assign out_2_58 = t_r2_c58_12 >> 4;

  assign t_r2_c59_0 = p_1_59 << 1;
  assign t_r2_c59_1 = p_2_58 << 1;
  assign t_r2_c59_2 = p_2_59 << 2;
  assign t_r2_c59_3 = p_2_60 << 1;
  assign t_r2_c59_4 = p_3_59 << 1;
  assign t_r2_c59_5 = t_r2_c59_0 + p_1_58;
  assign t_r2_c59_6 = t_r2_c59_1 + p_1_60;
  assign t_r2_c59_7 = t_r2_c59_2 + t_r2_c59_3;
  assign t_r2_c59_8 = t_r2_c59_4 + p_3_58;
  assign t_r2_c59_9 = t_r2_c59_5 + t_r2_c59_6;
  assign t_r2_c59_10 = t_r2_c59_7 + t_r2_c59_8;
  assign t_r2_c59_11 = t_r2_c59_9 + t_r2_c59_10;
  assign t_r2_c59_12 = t_r2_c59_11 + p_3_60;
  assign out_2_59 = t_r2_c59_12 >> 4;

  assign t_r2_c60_0 = p_1_60 << 1;
  assign t_r2_c60_1 = p_2_59 << 1;
  assign t_r2_c60_2 = p_2_60 << 2;
  assign t_r2_c60_3 = p_2_61 << 1;
  assign t_r2_c60_4 = p_3_60 << 1;
  assign t_r2_c60_5 = t_r2_c60_0 + p_1_59;
  assign t_r2_c60_6 = t_r2_c60_1 + p_1_61;
  assign t_r2_c60_7 = t_r2_c60_2 + t_r2_c60_3;
  assign t_r2_c60_8 = t_r2_c60_4 + p_3_59;
  assign t_r2_c60_9 = t_r2_c60_5 + t_r2_c60_6;
  assign t_r2_c60_10 = t_r2_c60_7 + t_r2_c60_8;
  assign t_r2_c60_11 = t_r2_c60_9 + t_r2_c60_10;
  assign t_r2_c60_12 = t_r2_c60_11 + p_3_61;
  assign out_2_60 = t_r2_c60_12 >> 4;

  assign t_r2_c61_0 = p_1_61 << 1;
  assign t_r2_c61_1 = p_2_60 << 1;
  assign t_r2_c61_2 = p_2_61 << 2;
  assign t_r2_c61_3 = p_2_62 << 1;
  assign t_r2_c61_4 = p_3_61 << 1;
  assign t_r2_c61_5 = t_r2_c61_0 + p_1_60;
  assign t_r2_c61_6 = t_r2_c61_1 + p_1_62;
  assign t_r2_c61_7 = t_r2_c61_2 + t_r2_c61_3;
  assign t_r2_c61_8 = t_r2_c61_4 + p_3_60;
  assign t_r2_c61_9 = t_r2_c61_5 + t_r2_c61_6;
  assign t_r2_c61_10 = t_r2_c61_7 + t_r2_c61_8;
  assign t_r2_c61_11 = t_r2_c61_9 + t_r2_c61_10;
  assign t_r2_c61_12 = t_r2_c61_11 + p_3_62;
  assign out_2_61 = t_r2_c61_12 >> 4;

  assign t_r2_c62_0 = p_1_62 << 1;
  assign t_r2_c62_1 = p_2_61 << 1;
  assign t_r2_c62_2 = p_2_62 << 2;
  assign t_r2_c62_3 = p_2_63 << 1;
  assign t_r2_c62_4 = p_3_62 << 1;
  assign t_r2_c62_5 = t_r2_c62_0 + p_1_61;
  assign t_r2_c62_6 = t_r2_c62_1 + p_1_63;
  assign t_r2_c62_7 = t_r2_c62_2 + t_r2_c62_3;
  assign t_r2_c62_8 = t_r2_c62_4 + p_3_61;
  assign t_r2_c62_9 = t_r2_c62_5 + t_r2_c62_6;
  assign t_r2_c62_10 = t_r2_c62_7 + t_r2_c62_8;
  assign t_r2_c62_11 = t_r2_c62_9 + t_r2_c62_10;
  assign t_r2_c62_12 = t_r2_c62_11 + p_3_63;
  assign out_2_62 = t_r2_c62_12 >> 4;

  assign t_r2_c63_0 = p_1_63 << 1;
  assign t_r2_c63_1 = p_2_62 << 1;
  assign t_r2_c63_2 = p_2_63 << 2;
  assign t_r2_c63_3 = p_2_64 << 1;
  assign t_r2_c63_4 = p_3_63 << 1;
  assign t_r2_c63_5 = t_r2_c63_0 + p_1_62;
  assign t_r2_c63_6 = t_r2_c63_1 + p_1_64;
  assign t_r2_c63_7 = t_r2_c63_2 + t_r2_c63_3;
  assign t_r2_c63_8 = t_r2_c63_4 + p_3_62;
  assign t_r2_c63_9 = t_r2_c63_5 + t_r2_c63_6;
  assign t_r2_c63_10 = t_r2_c63_7 + t_r2_c63_8;
  assign t_r2_c63_11 = t_r2_c63_9 + t_r2_c63_10;
  assign t_r2_c63_12 = t_r2_c63_11 + p_3_64;
  assign out_2_63 = t_r2_c63_12 >> 4;

  assign t_r2_c64_0 = p_1_64 << 1;
  assign t_r2_c64_1 = p_2_63 << 1;
  assign t_r2_c64_2 = p_2_64 << 2;
  assign t_r2_c64_3 = p_2_65 << 1;
  assign t_r2_c64_4 = p_3_64 << 1;
  assign t_r2_c64_5 = t_r2_c64_0 + p_1_63;
  assign t_r2_c64_6 = t_r2_c64_1 + p_1_65;
  assign t_r2_c64_7 = t_r2_c64_2 + t_r2_c64_3;
  assign t_r2_c64_8 = t_r2_c64_4 + p_3_63;
  assign t_r2_c64_9 = t_r2_c64_5 + t_r2_c64_6;
  assign t_r2_c64_10 = t_r2_c64_7 + t_r2_c64_8;
  assign t_r2_c64_11 = t_r2_c64_9 + t_r2_c64_10;
  assign t_r2_c64_12 = t_r2_c64_11 + p_3_65;
  assign out_2_64 = t_r2_c64_12 >> 4;

  assign t_r3_c1_0 = p_2_1 << 1;
  assign t_r3_c1_1 = p_3_0 << 1;
  assign t_r3_c1_2 = p_3_1 << 2;
  assign t_r3_c1_3 = p_3_2 << 1;
  assign t_r3_c1_4 = p_4_1 << 1;
  assign t_r3_c1_5 = t_r3_c1_0 + p_2_0;
  assign t_r3_c1_6 = t_r3_c1_1 + p_2_2;
  assign t_r3_c1_7 = t_r3_c1_2 + t_r3_c1_3;
  assign t_r3_c1_8 = t_r3_c1_4 + p_4_0;
  assign t_r3_c1_9 = t_r3_c1_5 + t_r3_c1_6;
  assign t_r3_c1_10 = t_r3_c1_7 + t_r3_c1_8;
  assign t_r3_c1_11 = t_r3_c1_9 + t_r3_c1_10;
  assign t_r3_c1_12 = t_r3_c1_11 + p_4_2;
  assign out_3_1 = t_r3_c1_12 >> 4;

  assign t_r3_c2_0 = p_2_2 << 1;
  assign t_r3_c2_1 = p_3_1 << 1;
  assign t_r3_c2_2 = p_3_2 << 2;
  assign t_r3_c2_3 = p_3_3 << 1;
  assign t_r3_c2_4 = p_4_2 << 1;
  assign t_r3_c2_5 = t_r3_c2_0 + p_2_1;
  assign t_r3_c2_6 = t_r3_c2_1 + p_2_3;
  assign t_r3_c2_7 = t_r3_c2_2 + t_r3_c2_3;
  assign t_r3_c2_8 = t_r3_c2_4 + p_4_1;
  assign t_r3_c2_9 = t_r3_c2_5 + t_r3_c2_6;
  assign t_r3_c2_10 = t_r3_c2_7 + t_r3_c2_8;
  assign t_r3_c2_11 = t_r3_c2_9 + t_r3_c2_10;
  assign t_r3_c2_12 = t_r3_c2_11 + p_4_3;
  assign out_3_2 = t_r3_c2_12 >> 4;

  assign t_r3_c3_0 = p_2_3 << 1;
  assign t_r3_c3_1 = p_3_2 << 1;
  assign t_r3_c3_2 = p_3_3 << 2;
  assign t_r3_c3_3 = p_3_4 << 1;
  assign t_r3_c3_4 = p_4_3 << 1;
  assign t_r3_c3_5 = t_r3_c3_0 + p_2_2;
  assign t_r3_c3_6 = t_r3_c3_1 + p_2_4;
  assign t_r3_c3_7 = t_r3_c3_2 + t_r3_c3_3;
  assign t_r3_c3_8 = t_r3_c3_4 + p_4_2;
  assign t_r3_c3_9 = t_r3_c3_5 + t_r3_c3_6;
  assign t_r3_c3_10 = t_r3_c3_7 + t_r3_c3_8;
  assign t_r3_c3_11 = t_r3_c3_9 + t_r3_c3_10;
  assign t_r3_c3_12 = t_r3_c3_11 + p_4_4;
  assign out_3_3 = t_r3_c3_12 >> 4;

  assign t_r3_c4_0 = p_2_4 << 1;
  assign t_r3_c4_1 = p_3_3 << 1;
  assign t_r3_c4_2 = p_3_4 << 2;
  assign t_r3_c4_3 = p_3_5 << 1;
  assign t_r3_c4_4 = p_4_4 << 1;
  assign t_r3_c4_5 = t_r3_c4_0 + p_2_3;
  assign t_r3_c4_6 = t_r3_c4_1 + p_2_5;
  assign t_r3_c4_7 = t_r3_c4_2 + t_r3_c4_3;
  assign t_r3_c4_8 = t_r3_c4_4 + p_4_3;
  assign t_r3_c4_9 = t_r3_c4_5 + t_r3_c4_6;
  assign t_r3_c4_10 = t_r3_c4_7 + t_r3_c4_8;
  assign t_r3_c4_11 = t_r3_c4_9 + t_r3_c4_10;
  assign t_r3_c4_12 = t_r3_c4_11 + p_4_5;
  assign out_3_4 = t_r3_c4_12 >> 4;

  assign t_r3_c5_0 = p_2_5 << 1;
  assign t_r3_c5_1 = p_3_4 << 1;
  assign t_r3_c5_2 = p_3_5 << 2;
  assign t_r3_c5_3 = p_3_6 << 1;
  assign t_r3_c5_4 = p_4_5 << 1;
  assign t_r3_c5_5 = t_r3_c5_0 + p_2_4;
  assign t_r3_c5_6 = t_r3_c5_1 + p_2_6;
  assign t_r3_c5_7 = t_r3_c5_2 + t_r3_c5_3;
  assign t_r3_c5_8 = t_r3_c5_4 + p_4_4;
  assign t_r3_c5_9 = t_r3_c5_5 + t_r3_c5_6;
  assign t_r3_c5_10 = t_r3_c5_7 + t_r3_c5_8;
  assign t_r3_c5_11 = t_r3_c5_9 + t_r3_c5_10;
  assign t_r3_c5_12 = t_r3_c5_11 + p_4_6;
  assign out_3_5 = t_r3_c5_12 >> 4;

  assign t_r3_c6_0 = p_2_6 << 1;
  assign t_r3_c6_1 = p_3_5 << 1;
  assign t_r3_c6_2 = p_3_6 << 2;
  assign t_r3_c6_3 = p_3_7 << 1;
  assign t_r3_c6_4 = p_4_6 << 1;
  assign t_r3_c6_5 = t_r3_c6_0 + p_2_5;
  assign t_r3_c6_6 = t_r3_c6_1 + p_2_7;
  assign t_r3_c6_7 = t_r3_c6_2 + t_r3_c6_3;
  assign t_r3_c6_8 = t_r3_c6_4 + p_4_5;
  assign t_r3_c6_9 = t_r3_c6_5 + t_r3_c6_6;
  assign t_r3_c6_10 = t_r3_c6_7 + t_r3_c6_8;
  assign t_r3_c6_11 = t_r3_c6_9 + t_r3_c6_10;
  assign t_r3_c6_12 = t_r3_c6_11 + p_4_7;
  assign out_3_6 = t_r3_c6_12 >> 4;

  assign t_r3_c7_0 = p_2_7 << 1;
  assign t_r3_c7_1 = p_3_6 << 1;
  assign t_r3_c7_2 = p_3_7 << 2;
  assign t_r3_c7_3 = p_3_8 << 1;
  assign t_r3_c7_4 = p_4_7 << 1;
  assign t_r3_c7_5 = t_r3_c7_0 + p_2_6;
  assign t_r3_c7_6 = t_r3_c7_1 + p_2_8;
  assign t_r3_c7_7 = t_r3_c7_2 + t_r3_c7_3;
  assign t_r3_c7_8 = t_r3_c7_4 + p_4_6;
  assign t_r3_c7_9 = t_r3_c7_5 + t_r3_c7_6;
  assign t_r3_c7_10 = t_r3_c7_7 + t_r3_c7_8;
  assign t_r3_c7_11 = t_r3_c7_9 + t_r3_c7_10;
  assign t_r3_c7_12 = t_r3_c7_11 + p_4_8;
  assign out_3_7 = t_r3_c7_12 >> 4;

  assign t_r3_c8_0 = p_2_8 << 1;
  assign t_r3_c8_1 = p_3_7 << 1;
  assign t_r3_c8_2 = p_3_8 << 2;
  assign t_r3_c8_3 = p_3_9 << 1;
  assign t_r3_c8_4 = p_4_8 << 1;
  assign t_r3_c8_5 = t_r3_c8_0 + p_2_7;
  assign t_r3_c8_6 = t_r3_c8_1 + p_2_9;
  assign t_r3_c8_7 = t_r3_c8_2 + t_r3_c8_3;
  assign t_r3_c8_8 = t_r3_c8_4 + p_4_7;
  assign t_r3_c8_9 = t_r3_c8_5 + t_r3_c8_6;
  assign t_r3_c8_10 = t_r3_c8_7 + t_r3_c8_8;
  assign t_r3_c8_11 = t_r3_c8_9 + t_r3_c8_10;
  assign t_r3_c8_12 = t_r3_c8_11 + p_4_9;
  assign out_3_8 = t_r3_c8_12 >> 4;

  assign t_r3_c9_0 = p_2_9 << 1;
  assign t_r3_c9_1 = p_3_8 << 1;
  assign t_r3_c9_2 = p_3_9 << 2;
  assign t_r3_c9_3 = p_3_10 << 1;
  assign t_r3_c9_4 = p_4_9 << 1;
  assign t_r3_c9_5 = t_r3_c9_0 + p_2_8;
  assign t_r3_c9_6 = t_r3_c9_1 + p_2_10;
  assign t_r3_c9_7 = t_r3_c9_2 + t_r3_c9_3;
  assign t_r3_c9_8 = t_r3_c9_4 + p_4_8;
  assign t_r3_c9_9 = t_r3_c9_5 + t_r3_c9_6;
  assign t_r3_c9_10 = t_r3_c9_7 + t_r3_c9_8;
  assign t_r3_c9_11 = t_r3_c9_9 + t_r3_c9_10;
  assign t_r3_c9_12 = t_r3_c9_11 + p_4_10;
  assign out_3_9 = t_r3_c9_12 >> 4;

  assign t_r3_c10_0 = p_2_10 << 1;
  assign t_r3_c10_1 = p_3_9 << 1;
  assign t_r3_c10_2 = p_3_10 << 2;
  assign t_r3_c10_3 = p_3_11 << 1;
  assign t_r3_c10_4 = p_4_10 << 1;
  assign t_r3_c10_5 = t_r3_c10_0 + p_2_9;
  assign t_r3_c10_6 = t_r3_c10_1 + p_2_11;
  assign t_r3_c10_7 = t_r3_c10_2 + t_r3_c10_3;
  assign t_r3_c10_8 = t_r3_c10_4 + p_4_9;
  assign t_r3_c10_9 = t_r3_c10_5 + t_r3_c10_6;
  assign t_r3_c10_10 = t_r3_c10_7 + t_r3_c10_8;
  assign t_r3_c10_11 = t_r3_c10_9 + t_r3_c10_10;
  assign t_r3_c10_12 = t_r3_c10_11 + p_4_11;
  assign out_3_10 = t_r3_c10_12 >> 4;

  assign t_r3_c11_0 = p_2_11 << 1;
  assign t_r3_c11_1 = p_3_10 << 1;
  assign t_r3_c11_2 = p_3_11 << 2;
  assign t_r3_c11_3 = p_3_12 << 1;
  assign t_r3_c11_4 = p_4_11 << 1;
  assign t_r3_c11_5 = t_r3_c11_0 + p_2_10;
  assign t_r3_c11_6 = t_r3_c11_1 + p_2_12;
  assign t_r3_c11_7 = t_r3_c11_2 + t_r3_c11_3;
  assign t_r3_c11_8 = t_r3_c11_4 + p_4_10;
  assign t_r3_c11_9 = t_r3_c11_5 + t_r3_c11_6;
  assign t_r3_c11_10 = t_r3_c11_7 + t_r3_c11_8;
  assign t_r3_c11_11 = t_r3_c11_9 + t_r3_c11_10;
  assign t_r3_c11_12 = t_r3_c11_11 + p_4_12;
  assign out_3_11 = t_r3_c11_12 >> 4;

  assign t_r3_c12_0 = p_2_12 << 1;
  assign t_r3_c12_1 = p_3_11 << 1;
  assign t_r3_c12_2 = p_3_12 << 2;
  assign t_r3_c12_3 = p_3_13 << 1;
  assign t_r3_c12_4 = p_4_12 << 1;
  assign t_r3_c12_5 = t_r3_c12_0 + p_2_11;
  assign t_r3_c12_6 = t_r3_c12_1 + p_2_13;
  assign t_r3_c12_7 = t_r3_c12_2 + t_r3_c12_3;
  assign t_r3_c12_8 = t_r3_c12_4 + p_4_11;
  assign t_r3_c12_9 = t_r3_c12_5 + t_r3_c12_6;
  assign t_r3_c12_10 = t_r3_c12_7 + t_r3_c12_8;
  assign t_r3_c12_11 = t_r3_c12_9 + t_r3_c12_10;
  assign t_r3_c12_12 = t_r3_c12_11 + p_4_13;
  assign out_3_12 = t_r3_c12_12 >> 4;

  assign t_r3_c13_0 = p_2_13 << 1;
  assign t_r3_c13_1 = p_3_12 << 1;
  assign t_r3_c13_2 = p_3_13 << 2;
  assign t_r3_c13_3 = p_3_14 << 1;
  assign t_r3_c13_4 = p_4_13 << 1;
  assign t_r3_c13_5 = t_r3_c13_0 + p_2_12;
  assign t_r3_c13_6 = t_r3_c13_1 + p_2_14;
  assign t_r3_c13_7 = t_r3_c13_2 + t_r3_c13_3;
  assign t_r3_c13_8 = t_r3_c13_4 + p_4_12;
  assign t_r3_c13_9 = t_r3_c13_5 + t_r3_c13_6;
  assign t_r3_c13_10 = t_r3_c13_7 + t_r3_c13_8;
  assign t_r3_c13_11 = t_r3_c13_9 + t_r3_c13_10;
  assign t_r3_c13_12 = t_r3_c13_11 + p_4_14;
  assign out_3_13 = t_r3_c13_12 >> 4;

  assign t_r3_c14_0 = p_2_14 << 1;
  assign t_r3_c14_1 = p_3_13 << 1;
  assign t_r3_c14_2 = p_3_14 << 2;
  assign t_r3_c14_3 = p_3_15 << 1;
  assign t_r3_c14_4 = p_4_14 << 1;
  assign t_r3_c14_5 = t_r3_c14_0 + p_2_13;
  assign t_r3_c14_6 = t_r3_c14_1 + p_2_15;
  assign t_r3_c14_7 = t_r3_c14_2 + t_r3_c14_3;
  assign t_r3_c14_8 = t_r3_c14_4 + p_4_13;
  assign t_r3_c14_9 = t_r3_c14_5 + t_r3_c14_6;
  assign t_r3_c14_10 = t_r3_c14_7 + t_r3_c14_8;
  assign t_r3_c14_11 = t_r3_c14_9 + t_r3_c14_10;
  assign t_r3_c14_12 = t_r3_c14_11 + p_4_15;
  assign out_3_14 = t_r3_c14_12 >> 4;

  assign t_r3_c15_0 = p_2_15 << 1;
  assign t_r3_c15_1 = p_3_14 << 1;
  assign t_r3_c15_2 = p_3_15 << 2;
  assign t_r3_c15_3 = p_3_16 << 1;
  assign t_r3_c15_4 = p_4_15 << 1;
  assign t_r3_c15_5 = t_r3_c15_0 + p_2_14;
  assign t_r3_c15_6 = t_r3_c15_1 + p_2_16;
  assign t_r3_c15_7 = t_r3_c15_2 + t_r3_c15_3;
  assign t_r3_c15_8 = t_r3_c15_4 + p_4_14;
  assign t_r3_c15_9 = t_r3_c15_5 + t_r3_c15_6;
  assign t_r3_c15_10 = t_r3_c15_7 + t_r3_c15_8;
  assign t_r3_c15_11 = t_r3_c15_9 + t_r3_c15_10;
  assign t_r3_c15_12 = t_r3_c15_11 + p_4_16;
  assign out_3_15 = t_r3_c15_12 >> 4;

  assign t_r3_c16_0 = p_2_16 << 1;
  assign t_r3_c16_1 = p_3_15 << 1;
  assign t_r3_c16_2 = p_3_16 << 2;
  assign t_r3_c16_3 = p_3_17 << 1;
  assign t_r3_c16_4 = p_4_16 << 1;
  assign t_r3_c16_5 = t_r3_c16_0 + p_2_15;
  assign t_r3_c16_6 = t_r3_c16_1 + p_2_17;
  assign t_r3_c16_7 = t_r3_c16_2 + t_r3_c16_3;
  assign t_r3_c16_8 = t_r3_c16_4 + p_4_15;
  assign t_r3_c16_9 = t_r3_c16_5 + t_r3_c16_6;
  assign t_r3_c16_10 = t_r3_c16_7 + t_r3_c16_8;
  assign t_r3_c16_11 = t_r3_c16_9 + t_r3_c16_10;
  assign t_r3_c16_12 = t_r3_c16_11 + p_4_17;
  assign out_3_16 = t_r3_c16_12 >> 4;

  assign t_r3_c17_0 = p_2_17 << 1;
  assign t_r3_c17_1 = p_3_16 << 1;
  assign t_r3_c17_2 = p_3_17 << 2;
  assign t_r3_c17_3 = p_3_18 << 1;
  assign t_r3_c17_4 = p_4_17 << 1;
  assign t_r3_c17_5 = t_r3_c17_0 + p_2_16;
  assign t_r3_c17_6 = t_r3_c17_1 + p_2_18;
  assign t_r3_c17_7 = t_r3_c17_2 + t_r3_c17_3;
  assign t_r3_c17_8 = t_r3_c17_4 + p_4_16;
  assign t_r3_c17_9 = t_r3_c17_5 + t_r3_c17_6;
  assign t_r3_c17_10 = t_r3_c17_7 + t_r3_c17_8;
  assign t_r3_c17_11 = t_r3_c17_9 + t_r3_c17_10;
  assign t_r3_c17_12 = t_r3_c17_11 + p_4_18;
  assign out_3_17 = t_r3_c17_12 >> 4;

  assign t_r3_c18_0 = p_2_18 << 1;
  assign t_r3_c18_1 = p_3_17 << 1;
  assign t_r3_c18_2 = p_3_18 << 2;
  assign t_r3_c18_3 = p_3_19 << 1;
  assign t_r3_c18_4 = p_4_18 << 1;
  assign t_r3_c18_5 = t_r3_c18_0 + p_2_17;
  assign t_r3_c18_6 = t_r3_c18_1 + p_2_19;
  assign t_r3_c18_7 = t_r3_c18_2 + t_r3_c18_3;
  assign t_r3_c18_8 = t_r3_c18_4 + p_4_17;
  assign t_r3_c18_9 = t_r3_c18_5 + t_r3_c18_6;
  assign t_r3_c18_10 = t_r3_c18_7 + t_r3_c18_8;
  assign t_r3_c18_11 = t_r3_c18_9 + t_r3_c18_10;
  assign t_r3_c18_12 = t_r3_c18_11 + p_4_19;
  assign out_3_18 = t_r3_c18_12 >> 4;

  assign t_r3_c19_0 = p_2_19 << 1;
  assign t_r3_c19_1 = p_3_18 << 1;
  assign t_r3_c19_2 = p_3_19 << 2;
  assign t_r3_c19_3 = p_3_20 << 1;
  assign t_r3_c19_4 = p_4_19 << 1;
  assign t_r3_c19_5 = t_r3_c19_0 + p_2_18;
  assign t_r3_c19_6 = t_r3_c19_1 + p_2_20;
  assign t_r3_c19_7 = t_r3_c19_2 + t_r3_c19_3;
  assign t_r3_c19_8 = t_r3_c19_4 + p_4_18;
  assign t_r3_c19_9 = t_r3_c19_5 + t_r3_c19_6;
  assign t_r3_c19_10 = t_r3_c19_7 + t_r3_c19_8;
  assign t_r3_c19_11 = t_r3_c19_9 + t_r3_c19_10;
  assign t_r3_c19_12 = t_r3_c19_11 + p_4_20;
  assign out_3_19 = t_r3_c19_12 >> 4;

  assign t_r3_c20_0 = p_2_20 << 1;
  assign t_r3_c20_1 = p_3_19 << 1;
  assign t_r3_c20_2 = p_3_20 << 2;
  assign t_r3_c20_3 = p_3_21 << 1;
  assign t_r3_c20_4 = p_4_20 << 1;
  assign t_r3_c20_5 = t_r3_c20_0 + p_2_19;
  assign t_r3_c20_6 = t_r3_c20_1 + p_2_21;
  assign t_r3_c20_7 = t_r3_c20_2 + t_r3_c20_3;
  assign t_r3_c20_8 = t_r3_c20_4 + p_4_19;
  assign t_r3_c20_9 = t_r3_c20_5 + t_r3_c20_6;
  assign t_r3_c20_10 = t_r3_c20_7 + t_r3_c20_8;
  assign t_r3_c20_11 = t_r3_c20_9 + t_r3_c20_10;
  assign t_r3_c20_12 = t_r3_c20_11 + p_4_21;
  assign out_3_20 = t_r3_c20_12 >> 4;

  assign t_r3_c21_0 = p_2_21 << 1;
  assign t_r3_c21_1 = p_3_20 << 1;
  assign t_r3_c21_2 = p_3_21 << 2;
  assign t_r3_c21_3 = p_3_22 << 1;
  assign t_r3_c21_4 = p_4_21 << 1;
  assign t_r3_c21_5 = t_r3_c21_0 + p_2_20;
  assign t_r3_c21_6 = t_r3_c21_1 + p_2_22;
  assign t_r3_c21_7 = t_r3_c21_2 + t_r3_c21_3;
  assign t_r3_c21_8 = t_r3_c21_4 + p_4_20;
  assign t_r3_c21_9 = t_r3_c21_5 + t_r3_c21_6;
  assign t_r3_c21_10 = t_r3_c21_7 + t_r3_c21_8;
  assign t_r3_c21_11 = t_r3_c21_9 + t_r3_c21_10;
  assign t_r3_c21_12 = t_r3_c21_11 + p_4_22;
  assign out_3_21 = t_r3_c21_12 >> 4;

  assign t_r3_c22_0 = p_2_22 << 1;
  assign t_r3_c22_1 = p_3_21 << 1;
  assign t_r3_c22_2 = p_3_22 << 2;
  assign t_r3_c22_3 = p_3_23 << 1;
  assign t_r3_c22_4 = p_4_22 << 1;
  assign t_r3_c22_5 = t_r3_c22_0 + p_2_21;
  assign t_r3_c22_6 = t_r3_c22_1 + p_2_23;
  assign t_r3_c22_7 = t_r3_c22_2 + t_r3_c22_3;
  assign t_r3_c22_8 = t_r3_c22_4 + p_4_21;
  assign t_r3_c22_9 = t_r3_c22_5 + t_r3_c22_6;
  assign t_r3_c22_10 = t_r3_c22_7 + t_r3_c22_8;
  assign t_r3_c22_11 = t_r3_c22_9 + t_r3_c22_10;
  assign t_r3_c22_12 = t_r3_c22_11 + p_4_23;
  assign out_3_22 = t_r3_c22_12 >> 4;

  assign t_r3_c23_0 = p_2_23 << 1;
  assign t_r3_c23_1 = p_3_22 << 1;
  assign t_r3_c23_2 = p_3_23 << 2;
  assign t_r3_c23_3 = p_3_24 << 1;
  assign t_r3_c23_4 = p_4_23 << 1;
  assign t_r3_c23_5 = t_r3_c23_0 + p_2_22;
  assign t_r3_c23_6 = t_r3_c23_1 + p_2_24;
  assign t_r3_c23_7 = t_r3_c23_2 + t_r3_c23_3;
  assign t_r3_c23_8 = t_r3_c23_4 + p_4_22;
  assign t_r3_c23_9 = t_r3_c23_5 + t_r3_c23_6;
  assign t_r3_c23_10 = t_r3_c23_7 + t_r3_c23_8;
  assign t_r3_c23_11 = t_r3_c23_9 + t_r3_c23_10;
  assign t_r3_c23_12 = t_r3_c23_11 + p_4_24;
  assign out_3_23 = t_r3_c23_12 >> 4;

  assign t_r3_c24_0 = p_2_24 << 1;
  assign t_r3_c24_1 = p_3_23 << 1;
  assign t_r3_c24_2 = p_3_24 << 2;
  assign t_r3_c24_3 = p_3_25 << 1;
  assign t_r3_c24_4 = p_4_24 << 1;
  assign t_r3_c24_5 = t_r3_c24_0 + p_2_23;
  assign t_r3_c24_6 = t_r3_c24_1 + p_2_25;
  assign t_r3_c24_7 = t_r3_c24_2 + t_r3_c24_3;
  assign t_r3_c24_8 = t_r3_c24_4 + p_4_23;
  assign t_r3_c24_9 = t_r3_c24_5 + t_r3_c24_6;
  assign t_r3_c24_10 = t_r3_c24_7 + t_r3_c24_8;
  assign t_r3_c24_11 = t_r3_c24_9 + t_r3_c24_10;
  assign t_r3_c24_12 = t_r3_c24_11 + p_4_25;
  assign out_3_24 = t_r3_c24_12 >> 4;

  assign t_r3_c25_0 = p_2_25 << 1;
  assign t_r3_c25_1 = p_3_24 << 1;
  assign t_r3_c25_2 = p_3_25 << 2;
  assign t_r3_c25_3 = p_3_26 << 1;
  assign t_r3_c25_4 = p_4_25 << 1;
  assign t_r3_c25_5 = t_r3_c25_0 + p_2_24;
  assign t_r3_c25_6 = t_r3_c25_1 + p_2_26;
  assign t_r3_c25_7 = t_r3_c25_2 + t_r3_c25_3;
  assign t_r3_c25_8 = t_r3_c25_4 + p_4_24;
  assign t_r3_c25_9 = t_r3_c25_5 + t_r3_c25_6;
  assign t_r3_c25_10 = t_r3_c25_7 + t_r3_c25_8;
  assign t_r3_c25_11 = t_r3_c25_9 + t_r3_c25_10;
  assign t_r3_c25_12 = t_r3_c25_11 + p_4_26;
  assign out_3_25 = t_r3_c25_12 >> 4;

  assign t_r3_c26_0 = p_2_26 << 1;
  assign t_r3_c26_1 = p_3_25 << 1;
  assign t_r3_c26_2 = p_3_26 << 2;
  assign t_r3_c26_3 = p_3_27 << 1;
  assign t_r3_c26_4 = p_4_26 << 1;
  assign t_r3_c26_5 = t_r3_c26_0 + p_2_25;
  assign t_r3_c26_6 = t_r3_c26_1 + p_2_27;
  assign t_r3_c26_7 = t_r3_c26_2 + t_r3_c26_3;
  assign t_r3_c26_8 = t_r3_c26_4 + p_4_25;
  assign t_r3_c26_9 = t_r3_c26_5 + t_r3_c26_6;
  assign t_r3_c26_10 = t_r3_c26_7 + t_r3_c26_8;
  assign t_r3_c26_11 = t_r3_c26_9 + t_r3_c26_10;
  assign t_r3_c26_12 = t_r3_c26_11 + p_4_27;
  assign out_3_26 = t_r3_c26_12 >> 4;

  assign t_r3_c27_0 = p_2_27 << 1;
  assign t_r3_c27_1 = p_3_26 << 1;
  assign t_r3_c27_2 = p_3_27 << 2;
  assign t_r3_c27_3 = p_3_28 << 1;
  assign t_r3_c27_4 = p_4_27 << 1;
  assign t_r3_c27_5 = t_r3_c27_0 + p_2_26;
  assign t_r3_c27_6 = t_r3_c27_1 + p_2_28;
  assign t_r3_c27_7 = t_r3_c27_2 + t_r3_c27_3;
  assign t_r3_c27_8 = t_r3_c27_4 + p_4_26;
  assign t_r3_c27_9 = t_r3_c27_5 + t_r3_c27_6;
  assign t_r3_c27_10 = t_r3_c27_7 + t_r3_c27_8;
  assign t_r3_c27_11 = t_r3_c27_9 + t_r3_c27_10;
  assign t_r3_c27_12 = t_r3_c27_11 + p_4_28;
  assign out_3_27 = t_r3_c27_12 >> 4;

  assign t_r3_c28_0 = p_2_28 << 1;
  assign t_r3_c28_1 = p_3_27 << 1;
  assign t_r3_c28_2 = p_3_28 << 2;
  assign t_r3_c28_3 = p_3_29 << 1;
  assign t_r3_c28_4 = p_4_28 << 1;
  assign t_r3_c28_5 = t_r3_c28_0 + p_2_27;
  assign t_r3_c28_6 = t_r3_c28_1 + p_2_29;
  assign t_r3_c28_7 = t_r3_c28_2 + t_r3_c28_3;
  assign t_r3_c28_8 = t_r3_c28_4 + p_4_27;
  assign t_r3_c28_9 = t_r3_c28_5 + t_r3_c28_6;
  assign t_r3_c28_10 = t_r3_c28_7 + t_r3_c28_8;
  assign t_r3_c28_11 = t_r3_c28_9 + t_r3_c28_10;
  assign t_r3_c28_12 = t_r3_c28_11 + p_4_29;
  assign out_3_28 = t_r3_c28_12 >> 4;

  assign t_r3_c29_0 = p_2_29 << 1;
  assign t_r3_c29_1 = p_3_28 << 1;
  assign t_r3_c29_2 = p_3_29 << 2;
  assign t_r3_c29_3 = p_3_30 << 1;
  assign t_r3_c29_4 = p_4_29 << 1;
  assign t_r3_c29_5 = t_r3_c29_0 + p_2_28;
  assign t_r3_c29_6 = t_r3_c29_1 + p_2_30;
  assign t_r3_c29_7 = t_r3_c29_2 + t_r3_c29_3;
  assign t_r3_c29_8 = t_r3_c29_4 + p_4_28;
  assign t_r3_c29_9 = t_r3_c29_5 + t_r3_c29_6;
  assign t_r3_c29_10 = t_r3_c29_7 + t_r3_c29_8;
  assign t_r3_c29_11 = t_r3_c29_9 + t_r3_c29_10;
  assign t_r3_c29_12 = t_r3_c29_11 + p_4_30;
  assign out_3_29 = t_r3_c29_12 >> 4;

  assign t_r3_c30_0 = p_2_30 << 1;
  assign t_r3_c30_1 = p_3_29 << 1;
  assign t_r3_c30_2 = p_3_30 << 2;
  assign t_r3_c30_3 = p_3_31 << 1;
  assign t_r3_c30_4 = p_4_30 << 1;
  assign t_r3_c30_5 = t_r3_c30_0 + p_2_29;
  assign t_r3_c30_6 = t_r3_c30_1 + p_2_31;
  assign t_r3_c30_7 = t_r3_c30_2 + t_r3_c30_3;
  assign t_r3_c30_8 = t_r3_c30_4 + p_4_29;
  assign t_r3_c30_9 = t_r3_c30_5 + t_r3_c30_6;
  assign t_r3_c30_10 = t_r3_c30_7 + t_r3_c30_8;
  assign t_r3_c30_11 = t_r3_c30_9 + t_r3_c30_10;
  assign t_r3_c30_12 = t_r3_c30_11 + p_4_31;
  assign out_3_30 = t_r3_c30_12 >> 4;

  assign t_r3_c31_0 = p_2_31 << 1;
  assign t_r3_c31_1 = p_3_30 << 1;
  assign t_r3_c31_2 = p_3_31 << 2;
  assign t_r3_c31_3 = p_3_32 << 1;
  assign t_r3_c31_4 = p_4_31 << 1;
  assign t_r3_c31_5 = t_r3_c31_0 + p_2_30;
  assign t_r3_c31_6 = t_r3_c31_1 + p_2_32;
  assign t_r3_c31_7 = t_r3_c31_2 + t_r3_c31_3;
  assign t_r3_c31_8 = t_r3_c31_4 + p_4_30;
  assign t_r3_c31_9 = t_r3_c31_5 + t_r3_c31_6;
  assign t_r3_c31_10 = t_r3_c31_7 + t_r3_c31_8;
  assign t_r3_c31_11 = t_r3_c31_9 + t_r3_c31_10;
  assign t_r3_c31_12 = t_r3_c31_11 + p_4_32;
  assign out_3_31 = t_r3_c31_12 >> 4;

  assign t_r3_c32_0 = p_2_32 << 1;
  assign t_r3_c32_1 = p_3_31 << 1;
  assign t_r3_c32_2 = p_3_32 << 2;
  assign t_r3_c32_3 = p_3_33 << 1;
  assign t_r3_c32_4 = p_4_32 << 1;
  assign t_r3_c32_5 = t_r3_c32_0 + p_2_31;
  assign t_r3_c32_6 = t_r3_c32_1 + p_2_33;
  assign t_r3_c32_7 = t_r3_c32_2 + t_r3_c32_3;
  assign t_r3_c32_8 = t_r3_c32_4 + p_4_31;
  assign t_r3_c32_9 = t_r3_c32_5 + t_r3_c32_6;
  assign t_r3_c32_10 = t_r3_c32_7 + t_r3_c32_8;
  assign t_r3_c32_11 = t_r3_c32_9 + t_r3_c32_10;
  assign t_r3_c32_12 = t_r3_c32_11 + p_4_33;
  assign out_3_32 = t_r3_c32_12 >> 4;

  assign t_r3_c33_0 = p_2_33 << 1;
  assign t_r3_c33_1 = p_3_32 << 1;
  assign t_r3_c33_2 = p_3_33 << 2;
  assign t_r3_c33_3 = p_3_34 << 1;
  assign t_r3_c33_4 = p_4_33 << 1;
  assign t_r3_c33_5 = t_r3_c33_0 + p_2_32;
  assign t_r3_c33_6 = t_r3_c33_1 + p_2_34;
  assign t_r3_c33_7 = t_r3_c33_2 + t_r3_c33_3;
  assign t_r3_c33_8 = t_r3_c33_4 + p_4_32;
  assign t_r3_c33_9 = t_r3_c33_5 + t_r3_c33_6;
  assign t_r3_c33_10 = t_r3_c33_7 + t_r3_c33_8;
  assign t_r3_c33_11 = t_r3_c33_9 + t_r3_c33_10;
  assign t_r3_c33_12 = t_r3_c33_11 + p_4_34;
  assign out_3_33 = t_r3_c33_12 >> 4;

  assign t_r3_c34_0 = p_2_34 << 1;
  assign t_r3_c34_1 = p_3_33 << 1;
  assign t_r3_c34_2 = p_3_34 << 2;
  assign t_r3_c34_3 = p_3_35 << 1;
  assign t_r3_c34_4 = p_4_34 << 1;
  assign t_r3_c34_5 = t_r3_c34_0 + p_2_33;
  assign t_r3_c34_6 = t_r3_c34_1 + p_2_35;
  assign t_r3_c34_7 = t_r3_c34_2 + t_r3_c34_3;
  assign t_r3_c34_8 = t_r3_c34_4 + p_4_33;
  assign t_r3_c34_9 = t_r3_c34_5 + t_r3_c34_6;
  assign t_r3_c34_10 = t_r3_c34_7 + t_r3_c34_8;
  assign t_r3_c34_11 = t_r3_c34_9 + t_r3_c34_10;
  assign t_r3_c34_12 = t_r3_c34_11 + p_4_35;
  assign out_3_34 = t_r3_c34_12 >> 4;

  assign t_r3_c35_0 = p_2_35 << 1;
  assign t_r3_c35_1 = p_3_34 << 1;
  assign t_r3_c35_2 = p_3_35 << 2;
  assign t_r3_c35_3 = p_3_36 << 1;
  assign t_r3_c35_4 = p_4_35 << 1;
  assign t_r3_c35_5 = t_r3_c35_0 + p_2_34;
  assign t_r3_c35_6 = t_r3_c35_1 + p_2_36;
  assign t_r3_c35_7 = t_r3_c35_2 + t_r3_c35_3;
  assign t_r3_c35_8 = t_r3_c35_4 + p_4_34;
  assign t_r3_c35_9 = t_r3_c35_5 + t_r3_c35_6;
  assign t_r3_c35_10 = t_r3_c35_7 + t_r3_c35_8;
  assign t_r3_c35_11 = t_r3_c35_9 + t_r3_c35_10;
  assign t_r3_c35_12 = t_r3_c35_11 + p_4_36;
  assign out_3_35 = t_r3_c35_12 >> 4;

  assign t_r3_c36_0 = p_2_36 << 1;
  assign t_r3_c36_1 = p_3_35 << 1;
  assign t_r3_c36_2 = p_3_36 << 2;
  assign t_r3_c36_3 = p_3_37 << 1;
  assign t_r3_c36_4 = p_4_36 << 1;
  assign t_r3_c36_5 = t_r3_c36_0 + p_2_35;
  assign t_r3_c36_6 = t_r3_c36_1 + p_2_37;
  assign t_r3_c36_7 = t_r3_c36_2 + t_r3_c36_3;
  assign t_r3_c36_8 = t_r3_c36_4 + p_4_35;
  assign t_r3_c36_9 = t_r3_c36_5 + t_r3_c36_6;
  assign t_r3_c36_10 = t_r3_c36_7 + t_r3_c36_8;
  assign t_r3_c36_11 = t_r3_c36_9 + t_r3_c36_10;
  assign t_r3_c36_12 = t_r3_c36_11 + p_4_37;
  assign out_3_36 = t_r3_c36_12 >> 4;

  assign t_r3_c37_0 = p_2_37 << 1;
  assign t_r3_c37_1 = p_3_36 << 1;
  assign t_r3_c37_2 = p_3_37 << 2;
  assign t_r3_c37_3 = p_3_38 << 1;
  assign t_r3_c37_4 = p_4_37 << 1;
  assign t_r3_c37_5 = t_r3_c37_0 + p_2_36;
  assign t_r3_c37_6 = t_r3_c37_1 + p_2_38;
  assign t_r3_c37_7 = t_r3_c37_2 + t_r3_c37_3;
  assign t_r3_c37_8 = t_r3_c37_4 + p_4_36;
  assign t_r3_c37_9 = t_r3_c37_5 + t_r3_c37_6;
  assign t_r3_c37_10 = t_r3_c37_7 + t_r3_c37_8;
  assign t_r3_c37_11 = t_r3_c37_9 + t_r3_c37_10;
  assign t_r3_c37_12 = t_r3_c37_11 + p_4_38;
  assign out_3_37 = t_r3_c37_12 >> 4;

  assign t_r3_c38_0 = p_2_38 << 1;
  assign t_r3_c38_1 = p_3_37 << 1;
  assign t_r3_c38_2 = p_3_38 << 2;
  assign t_r3_c38_3 = p_3_39 << 1;
  assign t_r3_c38_4 = p_4_38 << 1;
  assign t_r3_c38_5 = t_r3_c38_0 + p_2_37;
  assign t_r3_c38_6 = t_r3_c38_1 + p_2_39;
  assign t_r3_c38_7 = t_r3_c38_2 + t_r3_c38_3;
  assign t_r3_c38_8 = t_r3_c38_4 + p_4_37;
  assign t_r3_c38_9 = t_r3_c38_5 + t_r3_c38_6;
  assign t_r3_c38_10 = t_r3_c38_7 + t_r3_c38_8;
  assign t_r3_c38_11 = t_r3_c38_9 + t_r3_c38_10;
  assign t_r3_c38_12 = t_r3_c38_11 + p_4_39;
  assign out_3_38 = t_r3_c38_12 >> 4;

  assign t_r3_c39_0 = p_2_39 << 1;
  assign t_r3_c39_1 = p_3_38 << 1;
  assign t_r3_c39_2 = p_3_39 << 2;
  assign t_r3_c39_3 = p_3_40 << 1;
  assign t_r3_c39_4 = p_4_39 << 1;
  assign t_r3_c39_5 = t_r3_c39_0 + p_2_38;
  assign t_r3_c39_6 = t_r3_c39_1 + p_2_40;
  assign t_r3_c39_7 = t_r3_c39_2 + t_r3_c39_3;
  assign t_r3_c39_8 = t_r3_c39_4 + p_4_38;
  assign t_r3_c39_9 = t_r3_c39_5 + t_r3_c39_6;
  assign t_r3_c39_10 = t_r3_c39_7 + t_r3_c39_8;
  assign t_r3_c39_11 = t_r3_c39_9 + t_r3_c39_10;
  assign t_r3_c39_12 = t_r3_c39_11 + p_4_40;
  assign out_3_39 = t_r3_c39_12 >> 4;

  assign t_r3_c40_0 = p_2_40 << 1;
  assign t_r3_c40_1 = p_3_39 << 1;
  assign t_r3_c40_2 = p_3_40 << 2;
  assign t_r3_c40_3 = p_3_41 << 1;
  assign t_r3_c40_4 = p_4_40 << 1;
  assign t_r3_c40_5 = t_r3_c40_0 + p_2_39;
  assign t_r3_c40_6 = t_r3_c40_1 + p_2_41;
  assign t_r3_c40_7 = t_r3_c40_2 + t_r3_c40_3;
  assign t_r3_c40_8 = t_r3_c40_4 + p_4_39;
  assign t_r3_c40_9 = t_r3_c40_5 + t_r3_c40_6;
  assign t_r3_c40_10 = t_r3_c40_7 + t_r3_c40_8;
  assign t_r3_c40_11 = t_r3_c40_9 + t_r3_c40_10;
  assign t_r3_c40_12 = t_r3_c40_11 + p_4_41;
  assign out_3_40 = t_r3_c40_12 >> 4;

  assign t_r3_c41_0 = p_2_41 << 1;
  assign t_r3_c41_1 = p_3_40 << 1;
  assign t_r3_c41_2 = p_3_41 << 2;
  assign t_r3_c41_3 = p_3_42 << 1;
  assign t_r3_c41_4 = p_4_41 << 1;
  assign t_r3_c41_5 = t_r3_c41_0 + p_2_40;
  assign t_r3_c41_6 = t_r3_c41_1 + p_2_42;
  assign t_r3_c41_7 = t_r3_c41_2 + t_r3_c41_3;
  assign t_r3_c41_8 = t_r3_c41_4 + p_4_40;
  assign t_r3_c41_9 = t_r3_c41_5 + t_r3_c41_6;
  assign t_r3_c41_10 = t_r3_c41_7 + t_r3_c41_8;
  assign t_r3_c41_11 = t_r3_c41_9 + t_r3_c41_10;
  assign t_r3_c41_12 = t_r3_c41_11 + p_4_42;
  assign out_3_41 = t_r3_c41_12 >> 4;

  assign t_r3_c42_0 = p_2_42 << 1;
  assign t_r3_c42_1 = p_3_41 << 1;
  assign t_r3_c42_2 = p_3_42 << 2;
  assign t_r3_c42_3 = p_3_43 << 1;
  assign t_r3_c42_4 = p_4_42 << 1;
  assign t_r3_c42_5 = t_r3_c42_0 + p_2_41;
  assign t_r3_c42_6 = t_r3_c42_1 + p_2_43;
  assign t_r3_c42_7 = t_r3_c42_2 + t_r3_c42_3;
  assign t_r3_c42_8 = t_r3_c42_4 + p_4_41;
  assign t_r3_c42_9 = t_r3_c42_5 + t_r3_c42_6;
  assign t_r3_c42_10 = t_r3_c42_7 + t_r3_c42_8;
  assign t_r3_c42_11 = t_r3_c42_9 + t_r3_c42_10;
  assign t_r3_c42_12 = t_r3_c42_11 + p_4_43;
  assign out_3_42 = t_r3_c42_12 >> 4;

  assign t_r3_c43_0 = p_2_43 << 1;
  assign t_r3_c43_1 = p_3_42 << 1;
  assign t_r3_c43_2 = p_3_43 << 2;
  assign t_r3_c43_3 = p_3_44 << 1;
  assign t_r3_c43_4 = p_4_43 << 1;
  assign t_r3_c43_5 = t_r3_c43_0 + p_2_42;
  assign t_r3_c43_6 = t_r3_c43_1 + p_2_44;
  assign t_r3_c43_7 = t_r3_c43_2 + t_r3_c43_3;
  assign t_r3_c43_8 = t_r3_c43_4 + p_4_42;
  assign t_r3_c43_9 = t_r3_c43_5 + t_r3_c43_6;
  assign t_r3_c43_10 = t_r3_c43_7 + t_r3_c43_8;
  assign t_r3_c43_11 = t_r3_c43_9 + t_r3_c43_10;
  assign t_r3_c43_12 = t_r3_c43_11 + p_4_44;
  assign out_3_43 = t_r3_c43_12 >> 4;

  assign t_r3_c44_0 = p_2_44 << 1;
  assign t_r3_c44_1 = p_3_43 << 1;
  assign t_r3_c44_2 = p_3_44 << 2;
  assign t_r3_c44_3 = p_3_45 << 1;
  assign t_r3_c44_4 = p_4_44 << 1;
  assign t_r3_c44_5 = t_r3_c44_0 + p_2_43;
  assign t_r3_c44_6 = t_r3_c44_1 + p_2_45;
  assign t_r3_c44_7 = t_r3_c44_2 + t_r3_c44_3;
  assign t_r3_c44_8 = t_r3_c44_4 + p_4_43;
  assign t_r3_c44_9 = t_r3_c44_5 + t_r3_c44_6;
  assign t_r3_c44_10 = t_r3_c44_7 + t_r3_c44_8;
  assign t_r3_c44_11 = t_r3_c44_9 + t_r3_c44_10;
  assign t_r3_c44_12 = t_r3_c44_11 + p_4_45;
  assign out_3_44 = t_r3_c44_12 >> 4;

  assign t_r3_c45_0 = p_2_45 << 1;
  assign t_r3_c45_1 = p_3_44 << 1;
  assign t_r3_c45_2 = p_3_45 << 2;
  assign t_r3_c45_3 = p_3_46 << 1;
  assign t_r3_c45_4 = p_4_45 << 1;
  assign t_r3_c45_5 = t_r3_c45_0 + p_2_44;
  assign t_r3_c45_6 = t_r3_c45_1 + p_2_46;
  assign t_r3_c45_7 = t_r3_c45_2 + t_r3_c45_3;
  assign t_r3_c45_8 = t_r3_c45_4 + p_4_44;
  assign t_r3_c45_9 = t_r3_c45_5 + t_r3_c45_6;
  assign t_r3_c45_10 = t_r3_c45_7 + t_r3_c45_8;
  assign t_r3_c45_11 = t_r3_c45_9 + t_r3_c45_10;
  assign t_r3_c45_12 = t_r3_c45_11 + p_4_46;
  assign out_3_45 = t_r3_c45_12 >> 4;

  assign t_r3_c46_0 = p_2_46 << 1;
  assign t_r3_c46_1 = p_3_45 << 1;
  assign t_r3_c46_2 = p_3_46 << 2;
  assign t_r3_c46_3 = p_3_47 << 1;
  assign t_r3_c46_4 = p_4_46 << 1;
  assign t_r3_c46_5 = t_r3_c46_0 + p_2_45;
  assign t_r3_c46_6 = t_r3_c46_1 + p_2_47;
  assign t_r3_c46_7 = t_r3_c46_2 + t_r3_c46_3;
  assign t_r3_c46_8 = t_r3_c46_4 + p_4_45;
  assign t_r3_c46_9 = t_r3_c46_5 + t_r3_c46_6;
  assign t_r3_c46_10 = t_r3_c46_7 + t_r3_c46_8;
  assign t_r3_c46_11 = t_r3_c46_9 + t_r3_c46_10;
  assign t_r3_c46_12 = t_r3_c46_11 + p_4_47;
  assign out_3_46 = t_r3_c46_12 >> 4;

  assign t_r3_c47_0 = p_2_47 << 1;
  assign t_r3_c47_1 = p_3_46 << 1;
  assign t_r3_c47_2 = p_3_47 << 2;
  assign t_r3_c47_3 = p_3_48 << 1;
  assign t_r3_c47_4 = p_4_47 << 1;
  assign t_r3_c47_5 = t_r3_c47_0 + p_2_46;
  assign t_r3_c47_6 = t_r3_c47_1 + p_2_48;
  assign t_r3_c47_7 = t_r3_c47_2 + t_r3_c47_3;
  assign t_r3_c47_8 = t_r3_c47_4 + p_4_46;
  assign t_r3_c47_9 = t_r3_c47_5 + t_r3_c47_6;
  assign t_r3_c47_10 = t_r3_c47_7 + t_r3_c47_8;
  assign t_r3_c47_11 = t_r3_c47_9 + t_r3_c47_10;
  assign t_r3_c47_12 = t_r3_c47_11 + p_4_48;
  assign out_3_47 = t_r3_c47_12 >> 4;

  assign t_r3_c48_0 = p_2_48 << 1;
  assign t_r3_c48_1 = p_3_47 << 1;
  assign t_r3_c48_2 = p_3_48 << 2;
  assign t_r3_c48_3 = p_3_49 << 1;
  assign t_r3_c48_4 = p_4_48 << 1;
  assign t_r3_c48_5 = t_r3_c48_0 + p_2_47;
  assign t_r3_c48_6 = t_r3_c48_1 + p_2_49;
  assign t_r3_c48_7 = t_r3_c48_2 + t_r3_c48_3;
  assign t_r3_c48_8 = t_r3_c48_4 + p_4_47;
  assign t_r3_c48_9 = t_r3_c48_5 + t_r3_c48_6;
  assign t_r3_c48_10 = t_r3_c48_7 + t_r3_c48_8;
  assign t_r3_c48_11 = t_r3_c48_9 + t_r3_c48_10;
  assign t_r3_c48_12 = t_r3_c48_11 + p_4_49;
  assign out_3_48 = t_r3_c48_12 >> 4;

  assign t_r3_c49_0 = p_2_49 << 1;
  assign t_r3_c49_1 = p_3_48 << 1;
  assign t_r3_c49_2 = p_3_49 << 2;
  assign t_r3_c49_3 = p_3_50 << 1;
  assign t_r3_c49_4 = p_4_49 << 1;
  assign t_r3_c49_5 = t_r3_c49_0 + p_2_48;
  assign t_r3_c49_6 = t_r3_c49_1 + p_2_50;
  assign t_r3_c49_7 = t_r3_c49_2 + t_r3_c49_3;
  assign t_r3_c49_8 = t_r3_c49_4 + p_4_48;
  assign t_r3_c49_9 = t_r3_c49_5 + t_r3_c49_6;
  assign t_r3_c49_10 = t_r3_c49_7 + t_r3_c49_8;
  assign t_r3_c49_11 = t_r3_c49_9 + t_r3_c49_10;
  assign t_r3_c49_12 = t_r3_c49_11 + p_4_50;
  assign out_3_49 = t_r3_c49_12 >> 4;

  assign t_r3_c50_0 = p_2_50 << 1;
  assign t_r3_c50_1 = p_3_49 << 1;
  assign t_r3_c50_2 = p_3_50 << 2;
  assign t_r3_c50_3 = p_3_51 << 1;
  assign t_r3_c50_4 = p_4_50 << 1;
  assign t_r3_c50_5 = t_r3_c50_0 + p_2_49;
  assign t_r3_c50_6 = t_r3_c50_1 + p_2_51;
  assign t_r3_c50_7 = t_r3_c50_2 + t_r3_c50_3;
  assign t_r3_c50_8 = t_r3_c50_4 + p_4_49;
  assign t_r3_c50_9 = t_r3_c50_5 + t_r3_c50_6;
  assign t_r3_c50_10 = t_r3_c50_7 + t_r3_c50_8;
  assign t_r3_c50_11 = t_r3_c50_9 + t_r3_c50_10;
  assign t_r3_c50_12 = t_r3_c50_11 + p_4_51;
  assign out_3_50 = t_r3_c50_12 >> 4;

  assign t_r3_c51_0 = p_2_51 << 1;
  assign t_r3_c51_1 = p_3_50 << 1;
  assign t_r3_c51_2 = p_3_51 << 2;
  assign t_r3_c51_3 = p_3_52 << 1;
  assign t_r3_c51_4 = p_4_51 << 1;
  assign t_r3_c51_5 = t_r3_c51_0 + p_2_50;
  assign t_r3_c51_6 = t_r3_c51_1 + p_2_52;
  assign t_r3_c51_7 = t_r3_c51_2 + t_r3_c51_3;
  assign t_r3_c51_8 = t_r3_c51_4 + p_4_50;
  assign t_r3_c51_9 = t_r3_c51_5 + t_r3_c51_6;
  assign t_r3_c51_10 = t_r3_c51_7 + t_r3_c51_8;
  assign t_r3_c51_11 = t_r3_c51_9 + t_r3_c51_10;
  assign t_r3_c51_12 = t_r3_c51_11 + p_4_52;
  assign out_3_51 = t_r3_c51_12 >> 4;

  assign t_r3_c52_0 = p_2_52 << 1;
  assign t_r3_c52_1 = p_3_51 << 1;
  assign t_r3_c52_2 = p_3_52 << 2;
  assign t_r3_c52_3 = p_3_53 << 1;
  assign t_r3_c52_4 = p_4_52 << 1;
  assign t_r3_c52_5 = t_r3_c52_0 + p_2_51;
  assign t_r3_c52_6 = t_r3_c52_1 + p_2_53;
  assign t_r3_c52_7 = t_r3_c52_2 + t_r3_c52_3;
  assign t_r3_c52_8 = t_r3_c52_4 + p_4_51;
  assign t_r3_c52_9 = t_r3_c52_5 + t_r3_c52_6;
  assign t_r3_c52_10 = t_r3_c52_7 + t_r3_c52_8;
  assign t_r3_c52_11 = t_r3_c52_9 + t_r3_c52_10;
  assign t_r3_c52_12 = t_r3_c52_11 + p_4_53;
  assign out_3_52 = t_r3_c52_12 >> 4;

  assign t_r3_c53_0 = p_2_53 << 1;
  assign t_r3_c53_1 = p_3_52 << 1;
  assign t_r3_c53_2 = p_3_53 << 2;
  assign t_r3_c53_3 = p_3_54 << 1;
  assign t_r3_c53_4 = p_4_53 << 1;
  assign t_r3_c53_5 = t_r3_c53_0 + p_2_52;
  assign t_r3_c53_6 = t_r3_c53_1 + p_2_54;
  assign t_r3_c53_7 = t_r3_c53_2 + t_r3_c53_3;
  assign t_r3_c53_8 = t_r3_c53_4 + p_4_52;
  assign t_r3_c53_9 = t_r3_c53_5 + t_r3_c53_6;
  assign t_r3_c53_10 = t_r3_c53_7 + t_r3_c53_8;
  assign t_r3_c53_11 = t_r3_c53_9 + t_r3_c53_10;
  assign t_r3_c53_12 = t_r3_c53_11 + p_4_54;
  assign out_3_53 = t_r3_c53_12 >> 4;

  assign t_r3_c54_0 = p_2_54 << 1;
  assign t_r3_c54_1 = p_3_53 << 1;
  assign t_r3_c54_2 = p_3_54 << 2;
  assign t_r3_c54_3 = p_3_55 << 1;
  assign t_r3_c54_4 = p_4_54 << 1;
  assign t_r3_c54_5 = t_r3_c54_0 + p_2_53;
  assign t_r3_c54_6 = t_r3_c54_1 + p_2_55;
  assign t_r3_c54_7 = t_r3_c54_2 + t_r3_c54_3;
  assign t_r3_c54_8 = t_r3_c54_4 + p_4_53;
  assign t_r3_c54_9 = t_r3_c54_5 + t_r3_c54_6;
  assign t_r3_c54_10 = t_r3_c54_7 + t_r3_c54_8;
  assign t_r3_c54_11 = t_r3_c54_9 + t_r3_c54_10;
  assign t_r3_c54_12 = t_r3_c54_11 + p_4_55;
  assign out_3_54 = t_r3_c54_12 >> 4;

  assign t_r3_c55_0 = p_2_55 << 1;
  assign t_r3_c55_1 = p_3_54 << 1;
  assign t_r3_c55_2 = p_3_55 << 2;
  assign t_r3_c55_3 = p_3_56 << 1;
  assign t_r3_c55_4 = p_4_55 << 1;
  assign t_r3_c55_5 = t_r3_c55_0 + p_2_54;
  assign t_r3_c55_6 = t_r3_c55_1 + p_2_56;
  assign t_r3_c55_7 = t_r3_c55_2 + t_r3_c55_3;
  assign t_r3_c55_8 = t_r3_c55_4 + p_4_54;
  assign t_r3_c55_9 = t_r3_c55_5 + t_r3_c55_6;
  assign t_r3_c55_10 = t_r3_c55_7 + t_r3_c55_8;
  assign t_r3_c55_11 = t_r3_c55_9 + t_r3_c55_10;
  assign t_r3_c55_12 = t_r3_c55_11 + p_4_56;
  assign out_3_55 = t_r3_c55_12 >> 4;

  assign t_r3_c56_0 = p_2_56 << 1;
  assign t_r3_c56_1 = p_3_55 << 1;
  assign t_r3_c56_2 = p_3_56 << 2;
  assign t_r3_c56_3 = p_3_57 << 1;
  assign t_r3_c56_4 = p_4_56 << 1;
  assign t_r3_c56_5 = t_r3_c56_0 + p_2_55;
  assign t_r3_c56_6 = t_r3_c56_1 + p_2_57;
  assign t_r3_c56_7 = t_r3_c56_2 + t_r3_c56_3;
  assign t_r3_c56_8 = t_r3_c56_4 + p_4_55;
  assign t_r3_c56_9 = t_r3_c56_5 + t_r3_c56_6;
  assign t_r3_c56_10 = t_r3_c56_7 + t_r3_c56_8;
  assign t_r3_c56_11 = t_r3_c56_9 + t_r3_c56_10;
  assign t_r3_c56_12 = t_r3_c56_11 + p_4_57;
  assign out_3_56 = t_r3_c56_12 >> 4;

  assign t_r3_c57_0 = p_2_57 << 1;
  assign t_r3_c57_1 = p_3_56 << 1;
  assign t_r3_c57_2 = p_3_57 << 2;
  assign t_r3_c57_3 = p_3_58 << 1;
  assign t_r3_c57_4 = p_4_57 << 1;
  assign t_r3_c57_5 = t_r3_c57_0 + p_2_56;
  assign t_r3_c57_6 = t_r3_c57_1 + p_2_58;
  assign t_r3_c57_7 = t_r3_c57_2 + t_r3_c57_3;
  assign t_r3_c57_8 = t_r3_c57_4 + p_4_56;
  assign t_r3_c57_9 = t_r3_c57_5 + t_r3_c57_6;
  assign t_r3_c57_10 = t_r3_c57_7 + t_r3_c57_8;
  assign t_r3_c57_11 = t_r3_c57_9 + t_r3_c57_10;
  assign t_r3_c57_12 = t_r3_c57_11 + p_4_58;
  assign out_3_57 = t_r3_c57_12 >> 4;

  assign t_r3_c58_0 = p_2_58 << 1;
  assign t_r3_c58_1 = p_3_57 << 1;
  assign t_r3_c58_2 = p_3_58 << 2;
  assign t_r3_c58_3 = p_3_59 << 1;
  assign t_r3_c58_4 = p_4_58 << 1;
  assign t_r3_c58_5 = t_r3_c58_0 + p_2_57;
  assign t_r3_c58_6 = t_r3_c58_1 + p_2_59;
  assign t_r3_c58_7 = t_r3_c58_2 + t_r3_c58_3;
  assign t_r3_c58_8 = t_r3_c58_4 + p_4_57;
  assign t_r3_c58_9 = t_r3_c58_5 + t_r3_c58_6;
  assign t_r3_c58_10 = t_r3_c58_7 + t_r3_c58_8;
  assign t_r3_c58_11 = t_r3_c58_9 + t_r3_c58_10;
  assign t_r3_c58_12 = t_r3_c58_11 + p_4_59;
  assign out_3_58 = t_r3_c58_12 >> 4;

  assign t_r3_c59_0 = p_2_59 << 1;
  assign t_r3_c59_1 = p_3_58 << 1;
  assign t_r3_c59_2 = p_3_59 << 2;
  assign t_r3_c59_3 = p_3_60 << 1;
  assign t_r3_c59_4 = p_4_59 << 1;
  assign t_r3_c59_5 = t_r3_c59_0 + p_2_58;
  assign t_r3_c59_6 = t_r3_c59_1 + p_2_60;
  assign t_r3_c59_7 = t_r3_c59_2 + t_r3_c59_3;
  assign t_r3_c59_8 = t_r3_c59_4 + p_4_58;
  assign t_r3_c59_9 = t_r3_c59_5 + t_r3_c59_6;
  assign t_r3_c59_10 = t_r3_c59_7 + t_r3_c59_8;
  assign t_r3_c59_11 = t_r3_c59_9 + t_r3_c59_10;
  assign t_r3_c59_12 = t_r3_c59_11 + p_4_60;
  assign out_3_59 = t_r3_c59_12 >> 4;

  assign t_r3_c60_0 = p_2_60 << 1;
  assign t_r3_c60_1 = p_3_59 << 1;
  assign t_r3_c60_2 = p_3_60 << 2;
  assign t_r3_c60_3 = p_3_61 << 1;
  assign t_r3_c60_4 = p_4_60 << 1;
  assign t_r3_c60_5 = t_r3_c60_0 + p_2_59;
  assign t_r3_c60_6 = t_r3_c60_1 + p_2_61;
  assign t_r3_c60_7 = t_r3_c60_2 + t_r3_c60_3;
  assign t_r3_c60_8 = t_r3_c60_4 + p_4_59;
  assign t_r3_c60_9 = t_r3_c60_5 + t_r3_c60_6;
  assign t_r3_c60_10 = t_r3_c60_7 + t_r3_c60_8;
  assign t_r3_c60_11 = t_r3_c60_9 + t_r3_c60_10;
  assign t_r3_c60_12 = t_r3_c60_11 + p_4_61;
  assign out_3_60 = t_r3_c60_12 >> 4;

  assign t_r3_c61_0 = p_2_61 << 1;
  assign t_r3_c61_1 = p_3_60 << 1;
  assign t_r3_c61_2 = p_3_61 << 2;
  assign t_r3_c61_3 = p_3_62 << 1;
  assign t_r3_c61_4 = p_4_61 << 1;
  assign t_r3_c61_5 = t_r3_c61_0 + p_2_60;
  assign t_r3_c61_6 = t_r3_c61_1 + p_2_62;
  assign t_r3_c61_7 = t_r3_c61_2 + t_r3_c61_3;
  assign t_r3_c61_8 = t_r3_c61_4 + p_4_60;
  assign t_r3_c61_9 = t_r3_c61_5 + t_r3_c61_6;
  assign t_r3_c61_10 = t_r3_c61_7 + t_r3_c61_8;
  assign t_r3_c61_11 = t_r3_c61_9 + t_r3_c61_10;
  assign t_r3_c61_12 = t_r3_c61_11 + p_4_62;
  assign out_3_61 = t_r3_c61_12 >> 4;

  assign t_r3_c62_0 = p_2_62 << 1;
  assign t_r3_c62_1 = p_3_61 << 1;
  assign t_r3_c62_2 = p_3_62 << 2;
  assign t_r3_c62_3 = p_3_63 << 1;
  assign t_r3_c62_4 = p_4_62 << 1;
  assign t_r3_c62_5 = t_r3_c62_0 + p_2_61;
  assign t_r3_c62_6 = t_r3_c62_1 + p_2_63;
  assign t_r3_c62_7 = t_r3_c62_2 + t_r3_c62_3;
  assign t_r3_c62_8 = t_r3_c62_4 + p_4_61;
  assign t_r3_c62_9 = t_r3_c62_5 + t_r3_c62_6;
  assign t_r3_c62_10 = t_r3_c62_7 + t_r3_c62_8;
  assign t_r3_c62_11 = t_r3_c62_9 + t_r3_c62_10;
  assign t_r3_c62_12 = t_r3_c62_11 + p_4_63;
  assign out_3_62 = t_r3_c62_12 >> 4;

  assign t_r3_c63_0 = p_2_63 << 1;
  assign t_r3_c63_1 = p_3_62 << 1;
  assign t_r3_c63_2 = p_3_63 << 2;
  assign t_r3_c63_3 = p_3_64 << 1;
  assign t_r3_c63_4 = p_4_63 << 1;
  assign t_r3_c63_5 = t_r3_c63_0 + p_2_62;
  assign t_r3_c63_6 = t_r3_c63_1 + p_2_64;
  assign t_r3_c63_7 = t_r3_c63_2 + t_r3_c63_3;
  assign t_r3_c63_8 = t_r3_c63_4 + p_4_62;
  assign t_r3_c63_9 = t_r3_c63_5 + t_r3_c63_6;
  assign t_r3_c63_10 = t_r3_c63_7 + t_r3_c63_8;
  assign t_r3_c63_11 = t_r3_c63_9 + t_r3_c63_10;
  assign t_r3_c63_12 = t_r3_c63_11 + p_4_64;
  assign out_3_63 = t_r3_c63_12 >> 4;

  assign t_r3_c64_0 = p_2_64 << 1;
  assign t_r3_c64_1 = p_3_63 << 1;
  assign t_r3_c64_2 = p_3_64 << 2;
  assign t_r3_c64_3 = p_3_65 << 1;
  assign t_r3_c64_4 = p_4_64 << 1;
  assign t_r3_c64_5 = t_r3_c64_0 + p_2_63;
  assign t_r3_c64_6 = t_r3_c64_1 + p_2_65;
  assign t_r3_c64_7 = t_r3_c64_2 + t_r3_c64_3;
  assign t_r3_c64_8 = t_r3_c64_4 + p_4_63;
  assign t_r3_c64_9 = t_r3_c64_5 + t_r3_c64_6;
  assign t_r3_c64_10 = t_r3_c64_7 + t_r3_c64_8;
  assign t_r3_c64_11 = t_r3_c64_9 + t_r3_c64_10;
  assign t_r3_c64_12 = t_r3_c64_11 + p_4_65;
  assign out_3_64 = t_r3_c64_12 >> 4;

  assign t_r4_c1_0 = p_3_1 << 1;
  assign t_r4_c1_1 = p_4_0 << 1;
  assign t_r4_c1_2 = p_4_1 << 2;
  assign t_r4_c1_3 = p_4_2 << 1;
  assign t_r4_c1_4 = p_5_1 << 1;
  assign t_r4_c1_5 = t_r4_c1_0 + p_3_0;
  assign t_r4_c1_6 = t_r4_c1_1 + p_3_2;
  assign t_r4_c1_7 = t_r4_c1_2 + t_r4_c1_3;
  assign t_r4_c1_8 = t_r4_c1_4 + p_5_0;
  assign t_r4_c1_9 = t_r4_c1_5 + t_r4_c1_6;
  assign t_r4_c1_10 = t_r4_c1_7 + t_r4_c1_8;
  assign t_r4_c1_11 = t_r4_c1_9 + t_r4_c1_10;
  assign t_r4_c1_12 = t_r4_c1_11 + p_5_2;
  assign out_4_1 = t_r4_c1_12 >> 4;

  assign t_r4_c2_0 = p_3_2 << 1;
  assign t_r4_c2_1 = p_4_1 << 1;
  assign t_r4_c2_2 = p_4_2 << 2;
  assign t_r4_c2_3 = p_4_3 << 1;
  assign t_r4_c2_4 = p_5_2 << 1;
  assign t_r4_c2_5 = t_r4_c2_0 + p_3_1;
  assign t_r4_c2_6 = t_r4_c2_1 + p_3_3;
  assign t_r4_c2_7 = t_r4_c2_2 + t_r4_c2_3;
  assign t_r4_c2_8 = t_r4_c2_4 + p_5_1;
  assign t_r4_c2_9 = t_r4_c2_5 + t_r4_c2_6;
  assign t_r4_c2_10 = t_r4_c2_7 + t_r4_c2_8;
  assign t_r4_c2_11 = t_r4_c2_9 + t_r4_c2_10;
  assign t_r4_c2_12 = t_r4_c2_11 + p_5_3;
  assign out_4_2 = t_r4_c2_12 >> 4;

  assign t_r4_c3_0 = p_3_3 << 1;
  assign t_r4_c3_1 = p_4_2 << 1;
  assign t_r4_c3_2 = p_4_3 << 2;
  assign t_r4_c3_3 = p_4_4 << 1;
  assign t_r4_c3_4 = p_5_3 << 1;
  assign t_r4_c3_5 = t_r4_c3_0 + p_3_2;
  assign t_r4_c3_6 = t_r4_c3_1 + p_3_4;
  assign t_r4_c3_7 = t_r4_c3_2 + t_r4_c3_3;
  assign t_r4_c3_8 = t_r4_c3_4 + p_5_2;
  assign t_r4_c3_9 = t_r4_c3_5 + t_r4_c3_6;
  assign t_r4_c3_10 = t_r4_c3_7 + t_r4_c3_8;
  assign t_r4_c3_11 = t_r4_c3_9 + t_r4_c3_10;
  assign t_r4_c3_12 = t_r4_c3_11 + p_5_4;
  assign out_4_3 = t_r4_c3_12 >> 4;

  assign t_r4_c4_0 = p_3_4 << 1;
  assign t_r4_c4_1 = p_4_3 << 1;
  assign t_r4_c4_2 = p_4_4 << 2;
  assign t_r4_c4_3 = p_4_5 << 1;
  assign t_r4_c4_4 = p_5_4 << 1;
  assign t_r4_c4_5 = t_r4_c4_0 + p_3_3;
  assign t_r4_c4_6 = t_r4_c4_1 + p_3_5;
  assign t_r4_c4_7 = t_r4_c4_2 + t_r4_c4_3;
  assign t_r4_c4_8 = t_r4_c4_4 + p_5_3;
  assign t_r4_c4_9 = t_r4_c4_5 + t_r4_c4_6;
  assign t_r4_c4_10 = t_r4_c4_7 + t_r4_c4_8;
  assign t_r4_c4_11 = t_r4_c4_9 + t_r4_c4_10;
  assign t_r4_c4_12 = t_r4_c4_11 + p_5_5;
  assign out_4_4 = t_r4_c4_12 >> 4;

  assign t_r4_c5_0 = p_3_5 << 1;
  assign t_r4_c5_1 = p_4_4 << 1;
  assign t_r4_c5_2 = p_4_5 << 2;
  assign t_r4_c5_3 = p_4_6 << 1;
  assign t_r4_c5_4 = p_5_5 << 1;
  assign t_r4_c5_5 = t_r4_c5_0 + p_3_4;
  assign t_r4_c5_6 = t_r4_c5_1 + p_3_6;
  assign t_r4_c5_7 = t_r4_c5_2 + t_r4_c5_3;
  assign t_r4_c5_8 = t_r4_c5_4 + p_5_4;
  assign t_r4_c5_9 = t_r4_c5_5 + t_r4_c5_6;
  assign t_r4_c5_10 = t_r4_c5_7 + t_r4_c5_8;
  assign t_r4_c5_11 = t_r4_c5_9 + t_r4_c5_10;
  assign t_r4_c5_12 = t_r4_c5_11 + p_5_6;
  assign out_4_5 = t_r4_c5_12 >> 4;

  assign t_r4_c6_0 = p_3_6 << 1;
  assign t_r4_c6_1 = p_4_5 << 1;
  assign t_r4_c6_2 = p_4_6 << 2;
  assign t_r4_c6_3 = p_4_7 << 1;
  assign t_r4_c6_4 = p_5_6 << 1;
  assign t_r4_c6_5 = t_r4_c6_0 + p_3_5;
  assign t_r4_c6_6 = t_r4_c6_1 + p_3_7;
  assign t_r4_c6_7 = t_r4_c6_2 + t_r4_c6_3;
  assign t_r4_c6_8 = t_r4_c6_4 + p_5_5;
  assign t_r4_c6_9 = t_r4_c6_5 + t_r4_c6_6;
  assign t_r4_c6_10 = t_r4_c6_7 + t_r4_c6_8;
  assign t_r4_c6_11 = t_r4_c6_9 + t_r4_c6_10;
  assign t_r4_c6_12 = t_r4_c6_11 + p_5_7;
  assign out_4_6 = t_r4_c6_12 >> 4;

  assign t_r4_c7_0 = p_3_7 << 1;
  assign t_r4_c7_1 = p_4_6 << 1;
  assign t_r4_c7_2 = p_4_7 << 2;
  assign t_r4_c7_3 = p_4_8 << 1;
  assign t_r4_c7_4 = p_5_7 << 1;
  assign t_r4_c7_5 = t_r4_c7_0 + p_3_6;
  assign t_r4_c7_6 = t_r4_c7_1 + p_3_8;
  assign t_r4_c7_7 = t_r4_c7_2 + t_r4_c7_3;
  assign t_r4_c7_8 = t_r4_c7_4 + p_5_6;
  assign t_r4_c7_9 = t_r4_c7_5 + t_r4_c7_6;
  assign t_r4_c7_10 = t_r4_c7_7 + t_r4_c7_8;
  assign t_r4_c7_11 = t_r4_c7_9 + t_r4_c7_10;
  assign t_r4_c7_12 = t_r4_c7_11 + p_5_8;
  assign out_4_7 = t_r4_c7_12 >> 4;

  assign t_r4_c8_0 = p_3_8 << 1;
  assign t_r4_c8_1 = p_4_7 << 1;
  assign t_r4_c8_2 = p_4_8 << 2;
  assign t_r4_c8_3 = p_4_9 << 1;
  assign t_r4_c8_4 = p_5_8 << 1;
  assign t_r4_c8_5 = t_r4_c8_0 + p_3_7;
  assign t_r4_c8_6 = t_r4_c8_1 + p_3_9;
  assign t_r4_c8_7 = t_r4_c8_2 + t_r4_c8_3;
  assign t_r4_c8_8 = t_r4_c8_4 + p_5_7;
  assign t_r4_c8_9 = t_r4_c8_5 + t_r4_c8_6;
  assign t_r4_c8_10 = t_r4_c8_7 + t_r4_c8_8;
  assign t_r4_c8_11 = t_r4_c8_9 + t_r4_c8_10;
  assign t_r4_c8_12 = t_r4_c8_11 + p_5_9;
  assign out_4_8 = t_r4_c8_12 >> 4;

  assign t_r4_c9_0 = p_3_9 << 1;
  assign t_r4_c9_1 = p_4_8 << 1;
  assign t_r4_c9_2 = p_4_9 << 2;
  assign t_r4_c9_3 = p_4_10 << 1;
  assign t_r4_c9_4 = p_5_9 << 1;
  assign t_r4_c9_5 = t_r4_c9_0 + p_3_8;
  assign t_r4_c9_6 = t_r4_c9_1 + p_3_10;
  assign t_r4_c9_7 = t_r4_c9_2 + t_r4_c9_3;
  assign t_r4_c9_8 = t_r4_c9_4 + p_5_8;
  assign t_r4_c9_9 = t_r4_c9_5 + t_r4_c9_6;
  assign t_r4_c9_10 = t_r4_c9_7 + t_r4_c9_8;
  assign t_r4_c9_11 = t_r4_c9_9 + t_r4_c9_10;
  assign t_r4_c9_12 = t_r4_c9_11 + p_5_10;
  assign out_4_9 = t_r4_c9_12 >> 4;

  assign t_r4_c10_0 = p_3_10 << 1;
  assign t_r4_c10_1 = p_4_9 << 1;
  assign t_r4_c10_2 = p_4_10 << 2;
  assign t_r4_c10_3 = p_4_11 << 1;
  assign t_r4_c10_4 = p_5_10 << 1;
  assign t_r4_c10_5 = t_r4_c10_0 + p_3_9;
  assign t_r4_c10_6 = t_r4_c10_1 + p_3_11;
  assign t_r4_c10_7 = t_r4_c10_2 + t_r4_c10_3;
  assign t_r4_c10_8 = t_r4_c10_4 + p_5_9;
  assign t_r4_c10_9 = t_r4_c10_5 + t_r4_c10_6;
  assign t_r4_c10_10 = t_r4_c10_7 + t_r4_c10_8;
  assign t_r4_c10_11 = t_r4_c10_9 + t_r4_c10_10;
  assign t_r4_c10_12 = t_r4_c10_11 + p_5_11;
  assign out_4_10 = t_r4_c10_12 >> 4;

  assign t_r4_c11_0 = p_3_11 << 1;
  assign t_r4_c11_1 = p_4_10 << 1;
  assign t_r4_c11_2 = p_4_11 << 2;
  assign t_r4_c11_3 = p_4_12 << 1;
  assign t_r4_c11_4 = p_5_11 << 1;
  assign t_r4_c11_5 = t_r4_c11_0 + p_3_10;
  assign t_r4_c11_6 = t_r4_c11_1 + p_3_12;
  assign t_r4_c11_7 = t_r4_c11_2 + t_r4_c11_3;
  assign t_r4_c11_8 = t_r4_c11_4 + p_5_10;
  assign t_r4_c11_9 = t_r4_c11_5 + t_r4_c11_6;
  assign t_r4_c11_10 = t_r4_c11_7 + t_r4_c11_8;
  assign t_r4_c11_11 = t_r4_c11_9 + t_r4_c11_10;
  assign t_r4_c11_12 = t_r4_c11_11 + p_5_12;
  assign out_4_11 = t_r4_c11_12 >> 4;

  assign t_r4_c12_0 = p_3_12 << 1;
  assign t_r4_c12_1 = p_4_11 << 1;
  assign t_r4_c12_2 = p_4_12 << 2;
  assign t_r4_c12_3 = p_4_13 << 1;
  assign t_r4_c12_4 = p_5_12 << 1;
  assign t_r4_c12_5 = t_r4_c12_0 + p_3_11;
  assign t_r4_c12_6 = t_r4_c12_1 + p_3_13;
  assign t_r4_c12_7 = t_r4_c12_2 + t_r4_c12_3;
  assign t_r4_c12_8 = t_r4_c12_4 + p_5_11;
  assign t_r4_c12_9 = t_r4_c12_5 + t_r4_c12_6;
  assign t_r4_c12_10 = t_r4_c12_7 + t_r4_c12_8;
  assign t_r4_c12_11 = t_r4_c12_9 + t_r4_c12_10;
  assign t_r4_c12_12 = t_r4_c12_11 + p_5_13;
  assign out_4_12 = t_r4_c12_12 >> 4;

  assign t_r4_c13_0 = p_3_13 << 1;
  assign t_r4_c13_1 = p_4_12 << 1;
  assign t_r4_c13_2 = p_4_13 << 2;
  assign t_r4_c13_3 = p_4_14 << 1;
  assign t_r4_c13_4 = p_5_13 << 1;
  assign t_r4_c13_5 = t_r4_c13_0 + p_3_12;
  assign t_r4_c13_6 = t_r4_c13_1 + p_3_14;
  assign t_r4_c13_7 = t_r4_c13_2 + t_r4_c13_3;
  assign t_r4_c13_8 = t_r4_c13_4 + p_5_12;
  assign t_r4_c13_9 = t_r4_c13_5 + t_r4_c13_6;
  assign t_r4_c13_10 = t_r4_c13_7 + t_r4_c13_8;
  assign t_r4_c13_11 = t_r4_c13_9 + t_r4_c13_10;
  assign t_r4_c13_12 = t_r4_c13_11 + p_5_14;
  assign out_4_13 = t_r4_c13_12 >> 4;

  assign t_r4_c14_0 = p_3_14 << 1;
  assign t_r4_c14_1 = p_4_13 << 1;
  assign t_r4_c14_2 = p_4_14 << 2;
  assign t_r4_c14_3 = p_4_15 << 1;
  assign t_r4_c14_4 = p_5_14 << 1;
  assign t_r4_c14_5 = t_r4_c14_0 + p_3_13;
  assign t_r4_c14_6 = t_r4_c14_1 + p_3_15;
  assign t_r4_c14_7 = t_r4_c14_2 + t_r4_c14_3;
  assign t_r4_c14_8 = t_r4_c14_4 + p_5_13;
  assign t_r4_c14_9 = t_r4_c14_5 + t_r4_c14_6;
  assign t_r4_c14_10 = t_r4_c14_7 + t_r4_c14_8;
  assign t_r4_c14_11 = t_r4_c14_9 + t_r4_c14_10;
  assign t_r4_c14_12 = t_r4_c14_11 + p_5_15;
  assign out_4_14 = t_r4_c14_12 >> 4;

  assign t_r4_c15_0 = p_3_15 << 1;
  assign t_r4_c15_1 = p_4_14 << 1;
  assign t_r4_c15_2 = p_4_15 << 2;
  assign t_r4_c15_3 = p_4_16 << 1;
  assign t_r4_c15_4 = p_5_15 << 1;
  assign t_r4_c15_5 = t_r4_c15_0 + p_3_14;
  assign t_r4_c15_6 = t_r4_c15_1 + p_3_16;
  assign t_r4_c15_7 = t_r4_c15_2 + t_r4_c15_3;
  assign t_r4_c15_8 = t_r4_c15_4 + p_5_14;
  assign t_r4_c15_9 = t_r4_c15_5 + t_r4_c15_6;
  assign t_r4_c15_10 = t_r4_c15_7 + t_r4_c15_8;
  assign t_r4_c15_11 = t_r4_c15_9 + t_r4_c15_10;
  assign t_r4_c15_12 = t_r4_c15_11 + p_5_16;
  assign out_4_15 = t_r4_c15_12 >> 4;

  assign t_r4_c16_0 = p_3_16 << 1;
  assign t_r4_c16_1 = p_4_15 << 1;
  assign t_r4_c16_2 = p_4_16 << 2;
  assign t_r4_c16_3 = p_4_17 << 1;
  assign t_r4_c16_4 = p_5_16 << 1;
  assign t_r4_c16_5 = t_r4_c16_0 + p_3_15;
  assign t_r4_c16_6 = t_r4_c16_1 + p_3_17;
  assign t_r4_c16_7 = t_r4_c16_2 + t_r4_c16_3;
  assign t_r4_c16_8 = t_r4_c16_4 + p_5_15;
  assign t_r4_c16_9 = t_r4_c16_5 + t_r4_c16_6;
  assign t_r4_c16_10 = t_r4_c16_7 + t_r4_c16_8;
  assign t_r4_c16_11 = t_r4_c16_9 + t_r4_c16_10;
  assign t_r4_c16_12 = t_r4_c16_11 + p_5_17;
  assign out_4_16 = t_r4_c16_12 >> 4;

  assign t_r4_c17_0 = p_3_17 << 1;
  assign t_r4_c17_1 = p_4_16 << 1;
  assign t_r4_c17_2 = p_4_17 << 2;
  assign t_r4_c17_3 = p_4_18 << 1;
  assign t_r4_c17_4 = p_5_17 << 1;
  assign t_r4_c17_5 = t_r4_c17_0 + p_3_16;
  assign t_r4_c17_6 = t_r4_c17_1 + p_3_18;
  assign t_r4_c17_7 = t_r4_c17_2 + t_r4_c17_3;
  assign t_r4_c17_8 = t_r4_c17_4 + p_5_16;
  assign t_r4_c17_9 = t_r4_c17_5 + t_r4_c17_6;
  assign t_r4_c17_10 = t_r4_c17_7 + t_r4_c17_8;
  assign t_r4_c17_11 = t_r4_c17_9 + t_r4_c17_10;
  assign t_r4_c17_12 = t_r4_c17_11 + p_5_18;
  assign out_4_17 = t_r4_c17_12 >> 4;

  assign t_r4_c18_0 = p_3_18 << 1;
  assign t_r4_c18_1 = p_4_17 << 1;
  assign t_r4_c18_2 = p_4_18 << 2;
  assign t_r4_c18_3 = p_4_19 << 1;
  assign t_r4_c18_4 = p_5_18 << 1;
  assign t_r4_c18_5 = t_r4_c18_0 + p_3_17;
  assign t_r4_c18_6 = t_r4_c18_1 + p_3_19;
  assign t_r4_c18_7 = t_r4_c18_2 + t_r4_c18_3;
  assign t_r4_c18_8 = t_r4_c18_4 + p_5_17;
  assign t_r4_c18_9 = t_r4_c18_5 + t_r4_c18_6;
  assign t_r4_c18_10 = t_r4_c18_7 + t_r4_c18_8;
  assign t_r4_c18_11 = t_r4_c18_9 + t_r4_c18_10;
  assign t_r4_c18_12 = t_r4_c18_11 + p_5_19;
  assign out_4_18 = t_r4_c18_12 >> 4;

  assign t_r4_c19_0 = p_3_19 << 1;
  assign t_r4_c19_1 = p_4_18 << 1;
  assign t_r4_c19_2 = p_4_19 << 2;
  assign t_r4_c19_3 = p_4_20 << 1;
  assign t_r4_c19_4 = p_5_19 << 1;
  assign t_r4_c19_5 = t_r4_c19_0 + p_3_18;
  assign t_r4_c19_6 = t_r4_c19_1 + p_3_20;
  assign t_r4_c19_7 = t_r4_c19_2 + t_r4_c19_3;
  assign t_r4_c19_8 = t_r4_c19_4 + p_5_18;
  assign t_r4_c19_9 = t_r4_c19_5 + t_r4_c19_6;
  assign t_r4_c19_10 = t_r4_c19_7 + t_r4_c19_8;
  assign t_r4_c19_11 = t_r4_c19_9 + t_r4_c19_10;
  assign t_r4_c19_12 = t_r4_c19_11 + p_5_20;
  assign out_4_19 = t_r4_c19_12 >> 4;

  assign t_r4_c20_0 = p_3_20 << 1;
  assign t_r4_c20_1 = p_4_19 << 1;
  assign t_r4_c20_2 = p_4_20 << 2;
  assign t_r4_c20_3 = p_4_21 << 1;
  assign t_r4_c20_4 = p_5_20 << 1;
  assign t_r4_c20_5 = t_r4_c20_0 + p_3_19;
  assign t_r4_c20_6 = t_r4_c20_1 + p_3_21;
  assign t_r4_c20_7 = t_r4_c20_2 + t_r4_c20_3;
  assign t_r4_c20_8 = t_r4_c20_4 + p_5_19;
  assign t_r4_c20_9 = t_r4_c20_5 + t_r4_c20_6;
  assign t_r4_c20_10 = t_r4_c20_7 + t_r4_c20_8;
  assign t_r4_c20_11 = t_r4_c20_9 + t_r4_c20_10;
  assign t_r4_c20_12 = t_r4_c20_11 + p_5_21;
  assign out_4_20 = t_r4_c20_12 >> 4;

  assign t_r4_c21_0 = p_3_21 << 1;
  assign t_r4_c21_1 = p_4_20 << 1;
  assign t_r4_c21_2 = p_4_21 << 2;
  assign t_r4_c21_3 = p_4_22 << 1;
  assign t_r4_c21_4 = p_5_21 << 1;
  assign t_r4_c21_5 = t_r4_c21_0 + p_3_20;
  assign t_r4_c21_6 = t_r4_c21_1 + p_3_22;
  assign t_r4_c21_7 = t_r4_c21_2 + t_r4_c21_3;
  assign t_r4_c21_8 = t_r4_c21_4 + p_5_20;
  assign t_r4_c21_9 = t_r4_c21_5 + t_r4_c21_6;
  assign t_r4_c21_10 = t_r4_c21_7 + t_r4_c21_8;
  assign t_r4_c21_11 = t_r4_c21_9 + t_r4_c21_10;
  assign t_r4_c21_12 = t_r4_c21_11 + p_5_22;
  assign out_4_21 = t_r4_c21_12 >> 4;

  assign t_r4_c22_0 = p_3_22 << 1;
  assign t_r4_c22_1 = p_4_21 << 1;
  assign t_r4_c22_2 = p_4_22 << 2;
  assign t_r4_c22_3 = p_4_23 << 1;
  assign t_r4_c22_4 = p_5_22 << 1;
  assign t_r4_c22_5 = t_r4_c22_0 + p_3_21;
  assign t_r4_c22_6 = t_r4_c22_1 + p_3_23;
  assign t_r4_c22_7 = t_r4_c22_2 + t_r4_c22_3;
  assign t_r4_c22_8 = t_r4_c22_4 + p_5_21;
  assign t_r4_c22_9 = t_r4_c22_5 + t_r4_c22_6;
  assign t_r4_c22_10 = t_r4_c22_7 + t_r4_c22_8;
  assign t_r4_c22_11 = t_r4_c22_9 + t_r4_c22_10;
  assign t_r4_c22_12 = t_r4_c22_11 + p_5_23;
  assign out_4_22 = t_r4_c22_12 >> 4;

  assign t_r4_c23_0 = p_3_23 << 1;
  assign t_r4_c23_1 = p_4_22 << 1;
  assign t_r4_c23_2 = p_4_23 << 2;
  assign t_r4_c23_3 = p_4_24 << 1;
  assign t_r4_c23_4 = p_5_23 << 1;
  assign t_r4_c23_5 = t_r4_c23_0 + p_3_22;
  assign t_r4_c23_6 = t_r4_c23_1 + p_3_24;
  assign t_r4_c23_7 = t_r4_c23_2 + t_r4_c23_3;
  assign t_r4_c23_8 = t_r4_c23_4 + p_5_22;
  assign t_r4_c23_9 = t_r4_c23_5 + t_r4_c23_6;
  assign t_r4_c23_10 = t_r4_c23_7 + t_r4_c23_8;
  assign t_r4_c23_11 = t_r4_c23_9 + t_r4_c23_10;
  assign t_r4_c23_12 = t_r4_c23_11 + p_5_24;
  assign out_4_23 = t_r4_c23_12 >> 4;

  assign t_r4_c24_0 = p_3_24 << 1;
  assign t_r4_c24_1 = p_4_23 << 1;
  assign t_r4_c24_2 = p_4_24 << 2;
  assign t_r4_c24_3 = p_4_25 << 1;
  assign t_r4_c24_4 = p_5_24 << 1;
  assign t_r4_c24_5 = t_r4_c24_0 + p_3_23;
  assign t_r4_c24_6 = t_r4_c24_1 + p_3_25;
  assign t_r4_c24_7 = t_r4_c24_2 + t_r4_c24_3;
  assign t_r4_c24_8 = t_r4_c24_4 + p_5_23;
  assign t_r4_c24_9 = t_r4_c24_5 + t_r4_c24_6;
  assign t_r4_c24_10 = t_r4_c24_7 + t_r4_c24_8;
  assign t_r4_c24_11 = t_r4_c24_9 + t_r4_c24_10;
  assign t_r4_c24_12 = t_r4_c24_11 + p_5_25;
  assign out_4_24 = t_r4_c24_12 >> 4;

  assign t_r4_c25_0 = p_3_25 << 1;
  assign t_r4_c25_1 = p_4_24 << 1;
  assign t_r4_c25_2 = p_4_25 << 2;
  assign t_r4_c25_3 = p_4_26 << 1;
  assign t_r4_c25_4 = p_5_25 << 1;
  assign t_r4_c25_5 = t_r4_c25_0 + p_3_24;
  assign t_r4_c25_6 = t_r4_c25_1 + p_3_26;
  assign t_r4_c25_7 = t_r4_c25_2 + t_r4_c25_3;
  assign t_r4_c25_8 = t_r4_c25_4 + p_5_24;
  assign t_r4_c25_9 = t_r4_c25_5 + t_r4_c25_6;
  assign t_r4_c25_10 = t_r4_c25_7 + t_r4_c25_8;
  assign t_r4_c25_11 = t_r4_c25_9 + t_r4_c25_10;
  assign t_r4_c25_12 = t_r4_c25_11 + p_5_26;
  assign out_4_25 = t_r4_c25_12 >> 4;

  assign t_r4_c26_0 = p_3_26 << 1;
  assign t_r4_c26_1 = p_4_25 << 1;
  assign t_r4_c26_2 = p_4_26 << 2;
  assign t_r4_c26_3 = p_4_27 << 1;
  assign t_r4_c26_4 = p_5_26 << 1;
  assign t_r4_c26_5 = t_r4_c26_0 + p_3_25;
  assign t_r4_c26_6 = t_r4_c26_1 + p_3_27;
  assign t_r4_c26_7 = t_r4_c26_2 + t_r4_c26_3;
  assign t_r4_c26_8 = t_r4_c26_4 + p_5_25;
  assign t_r4_c26_9 = t_r4_c26_5 + t_r4_c26_6;
  assign t_r4_c26_10 = t_r4_c26_7 + t_r4_c26_8;
  assign t_r4_c26_11 = t_r4_c26_9 + t_r4_c26_10;
  assign t_r4_c26_12 = t_r4_c26_11 + p_5_27;
  assign out_4_26 = t_r4_c26_12 >> 4;

  assign t_r4_c27_0 = p_3_27 << 1;
  assign t_r4_c27_1 = p_4_26 << 1;
  assign t_r4_c27_2 = p_4_27 << 2;
  assign t_r4_c27_3 = p_4_28 << 1;
  assign t_r4_c27_4 = p_5_27 << 1;
  assign t_r4_c27_5 = t_r4_c27_0 + p_3_26;
  assign t_r4_c27_6 = t_r4_c27_1 + p_3_28;
  assign t_r4_c27_7 = t_r4_c27_2 + t_r4_c27_3;
  assign t_r4_c27_8 = t_r4_c27_4 + p_5_26;
  assign t_r4_c27_9 = t_r4_c27_5 + t_r4_c27_6;
  assign t_r4_c27_10 = t_r4_c27_7 + t_r4_c27_8;
  assign t_r4_c27_11 = t_r4_c27_9 + t_r4_c27_10;
  assign t_r4_c27_12 = t_r4_c27_11 + p_5_28;
  assign out_4_27 = t_r4_c27_12 >> 4;

  assign t_r4_c28_0 = p_3_28 << 1;
  assign t_r4_c28_1 = p_4_27 << 1;
  assign t_r4_c28_2 = p_4_28 << 2;
  assign t_r4_c28_3 = p_4_29 << 1;
  assign t_r4_c28_4 = p_5_28 << 1;
  assign t_r4_c28_5 = t_r4_c28_0 + p_3_27;
  assign t_r4_c28_6 = t_r4_c28_1 + p_3_29;
  assign t_r4_c28_7 = t_r4_c28_2 + t_r4_c28_3;
  assign t_r4_c28_8 = t_r4_c28_4 + p_5_27;
  assign t_r4_c28_9 = t_r4_c28_5 + t_r4_c28_6;
  assign t_r4_c28_10 = t_r4_c28_7 + t_r4_c28_8;
  assign t_r4_c28_11 = t_r4_c28_9 + t_r4_c28_10;
  assign t_r4_c28_12 = t_r4_c28_11 + p_5_29;
  assign out_4_28 = t_r4_c28_12 >> 4;

  assign t_r4_c29_0 = p_3_29 << 1;
  assign t_r4_c29_1 = p_4_28 << 1;
  assign t_r4_c29_2 = p_4_29 << 2;
  assign t_r4_c29_3 = p_4_30 << 1;
  assign t_r4_c29_4 = p_5_29 << 1;
  assign t_r4_c29_5 = t_r4_c29_0 + p_3_28;
  assign t_r4_c29_6 = t_r4_c29_1 + p_3_30;
  assign t_r4_c29_7 = t_r4_c29_2 + t_r4_c29_3;
  assign t_r4_c29_8 = t_r4_c29_4 + p_5_28;
  assign t_r4_c29_9 = t_r4_c29_5 + t_r4_c29_6;
  assign t_r4_c29_10 = t_r4_c29_7 + t_r4_c29_8;
  assign t_r4_c29_11 = t_r4_c29_9 + t_r4_c29_10;
  assign t_r4_c29_12 = t_r4_c29_11 + p_5_30;
  assign out_4_29 = t_r4_c29_12 >> 4;

  assign t_r4_c30_0 = p_3_30 << 1;
  assign t_r4_c30_1 = p_4_29 << 1;
  assign t_r4_c30_2 = p_4_30 << 2;
  assign t_r4_c30_3 = p_4_31 << 1;
  assign t_r4_c30_4 = p_5_30 << 1;
  assign t_r4_c30_5 = t_r4_c30_0 + p_3_29;
  assign t_r4_c30_6 = t_r4_c30_1 + p_3_31;
  assign t_r4_c30_7 = t_r4_c30_2 + t_r4_c30_3;
  assign t_r4_c30_8 = t_r4_c30_4 + p_5_29;
  assign t_r4_c30_9 = t_r4_c30_5 + t_r4_c30_6;
  assign t_r4_c30_10 = t_r4_c30_7 + t_r4_c30_8;
  assign t_r4_c30_11 = t_r4_c30_9 + t_r4_c30_10;
  assign t_r4_c30_12 = t_r4_c30_11 + p_5_31;
  assign out_4_30 = t_r4_c30_12 >> 4;

  assign t_r4_c31_0 = p_3_31 << 1;
  assign t_r4_c31_1 = p_4_30 << 1;
  assign t_r4_c31_2 = p_4_31 << 2;
  assign t_r4_c31_3 = p_4_32 << 1;
  assign t_r4_c31_4 = p_5_31 << 1;
  assign t_r4_c31_5 = t_r4_c31_0 + p_3_30;
  assign t_r4_c31_6 = t_r4_c31_1 + p_3_32;
  assign t_r4_c31_7 = t_r4_c31_2 + t_r4_c31_3;
  assign t_r4_c31_8 = t_r4_c31_4 + p_5_30;
  assign t_r4_c31_9 = t_r4_c31_5 + t_r4_c31_6;
  assign t_r4_c31_10 = t_r4_c31_7 + t_r4_c31_8;
  assign t_r4_c31_11 = t_r4_c31_9 + t_r4_c31_10;
  assign t_r4_c31_12 = t_r4_c31_11 + p_5_32;
  assign out_4_31 = t_r4_c31_12 >> 4;

  assign t_r4_c32_0 = p_3_32 << 1;
  assign t_r4_c32_1 = p_4_31 << 1;
  assign t_r4_c32_2 = p_4_32 << 2;
  assign t_r4_c32_3 = p_4_33 << 1;
  assign t_r4_c32_4 = p_5_32 << 1;
  assign t_r4_c32_5 = t_r4_c32_0 + p_3_31;
  assign t_r4_c32_6 = t_r4_c32_1 + p_3_33;
  assign t_r4_c32_7 = t_r4_c32_2 + t_r4_c32_3;
  assign t_r4_c32_8 = t_r4_c32_4 + p_5_31;
  assign t_r4_c32_9 = t_r4_c32_5 + t_r4_c32_6;
  assign t_r4_c32_10 = t_r4_c32_7 + t_r4_c32_8;
  assign t_r4_c32_11 = t_r4_c32_9 + t_r4_c32_10;
  assign t_r4_c32_12 = t_r4_c32_11 + p_5_33;
  assign out_4_32 = t_r4_c32_12 >> 4;

  assign t_r4_c33_0 = p_3_33 << 1;
  assign t_r4_c33_1 = p_4_32 << 1;
  assign t_r4_c33_2 = p_4_33 << 2;
  assign t_r4_c33_3 = p_4_34 << 1;
  assign t_r4_c33_4 = p_5_33 << 1;
  assign t_r4_c33_5 = t_r4_c33_0 + p_3_32;
  assign t_r4_c33_6 = t_r4_c33_1 + p_3_34;
  assign t_r4_c33_7 = t_r4_c33_2 + t_r4_c33_3;
  assign t_r4_c33_8 = t_r4_c33_4 + p_5_32;
  assign t_r4_c33_9 = t_r4_c33_5 + t_r4_c33_6;
  assign t_r4_c33_10 = t_r4_c33_7 + t_r4_c33_8;
  assign t_r4_c33_11 = t_r4_c33_9 + t_r4_c33_10;
  assign t_r4_c33_12 = t_r4_c33_11 + p_5_34;
  assign out_4_33 = t_r4_c33_12 >> 4;

  assign t_r4_c34_0 = p_3_34 << 1;
  assign t_r4_c34_1 = p_4_33 << 1;
  assign t_r4_c34_2 = p_4_34 << 2;
  assign t_r4_c34_3 = p_4_35 << 1;
  assign t_r4_c34_4 = p_5_34 << 1;
  assign t_r4_c34_5 = t_r4_c34_0 + p_3_33;
  assign t_r4_c34_6 = t_r4_c34_1 + p_3_35;
  assign t_r4_c34_7 = t_r4_c34_2 + t_r4_c34_3;
  assign t_r4_c34_8 = t_r4_c34_4 + p_5_33;
  assign t_r4_c34_9 = t_r4_c34_5 + t_r4_c34_6;
  assign t_r4_c34_10 = t_r4_c34_7 + t_r4_c34_8;
  assign t_r4_c34_11 = t_r4_c34_9 + t_r4_c34_10;
  assign t_r4_c34_12 = t_r4_c34_11 + p_5_35;
  assign out_4_34 = t_r4_c34_12 >> 4;

  assign t_r4_c35_0 = p_3_35 << 1;
  assign t_r4_c35_1 = p_4_34 << 1;
  assign t_r4_c35_2 = p_4_35 << 2;
  assign t_r4_c35_3 = p_4_36 << 1;
  assign t_r4_c35_4 = p_5_35 << 1;
  assign t_r4_c35_5 = t_r4_c35_0 + p_3_34;
  assign t_r4_c35_6 = t_r4_c35_1 + p_3_36;
  assign t_r4_c35_7 = t_r4_c35_2 + t_r4_c35_3;
  assign t_r4_c35_8 = t_r4_c35_4 + p_5_34;
  assign t_r4_c35_9 = t_r4_c35_5 + t_r4_c35_6;
  assign t_r4_c35_10 = t_r4_c35_7 + t_r4_c35_8;
  assign t_r4_c35_11 = t_r4_c35_9 + t_r4_c35_10;
  assign t_r4_c35_12 = t_r4_c35_11 + p_5_36;
  assign out_4_35 = t_r4_c35_12 >> 4;

  assign t_r4_c36_0 = p_3_36 << 1;
  assign t_r4_c36_1 = p_4_35 << 1;
  assign t_r4_c36_2 = p_4_36 << 2;
  assign t_r4_c36_3 = p_4_37 << 1;
  assign t_r4_c36_4 = p_5_36 << 1;
  assign t_r4_c36_5 = t_r4_c36_0 + p_3_35;
  assign t_r4_c36_6 = t_r4_c36_1 + p_3_37;
  assign t_r4_c36_7 = t_r4_c36_2 + t_r4_c36_3;
  assign t_r4_c36_8 = t_r4_c36_4 + p_5_35;
  assign t_r4_c36_9 = t_r4_c36_5 + t_r4_c36_6;
  assign t_r4_c36_10 = t_r4_c36_7 + t_r4_c36_8;
  assign t_r4_c36_11 = t_r4_c36_9 + t_r4_c36_10;
  assign t_r4_c36_12 = t_r4_c36_11 + p_5_37;
  assign out_4_36 = t_r4_c36_12 >> 4;

  assign t_r4_c37_0 = p_3_37 << 1;
  assign t_r4_c37_1 = p_4_36 << 1;
  assign t_r4_c37_2 = p_4_37 << 2;
  assign t_r4_c37_3 = p_4_38 << 1;
  assign t_r4_c37_4 = p_5_37 << 1;
  assign t_r4_c37_5 = t_r4_c37_0 + p_3_36;
  assign t_r4_c37_6 = t_r4_c37_1 + p_3_38;
  assign t_r4_c37_7 = t_r4_c37_2 + t_r4_c37_3;
  assign t_r4_c37_8 = t_r4_c37_4 + p_5_36;
  assign t_r4_c37_9 = t_r4_c37_5 + t_r4_c37_6;
  assign t_r4_c37_10 = t_r4_c37_7 + t_r4_c37_8;
  assign t_r4_c37_11 = t_r4_c37_9 + t_r4_c37_10;
  assign t_r4_c37_12 = t_r4_c37_11 + p_5_38;
  assign out_4_37 = t_r4_c37_12 >> 4;

  assign t_r4_c38_0 = p_3_38 << 1;
  assign t_r4_c38_1 = p_4_37 << 1;
  assign t_r4_c38_2 = p_4_38 << 2;
  assign t_r4_c38_3 = p_4_39 << 1;
  assign t_r4_c38_4 = p_5_38 << 1;
  assign t_r4_c38_5 = t_r4_c38_0 + p_3_37;
  assign t_r4_c38_6 = t_r4_c38_1 + p_3_39;
  assign t_r4_c38_7 = t_r4_c38_2 + t_r4_c38_3;
  assign t_r4_c38_8 = t_r4_c38_4 + p_5_37;
  assign t_r4_c38_9 = t_r4_c38_5 + t_r4_c38_6;
  assign t_r4_c38_10 = t_r4_c38_7 + t_r4_c38_8;
  assign t_r4_c38_11 = t_r4_c38_9 + t_r4_c38_10;
  assign t_r4_c38_12 = t_r4_c38_11 + p_5_39;
  assign out_4_38 = t_r4_c38_12 >> 4;

  assign t_r4_c39_0 = p_3_39 << 1;
  assign t_r4_c39_1 = p_4_38 << 1;
  assign t_r4_c39_2 = p_4_39 << 2;
  assign t_r4_c39_3 = p_4_40 << 1;
  assign t_r4_c39_4 = p_5_39 << 1;
  assign t_r4_c39_5 = t_r4_c39_0 + p_3_38;
  assign t_r4_c39_6 = t_r4_c39_1 + p_3_40;
  assign t_r4_c39_7 = t_r4_c39_2 + t_r4_c39_3;
  assign t_r4_c39_8 = t_r4_c39_4 + p_5_38;
  assign t_r4_c39_9 = t_r4_c39_5 + t_r4_c39_6;
  assign t_r4_c39_10 = t_r4_c39_7 + t_r4_c39_8;
  assign t_r4_c39_11 = t_r4_c39_9 + t_r4_c39_10;
  assign t_r4_c39_12 = t_r4_c39_11 + p_5_40;
  assign out_4_39 = t_r4_c39_12 >> 4;

  assign t_r4_c40_0 = p_3_40 << 1;
  assign t_r4_c40_1 = p_4_39 << 1;
  assign t_r4_c40_2 = p_4_40 << 2;
  assign t_r4_c40_3 = p_4_41 << 1;
  assign t_r4_c40_4 = p_5_40 << 1;
  assign t_r4_c40_5 = t_r4_c40_0 + p_3_39;
  assign t_r4_c40_6 = t_r4_c40_1 + p_3_41;
  assign t_r4_c40_7 = t_r4_c40_2 + t_r4_c40_3;
  assign t_r4_c40_8 = t_r4_c40_4 + p_5_39;
  assign t_r4_c40_9 = t_r4_c40_5 + t_r4_c40_6;
  assign t_r4_c40_10 = t_r4_c40_7 + t_r4_c40_8;
  assign t_r4_c40_11 = t_r4_c40_9 + t_r4_c40_10;
  assign t_r4_c40_12 = t_r4_c40_11 + p_5_41;
  assign out_4_40 = t_r4_c40_12 >> 4;

  assign t_r4_c41_0 = p_3_41 << 1;
  assign t_r4_c41_1 = p_4_40 << 1;
  assign t_r4_c41_2 = p_4_41 << 2;
  assign t_r4_c41_3 = p_4_42 << 1;
  assign t_r4_c41_4 = p_5_41 << 1;
  assign t_r4_c41_5 = t_r4_c41_0 + p_3_40;
  assign t_r4_c41_6 = t_r4_c41_1 + p_3_42;
  assign t_r4_c41_7 = t_r4_c41_2 + t_r4_c41_3;
  assign t_r4_c41_8 = t_r4_c41_4 + p_5_40;
  assign t_r4_c41_9 = t_r4_c41_5 + t_r4_c41_6;
  assign t_r4_c41_10 = t_r4_c41_7 + t_r4_c41_8;
  assign t_r4_c41_11 = t_r4_c41_9 + t_r4_c41_10;
  assign t_r4_c41_12 = t_r4_c41_11 + p_5_42;
  assign out_4_41 = t_r4_c41_12 >> 4;

  assign t_r4_c42_0 = p_3_42 << 1;
  assign t_r4_c42_1 = p_4_41 << 1;
  assign t_r4_c42_2 = p_4_42 << 2;
  assign t_r4_c42_3 = p_4_43 << 1;
  assign t_r4_c42_4 = p_5_42 << 1;
  assign t_r4_c42_5 = t_r4_c42_0 + p_3_41;
  assign t_r4_c42_6 = t_r4_c42_1 + p_3_43;
  assign t_r4_c42_7 = t_r4_c42_2 + t_r4_c42_3;
  assign t_r4_c42_8 = t_r4_c42_4 + p_5_41;
  assign t_r4_c42_9 = t_r4_c42_5 + t_r4_c42_6;
  assign t_r4_c42_10 = t_r4_c42_7 + t_r4_c42_8;
  assign t_r4_c42_11 = t_r4_c42_9 + t_r4_c42_10;
  assign t_r4_c42_12 = t_r4_c42_11 + p_5_43;
  assign out_4_42 = t_r4_c42_12 >> 4;

  assign t_r4_c43_0 = p_3_43 << 1;
  assign t_r4_c43_1 = p_4_42 << 1;
  assign t_r4_c43_2 = p_4_43 << 2;
  assign t_r4_c43_3 = p_4_44 << 1;
  assign t_r4_c43_4 = p_5_43 << 1;
  assign t_r4_c43_5 = t_r4_c43_0 + p_3_42;
  assign t_r4_c43_6 = t_r4_c43_1 + p_3_44;
  assign t_r4_c43_7 = t_r4_c43_2 + t_r4_c43_3;
  assign t_r4_c43_8 = t_r4_c43_4 + p_5_42;
  assign t_r4_c43_9 = t_r4_c43_5 + t_r4_c43_6;
  assign t_r4_c43_10 = t_r4_c43_7 + t_r4_c43_8;
  assign t_r4_c43_11 = t_r4_c43_9 + t_r4_c43_10;
  assign t_r4_c43_12 = t_r4_c43_11 + p_5_44;
  assign out_4_43 = t_r4_c43_12 >> 4;

  assign t_r4_c44_0 = p_3_44 << 1;
  assign t_r4_c44_1 = p_4_43 << 1;
  assign t_r4_c44_2 = p_4_44 << 2;
  assign t_r4_c44_3 = p_4_45 << 1;
  assign t_r4_c44_4 = p_5_44 << 1;
  assign t_r4_c44_5 = t_r4_c44_0 + p_3_43;
  assign t_r4_c44_6 = t_r4_c44_1 + p_3_45;
  assign t_r4_c44_7 = t_r4_c44_2 + t_r4_c44_3;
  assign t_r4_c44_8 = t_r4_c44_4 + p_5_43;
  assign t_r4_c44_9 = t_r4_c44_5 + t_r4_c44_6;
  assign t_r4_c44_10 = t_r4_c44_7 + t_r4_c44_8;
  assign t_r4_c44_11 = t_r4_c44_9 + t_r4_c44_10;
  assign t_r4_c44_12 = t_r4_c44_11 + p_5_45;
  assign out_4_44 = t_r4_c44_12 >> 4;

  assign t_r4_c45_0 = p_3_45 << 1;
  assign t_r4_c45_1 = p_4_44 << 1;
  assign t_r4_c45_2 = p_4_45 << 2;
  assign t_r4_c45_3 = p_4_46 << 1;
  assign t_r4_c45_4 = p_5_45 << 1;
  assign t_r4_c45_5 = t_r4_c45_0 + p_3_44;
  assign t_r4_c45_6 = t_r4_c45_1 + p_3_46;
  assign t_r4_c45_7 = t_r4_c45_2 + t_r4_c45_3;
  assign t_r4_c45_8 = t_r4_c45_4 + p_5_44;
  assign t_r4_c45_9 = t_r4_c45_5 + t_r4_c45_6;
  assign t_r4_c45_10 = t_r4_c45_7 + t_r4_c45_8;
  assign t_r4_c45_11 = t_r4_c45_9 + t_r4_c45_10;
  assign t_r4_c45_12 = t_r4_c45_11 + p_5_46;
  assign out_4_45 = t_r4_c45_12 >> 4;

  assign t_r4_c46_0 = p_3_46 << 1;
  assign t_r4_c46_1 = p_4_45 << 1;
  assign t_r4_c46_2 = p_4_46 << 2;
  assign t_r4_c46_3 = p_4_47 << 1;
  assign t_r4_c46_4 = p_5_46 << 1;
  assign t_r4_c46_5 = t_r4_c46_0 + p_3_45;
  assign t_r4_c46_6 = t_r4_c46_1 + p_3_47;
  assign t_r4_c46_7 = t_r4_c46_2 + t_r4_c46_3;
  assign t_r4_c46_8 = t_r4_c46_4 + p_5_45;
  assign t_r4_c46_9 = t_r4_c46_5 + t_r4_c46_6;
  assign t_r4_c46_10 = t_r4_c46_7 + t_r4_c46_8;
  assign t_r4_c46_11 = t_r4_c46_9 + t_r4_c46_10;
  assign t_r4_c46_12 = t_r4_c46_11 + p_5_47;
  assign out_4_46 = t_r4_c46_12 >> 4;

  assign t_r4_c47_0 = p_3_47 << 1;
  assign t_r4_c47_1 = p_4_46 << 1;
  assign t_r4_c47_2 = p_4_47 << 2;
  assign t_r4_c47_3 = p_4_48 << 1;
  assign t_r4_c47_4 = p_5_47 << 1;
  assign t_r4_c47_5 = t_r4_c47_0 + p_3_46;
  assign t_r4_c47_6 = t_r4_c47_1 + p_3_48;
  assign t_r4_c47_7 = t_r4_c47_2 + t_r4_c47_3;
  assign t_r4_c47_8 = t_r4_c47_4 + p_5_46;
  assign t_r4_c47_9 = t_r4_c47_5 + t_r4_c47_6;
  assign t_r4_c47_10 = t_r4_c47_7 + t_r4_c47_8;
  assign t_r4_c47_11 = t_r4_c47_9 + t_r4_c47_10;
  assign t_r4_c47_12 = t_r4_c47_11 + p_5_48;
  assign out_4_47 = t_r4_c47_12 >> 4;

  assign t_r4_c48_0 = p_3_48 << 1;
  assign t_r4_c48_1 = p_4_47 << 1;
  assign t_r4_c48_2 = p_4_48 << 2;
  assign t_r4_c48_3 = p_4_49 << 1;
  assign t_r4_c48_4 = p_5_48 << 1;
  assign t_r4_c48_5 = t_r4_c48_0 + p_3_47;
  assign t_r4_c48_6 = t_r4_c48_1 + p_3_49;
  assign t_r4_c48_7 = t_r4_c48_2 + t_r4_c48_3;
  assign t_r4_c48_8 = t_r4_c48_4 + p_5_47;
  assign t_r4_c48_9 = t_r4_c48_5 + t_r4_c48_6;
  assign t_r4_c48_10 = t_r4_c48_7 + t_r4_c48_8;
  assign t_r4_c48_11 = t_r4_c48_9 + t_r4_c48_10;
  assign t_r4_c48_12 = t_r4_c48_11 + p_5_49;
  assign out_4_48 = t_r4_c48_12 >> 4;

  assign t_r4_c49_0 = p_3_49 << 1;
  assign t_r4_c49_1 = p_4_48 << 1;
  assign t_r4_c49_2 = p_4_49 << 2;
  assign t_r4_c49_3 = p_4_50 << 1;
  assign t_r4_c49_4 = p_5_49 << 1;
  assign t_r4_c49_5 = t_r4_c49_0 + p_3_48;
  assign t_r4_c49_6 = t_r4_c49_1 + p_3_50;
  assign t_r4_c49_7 = t_r4_c49_2 + t_r4_c49_3;
  assign t_r4_c49_8 = t_r4_c49_4 + p_5_48;
  assign t_r4_c49_9 = t_r4_c49_5 + t_r4_c49_6;
  assign t_r4_c49_10 = t_r4_c49_7 + t_r4_c49_8;
  assign t_r4_c49_11 = t_r4_c49_9 + t_r4_c49_10;
  assign t_r4_c49_12 = t_r4_c49_11 + p_5_50;
  assign out_4_49 = t_r4_c49_12 >> 4;

  assign t_r4_c50_0 = p_3_50 << 1;
  assign t_r4_c50_1 = p_4_49 << 1;
  assign t_r4_c50_2 = p_4_50 << 2;
  assign t_r4_c50_3 = p_4_51 << 1;
  assign t_r4_c50_4 = p_5_50 << 1;
  assign t_r4_c50_5 = t_r4_c50_0 + p_3_49;
  assign t_r4_c50_6 = t_r4_c50_1 + p_3_51;
  assign t_r4_c50_7 = t_r4_c50_2 + t_r4_c50_3;
  assign t_r4_c50_8 = t_r4_c50_4 + p_5_49;
  assign t_r4_c50_9 = t_r4_c50_5 + t_r4_c50_6;
  assign t_r4_c50_10 = t_r4_c50_7 + t_r4_c50_8;
  assign t_r4_c50_11 = t_r4_c50_9 + t_r4_c50_10;
  assign t_r4_c50_12 = t_r4_c50_11 + p_5_51;
  assign out_4_50 = t_r4_c50_12 >> 4;

  assign t_r4_c51_0 = p_3_51 << 1;
  assign t_r4_c51_1 = p_4_50 << 1;
  assign t_r4_c51_2 = p_4_51 << 2;
  assign t_r4_c51_3 = p_4_52 << 1;
  assign t_r4_c51_4 = p_5_51 << 1;
  assign t_r4_c51_5 = t_r4_c51_0 + p_3_50;
  assign t_r4_c51_6 = t_r4_c51_1 + p_3_52;
  assign t_r4_c51_7 = t_r4_c51_2 + t_r4_c51_3;
  assign t_r4_c51_8 = t_r4_c51_4 + p_5_50;
  assign t_r4_c51_9 = t_r4_c51_5 + t_r4_c51_6;
  assign t_r4_c51_10 = t_r4_c51_7 + t_r4_c51_8;
  assign t_r4_c51_11 = t_r4_c51_9 + t_r4_c51_10;
  assign t_r4_c51_12 = t_r4_c51_11 + p_5_52;
  assign out_4_51 = t_r4_c51_12 >> 4;

  assign t_r4_c52_0 = p_3_52 << 1;
  assign t_r4_c52_1 = p_4_51 << 1;
  assign t_r4_c52_2 = p_4_52 << 2;
  assign t_r4_c52_3 = p_4_53 << 1;
  assign t_r4_c52_4 = p_5_52 << 1;
  assign t_r4_c52_5 = t_r4_c52_0 + p_3_51;
  assign t_r4_c52_6 = t_r4_c52_1 + p_3_53;
  assign t_r4_c52_7 = t_r4_c52_2 + t_r4_c52_3;
  assign t_r4_c52_8 = t_r4_c52_4 + p_5_51;
  assign t_r4_c52_9 = t_r4_c52_5 + t_r4_c52_6;
  assign t_r4_c52_10 = t_r4_c52_7 + t_r4_c52_8;
  assign t_r4_c52_11 = t_r4_c52_9 + t_r4_c52_10;
  assign t_r4_c52_12 = t_r4_c52_11 + p_5_53;
  assign out_4_52 = t_r4_c52_12 >> 4;

  assign t_r4_c53_0 = p_3_53 << 1;
  assign t_r4_c53_1 = p_4_52 << 1;
  assign t_r4_c53_2 = p_4_53 << 2;
  assign t_r4_c53_3 = p_4_54 << 1;
  assign t_r4_c53_4 = p_5_53 << 1;
  assign t_r4_c53_5 = t_r4_c53_0 + p_3_52;
  assign t_r4_c53_6 = t_r4_c53_1 + p_3_54;
  assign t_r4_c53_7 = t_r4_c53_2 + t_r4_c53_3;
  assign t_r4_c53_8 = t_r4_c53_4 + p_5_52;
  assign t_r4_c53_9 = t_r4_c53_5 + t_r4_c53_6;
  assign t_r4_c53_10 = t_r4_c53_7 + t_r4_c53_8;
  assign t_r4_c53_11 = t_r4_c53_9 + t_r4_c53_10;
  assign t_r4_c53_12 = t_r4_c53_11 + p_5_54;
  assign out_4_53 = t_r4_c53_12 >> 4;

  assign t_r4_c54_0 = p_3_54 << 1;
  assign t_r4_c54_1 = p_4_53 << 1;
  assign t_r4_c54_2 = p_4_54 << 2;
  assign t_r4_c54_3 = p_4_55 << 1;
  assign t_r4_c54_4 = p_5_54 << 1;
  assign t_r4_c54_5 = t_r4_c54_0 + p_3_53;
  assign t_r4_c54_6 = t_r4_c54_1 + p_3_55;
  assign t_r4_c54_7 = t_r4_c54_2 + t_r4_c54_3;
  assign t_r4_c54_8 = t_r4_c54_4 + p_5_53;
  assign t_r4_c54_9 = t_r4_c54_5 + t_r4_c54_6;
  assign t_r4_c54_10 = t_r4_c54_7 + t_r4_c54_8;
  assign t_r4_c54_11 = t_r4_c54_9 + t_r4_c54_10;
  assign t_r4_c54_12 = t_r4_c54_11 + p_5_55;
  assign out_4_54 = t_r4_c54_12 >> 4;

  assign t_r4_c55_0 = p_3_55 << 1;
  assign t_r4_c55_1 = p_4_54 << 1;
  assign t_r4_c55_2 = p_4_55 << 2;
  assign t_r4_c55_3 = p_4_56 << 1;
  assign t_r4_c55_4 = p_5_55 << 1;
  assign t_r4_c55_5 = t_r4_c55_0 + p_3_54;
  assign t_r4_c55_6 = t_r4_c55_1 + p_3_56;
  assign t_r4_c55_7 = t_r4_c55_2 + t_r4_c55_3;
  assign t_r4_c55_8 = t_r4_c55_4 + p_5_54;
  assign t_r4_c55_9 = t_r4_c55_5 + t_r4_c55_6;
  assign t_r4_c55_10 = t_r4_c55_7 + t_r4_c55_8;
  assign t_r4_c55_11 = t_r4_c55_9 + t_r4_c55_10;
  assign t_r4_c55_12 = t_r4_c55_11 + p_5_56;
  assign out_4_55 = t_r4_c55_12 >> 4;

  assign t_r4_c56_0 = p_3_56 << 1;
  assign t_r4_c56_1 = p_4_55 << 1;
  assign t_r4_c56_2 = p_4_56 << 2;
  assign t_r4_c56_3 = p_4_57 << 1;
  assign t_r4_c56_4 = p_5_56 << 1;
  assign t_r4_c56_5 = t_r4_c56_0 + p_3_55;
  assign t_r4_c56_6 = t_r4_c56_1 + p_3_57;
  assign t_r4_c56_7 = t_r4_c56_2 + t_r4_c56_3;
  assign t_r4_c56_8 = t_r4_c56_4 + p_5_55;
  assign t_r4_c56_9 = t_r4_c56_5 + t_r4_c56_6;
  assign t_r4_c56_10 = t_r4_c56_7 + t_r4_c56_8;
  assign t_r4_c56_11 = t_r4_c56_9 + t_r4_c56_10;
  assign t_r4_c56_12 = t_r4_c56_11 + p_5_57;
  assign out_4_56 = t_r4_c56_12 >> 4;

  assign t_r4_c57_0 = p_3_57 << 1;
  assign t_r4_c57_1 = p_4_56 << 1;
  assign t_r4_c57_2 = p_4_57 << 2;
  assign t_r4_c57_3 = p_4_58 << 1;
  assign t_r4_c57_4 = p_5_57 << 1;
  assign t_r4_c57_5 = t_r4_c57_0 + p_3_56;
  assign t_r4_c57_6 = t_r4_c57_1 + p_3_58;
  assign t_r4_c57_7 = t_r4_c57_2 + t_r4_c57_3;
  assign t_r4_c57_8 = t_r4_c57_4 + p_5_56;
  assign t_r4_c57_9 = t_r4_c57_5 + t_r4_c57_6;
  assign t_r4_c57_10 = t_r4_c57_7 + t_r4_c57_8;
  assign t_r4_c57_11 = t_r4_c57_9 + t_r4_c57_10;
  assign t_r4_c57_12 = t_r4_c57_11 + p_5_58;
  assign out_4_57 = t_r4_c57_12 >> 4;

  assign t_r4_c58_0 = p_3_58 << 1;
  assign t_r4_c58_1 = p_4_57 << 1;
  assign t_r4_c58_2 = p_4_58 << 2;
  assign t_r4_c58_3 = p_4_59 << 1;
  assign t_r4_c58_4 = p_5_58 << 1;
  assign t_r4_c58_5 = t_r4_c58_0 + p_3_57;
  assign t_r4_c58_6 = t_r4_c58_1 + p_3_59;
  assign t_r4_c58_7 = t_r4_c58_2 + t_r4_c58_3;
  assign t_r4_c58_8 = t_r4_c58_4 + p_5_57;
  assign t_r4_c58_9 = t_r4_c58_5 + t_r4_c58_6;
  assign t_r4_c58_10 = t_r4_c58_7 + t_r4_c58_8;
  assign t_r4_c58_11 = t_r4_c58_9 + t_r4_c58_10;
  assign t_r4_c58_12 = t_r4_c58_11 + p_5_59;
  assign out_4_58 = t_r4_c58_12 >> 4;

  assign t_r4_c59_0 = p_3_59 << 1;
  assign t_r4_c59_1 = p_4_58 << 1;
  assign t_r4_c59_2 = p_4_59 << 2;
  assign t_r4_c59_3 = p_4_60 << 1;
  assign t_r4_c59_4 = p_5_59 << 1;
  assign t_r4_c59_5 = t_r4_c59_0 + p_3_58;
  assign t_r4_c59_6 = t_r4_c59_1 + p_3_60;
  assign t_r4_c59_7 = t_r4_c59_2 + t_r4_c59_3;
  assign t_r4_c59_8 = t_r4_c59_4 + p_5_58;
  assign t_r4_c59_9 = t_r4_c59_5 + t_r4_c59_6;
  assign t_r4_c59_10 = t_r4_c59_7 + t_r4_c59_8;
  assign t_r4_c59_11 = t_r4_c59_9 + t_r4_c59_10;
  assign t_r4_c59_12 = t_r4_c59_11 + p_5_60;
  assign out_4_59 = t_r4_c59_12 >> 4;

  assign t_r4_c60_0 = p_3_60 << 1;
  assign t_r4_c60_1 = p_4_59 << 1;
  assign t_r4_c60_2 = p_4_60 << 2;
  assign t_r4_c60_3 = p_4_61 << 1;
  assign t_r4_c60_4 = p_5_60 << 1;
  assign t_r4_c60_5 = t_r4_c60_0 + p_3_59;
  assign t_r4_c60_6 = t_r4_c60_1 + p_3_61;
  assign t_r4_c60_7 = t_r4_c60_2 + t_r4_c60_3;
  assign t_r4_c60_8 = t_r4_c60_4 + p_5_59;
  assign t_r4_c60_9 = t_r4_c60_5 + t_r4_c60_6;
  assign t_r4_c60_10 = t_r4_c60_7 + t_r4_c60_8;
  assign t_r4_c60_11 = t_r4_c60_9 + t_r4_c60_10;
  assign t_r4_c60_12 = t_r4_c60_11 + p_5_61;
  assign out_4_60 = t_r4_c60_12 >> 4;

  assign t_r4_c61_0 = p_3_61 << 1;
  assign t_r4_c61_1 = p_4_60 << 1;
  assign t_r4_c61_2 = p_4_61 << 2;
  assign t_r4_c61_3 = p_4_62 << 1;
  assign t_r4_c61_4 = p_5_61 << 1;
  assign t_r4_c61_5 = t_r4_c61_0 + p_3_60;
  assign t_r4_c61_6 = t_r4_c61_1 + p_3_62;
  assign t_r4_c61_7 = t_r4_c61_2 + t_r4_c61_3;
  assign t_r4_c61_8 = t_r4_c61_4 + p_5_60;
  assign t_r4_c61_9 = t_r4_c61_5 + t_r4_c61_6;
  assign t_r4_c61_10 = t_r4_c61_7 + t_r4_c61_8;
  assign t_r4_c61_11 = t_r4_c61_9 + t_r4_c61_10;
  assign t_r4_c61_12 = t_r4_c61_11 + p_5_62;
  assign out_4_61 = t_r4_c61_12 >> 4;

  assign t_r4_c62_0 = p_3_62 << 1;
  assign t_r4_c62_1 = p_4_61 << 1;
  assign t_r4_c62_2 = p_4_62 << 2;
  assign t_r4_c62_3 = p_4_63 << 1;
  assign t_r4_c62_4 = p_5_62 << 1;
  assign t_r4_c62_5 = t_r4_c62_0 + p_3_61;
  assign t_r4_c62_6 = t_r4_c62_1 + p_3_63;
  assign t_r4_c62_7 = t_r4_c62_2 + t_r4_c62_3;
  assign t_r4_c62_8 = t_r4_c62_4 + p_5_61;
  assign t_r4_c62_9 = t_r4_c62_5 + t_r4_c62_6;
  assign t_r4_c62_10 = t_r4_c62_7 + t_r4_c62_8;
  assign t_r4_c62_11 = t_r4_c62_9 + t_r4_c62_10;
  assign t_r4_c62_12 = t_r4_c62_11 + p_5_63;
  assign out_4_62 = t_r4_c62_12 >> 4;

  assign t_r4_c63_0 = p_3_63 << 1;
  assign t_r4_c63_1 = p_4_62 << 1;
  assign t_r4_c63_2 = p_4_63 << 2;
  assign t_r4_c63_3 = p_4_64 << 1;
  assign t_r4_c63_4 = p_5_63 << 1;
  assign t_r4_c63_5 = t_r4_c63_0 + p_3_62;
  assign t_r4_c63_6 = t_r4_c63_1 + p_3_64;
  assign t_r4_c63_7 = t_r4_c63_2 + t_r4_c63_3;
  assign t_r4_c63_8 = t_r4_c63_4 + p_5_62;
  assign t_r4_c63_9 = t_r4_c63_5 + t_r4_c63_6;
  assign t_r4_c63_10 = t_r4_c63_7 + t_r4_c63_8;
  assign t_r4_c63_11 = t_r4_c63_9 + t_r4_c63_10;
  assign t_r4_c63_12 = t_r4_c63_11 + p_5_64;
  assign out_4_63 = t_r4_c63_12 >> 4;

  assign t_r4_c64_0 = p_3_64 << 1;
  assign t_r4_c64_1 = p_4_63 << 1;
  assign t_r4_c64_2 = p_4_64 << 2;
  assign t_r4_c64_3 = p_4_65 << 1;
  assign t_r4_c64_4 = p_5_64 << 1;
  assign t_r4_c64_5 = t_r4_c64_0 + p_3_63;
  assign t_r4_c64_6 = t_r4_c64_1 + p_3_65;
  assign t_r4_c64_7 = t_r4_c64_2 + t_r4_c64_3;
  assign t_r4_c64_8 = t_r4_c64_4 + p_5_63;
  assign t_r4_c64_9 = t_r4_c64_5 + t_r4_c64_6;
  assign t_r4_c64_10 = t_r4_c64_7 + t_r4_c64_8;
  assign t_r4_c64_11 = t_r4_c64_9 + t_r4_c64_10;
  assign t_r4_c64_12 = t_r4_c64_11 + p_5_65;
  assign out_4_64 = t_r4_c64_12 >> 4;

  assign t_r5_c1_0 = p_4_1 << 1;
  assign t_r5_c1_1 = p_5_0 << 1;
  assign t_r5_c1_2 = p_5_1 << 2;
  assign t_r5_c1_3 = p_5_2 << 1;
  assign t_r5_c1_4 = p_6_1 << 1;
  assign t_r5_c1_5 = t_r5_c1_0 + p_4_0;
  assign t_r5_c1_6 = t_r5_c1_1 + p_4_2;
  assign t_r5_c1_7 = t_r5_c1_2 + t_r5_c1_3;
  assign t_r5_c1_8 = t_r5_c1_4 + p_6_0;
  assign t_r5_c1_9 = t_r5_c1_5 + t_r5_c1_6;
  assign t_r5_c1_10 = t_r5_c1_7 + t_r5_c1_8;
  assign t_r5_c1_11 = t_r5_c1_9 + t_r5_c1_10;
  assign t_r5_c1_12 = t_r5_c1_11 + p_6_2;
  assign out_5_1 = t_r5_c1_12 >> 4;

  assign t_r5_c2_0 = p_4_2 << 1;
  assign t_r5_c2_1 = p_5_1 << 1;
  assign t_r5_c2_2 = p_5_2 << 2;
  assign t_r5_c2_3 = p_5_3 << 1;
  assign t_r5_c2_4 = p_6_2 << 1;
  assign t_r5_c2_5 = t_r5_c2_0 + p_4_1;
  assign t_r5_c2_6 = t_r5_c2_1 + p_4_3;
  assign t_r5_c2_7 = t_r5_c2_2 + t_r5_c2_3;
  assign t_r5_c2_8 = t_r5_c2_4 + p_6_1;
  assign t_r5_c2_9 = t_r5_c2_5 + t_r5_c2_6;
  assign t_r5_c2_10 = t_r5_c2_7 + t_r5_c2_8;
  assign t_r5_c2_11 = t_r5_c2_9 + t_r5_c2_10;
  assign t_r5_c2_12 = t_r5_c2_11 + p_6_3;
  assign out_5_2 = t_r5_c2_12 >> 4;

  assign t_r5_c3_0 = p_4_3 << 1;
  assign t_r5_c3_1 = p_5_2 << 1;
  assign t_r5_c3_2 = p_5_3 << 2;
  assign t_r5_c3_3 = p_5_4 << 1;
  assign t_r5_c3_4 = p_6_3 << 1;
  assign t_r5_c3_5 = t_r5_c3_0 + p_4_2;
  assign t_r5_c3_6 = t_r5_c3_1 + p_4_4;
  assign t_r5_c3_7 = t_r5_c3_2 + t_r5_c3_3;
  assign t_r5_c3_8 = t_r5_c3_4 + p_6_2;
  assign t_r5_c3_9 = t_r5_c3_5 + t_r5_c3_6;
  assign t_r5_c3_10 = t_r5_c3_7 + t_r5_c3_8;
  assign t_r5_c3_11 = t_r5_c3_9 + t_r5_c3_10;
  assign t_r5_c3_12 = t_r5_c3_11 + p_6_4;
  assign out_5_3 = t_r5_c3_12 >> 4;

  assign t_r5_c4_0 = p_4_4 << 1;
  assign t_r5_c4_1 = p_5_3 << 1;
  assign t_r5_c4_2 = p_5_4 << 2;
  assign t_r5_c4_3 = p_5_5 << 1;
  assign t_r5_c4_4 = p_6_4 << 1;
  assign t_r5_c4_5 = t_r5_c4_0 + p_4_3;
  assign t_r5_c4_6 = t_r5_c4_1 + p_4_5;
  assign t_r5_c4_7 = t_r5_c4_2 + t_r5_c4_3;
  assign t_r5_c4_8 = t_r5_c4_4 + p_6_3;
  assign t_r5_c4_9 = t_r5_c4_5 + t_r5_c4_6;
  assign t_r5_c4_10 = t_r5_c4_7 + t_r5_c4_8;
  assign t_r5_c4_11 = t_r5_c4_9 + t_r5_c4_10;
  assign t_r5_c4_12 = t_r5_c4_11 + p_6_5;
  assign out_5_4 = t_r5_c4_12 >> 4;

  assign t_r5_c5_0 = p_4_5 << 1;
  assign t_r5_c5_1 = p_5_4 << 1;
  assign t_r5_c5_2 = p_5_5 << 2;
  assign t_r5_c5_3 = p_5_6 << 1;
  assign t_r5_c5_4 = p_6_5 << 1;
  assign t_r5_c5_5 = t_r5_c5_0 + p_4_4;
  assign t_r5_c5_6 = t_r5_c5_1 + p_4_6;
  assign t_r5_c5_7 = t_r5_c5_2 + t_r5_c5_3;
  assign t_r5_c5_8 = t_r5_c5_4 + p_6_4;
  assign t_r5_c5_9 = t_r5_c5_5 + t_r5_c5_6;
  assign t_r5_c5_10 = t_r5_c5_7 + t_r5_c5_8;
  assign t_r5_c5_11 = t_r5_c5_9 + t_r5_c5_10;
  assign t_r5_c5_12 = t_r5_c5_11 + p_6_6;
  assign out_5_5 = t_r5_c5_12 >> 4;

  assign t_r5_c6_0 = p_4_6 << 1;
  assign t_r5_c6_1 = p_5_5 << 1;
  assign t_r5_c6_2 = p_5_6 << 2;
  assign t_r5_c6_3 = p_5_7 << 1;
  assign t_r5_c6_4 = p_6_6 << 1;
  assign t_r5_c6_5 = t_r5_c6_0 + p_4_5;
  assign t_r5_c6_6 = t_r5_c6_1 + p_4_7;
  assign t_r5_c6_7 = t_r5_c6_2 + t_r5_c6_3;
  assign t_r5_c6_8 = t_r5_c6_4 + p_6_5;
  assign t_r5_c6_9 = t_r5_c6_5 + t_r5_c6_6;
  assign t_r5_c6_10 = t_r5_c6_7 + t_r5_c6_8;
  assign t_r5_c6_11 = t_r5_c6_9 + t_r5_c6_10;
  assign t_r5_c6_12 = t_r5_c6_11 + p_6_7;
  assign out_5_6 = t_r5_c6_12 >> 4;

  assign t_r5_c7_0 = p_4_7 << 1;
  assign t_r5_c7_1 = p_5_6 << 1;
  assign t_r5_c7_2 = p_5_7 << 2;
  assign t_r5_c7_3 = p_5_8 << 1;
  assign t_r5_c7_4 = p_6_7 << 1;
  assign t_r5_c7_5 = t_r5_c7_0 + p_4_6;
  assign t_r5_c7_6 = t_r5_c7_1 + p_4_8;
  assign t_r5_c7_7 = t_r5_c7_2 + t_r5_c7_3;
  assign t_r5_c7_8 = t_r5_c7_4 + p_6_6;
  assign t_r5_c7_9 = t_r5_c7_5 + t_r5_c7_6;
  assign t_r5_c7_10 = t_r5_c7_7 + t_r5_c7_8;
  assign t_r5_c7_11 = t_r5_c7_9 + t_r5_c7_10;
  assign t_r5_c7_12 = t_r5_c7_11 + p_6_8;
  assign out_5_7 = t_r5_c7_12 >> 4;

  assign t_r5_c8_0 = p_4_8 << 1;
  assign t_r5_c8_1 = p_5_7 << 1;
  assign t_r5_c8_2 = p_5_8 << 2;
  assign t_r5_c8_3 = p_5_9 << 1;
  assign t_r5_c8_4 = p_6_8 << 1;
  assign t_r5_c8_5 = t_r5_c8_0 + p_4_7;
  assign t_r5_c8_6 = t_r5_c8_1 + p_4_9;
  assign t_r5_c8_7 = t_r5_c8_2 + t_r5_c8_3;
  assign t_r5_c8_8 = t_r5_c8_4 + p_6_7;
  assign t_r5_c8_9 = t_r5_c8_5 + t_r5_c8_6;
  assign t_r5_c8_10 = t_r5_c8_7 + t_r5_c8_8;
  assign t_r5_c8_11 = t_r5_c8_9 + t_r5_c8_10;
  assign t_r5_c8_12 = t_r5_c8_11 + p_6_9;
  assign out_5_8 = t_r5_c8_12 >> 4;

  assign t_r5_c9_0 = p_4_9 << 1;
  assign t_r5_c9_1 = p_5_8 << 1;
  assign t_r5_c9_2 = p_5_9 << 2;
  assign t_r5_c9_3 = p_5_10 << 1;
  assign t_r5_c9_4 = p_6_9 << 1;
  assign t_r5_c9_5 = t_r5_c9_0 + p_4_8;
  assign t_r5_c9_6 = t_r5_c9_1 + p_4_10;
  assign t_r5_c9_7 = t_r5_c9_2 + t_r5_c9_3;
  assign t_r5_c9_8 = t_r5_c9_4 + p_6_8;
  assign t_r5_c9_9 = t_r5_c9_5 + t_r5_c9_6;
  assign t_r5_c9_10 = t_r5_c9_7 + t_r5_c9_8;
  assign t_r5_c9_11 = t_r5_c9_9 + t_r5_c9_10;
  assign t_r5_c9_12 = t_r5_c9_11 + p_6_10;
  assign out_5_9 = t_r5_c9_12 >> 4;

  assign t_r5_c10_0 = p_4_10 << 1;
  assign t_r5_c10_1 = p_5_9 << 1;
  assign t_r5_c10_2 = p_5_10 << 2;
  assign t_r5_c10_3 = p_5_11 << 1;
  assign t_r5_c10_4 = p_6_10 << 1;
  assign t_r5_c10_5 = t_r5_c10_0 + p_4_9;
  assign t_r5_c10_6 = t_r5_c10_1 + p_4_11;
  assign t_r5_c10_7 = t_r5_c10_2 + t_r5_c10_3;
  assign t_r5_c10_8 = t_r5_c10_4 + p_6_9;
  assign t_r5_c10_9 = t_r5_c10_5 + t_r5_c10_6;
  assign t_r5_c10_10 = t_r5_c10_7 + t_r5_c10_8;
  assign t_r5_c10_11 = t_r5_c10_9 + t_r5_c10_10;
  assign t_r5_c10_12 = t_r5_c10_11 + p_6_11;
  assign out_5_10 = t_r5_c10_12 >> 4;

  assign t_r5_c11_0 = p_4_11 << 1;
  assign t_r5_c11_1 = p_5_10 << 1;
  assign t_r5_c11_2 = p_5_11 << 2;
  assign t_r5_c11_3 = p_5_12 << 1;
  assign t_r5_c11_4 = p_6_11 << 1;
  assign t_r5_c11_5 = t_r5_c11_0 + p_4_10;
  assign t_r5_c11_6 = t_r5_c11_1 + p_4_12;
  assign t_r5_c11_7 = t_r5_c11_2 + t_r5_c11_3;
  assign t_r5_c11_8 = t_r5_c11_4 + p_6_10;
  assign t_r5_c11_9 = t_r5_c11_5 + t_r5_c11_6;
  assign t_r5_c11_10 = t_r5_c11_7 + t_r5_c11_8;
  assign t_r5_c11_11 = t_r5_c11_9 + t_r5_c11_10;
  assign t_r5_c11_12 = t_r5_c11_11 + p_6_12;
  assign out_5_11 = t_r5_c11_12 >> 4;

  assign t_r5_c12_0 = p_4_12 << 1;
  assign t_r5_c12_1 = p_5_11 << 1;
  assign t_r5_c12_2 = p_5_12 << 2;
  assign t_r5_c12_3 = p_5_13 << 1;
  assign t_r5_c12_4 = p_6_12 << 1;
  assign t_r5_c12_5 = t_r5_c12_0 + p_4_11;
  assign t_r5_c12_6 = t_r5_c12_1 + p_4_13;
  assign t_r5_c12_7 = t_r5_c12_2 + t_r5_c12_3;
  assign t_r5_c12_8 = t_r5_c12_4 + p_6_11;
  assign t_r5_c12_9 = t_r5_c12_5 + t_r5_c12_6;
  assign t_r5_c12_10 = t_r5_c12_7 + t_r5_c12_8;
  assign t_r5_c12_11 = t_r5_c12_9 + t_r5_c12_10;
  assign t_r5_c12_12 = t_r5_c12_11 + p_6_13;
  assign out_5_12 = t_r5_c12_12 >> 4;

  assign t_r5_c13_0 = p_4_13 << 1;
  assign t_r5_c13_1 = p_5_12 << 1;
  assign t_r5_c13_2 = p_5_13 << 2;
  assign t_r5_c13_3 = p_5_14 << 1;
  assign t_r5_c13_4 = p_6_13 << 1;
  assign t_r5_c13_5 = t_r5_c13_0 + p_4_12;
  assign t_r5_c13_6 = t_r5_c13_1 + p_4_14;
  assign t_r5_c13_7 = t_r5_c13_2 + t_r5_c13_3;
  assign t_r5_c13_8 = t_r5_c13_4 + p_6_12;
  assign t_r5_c13_9 = t_r5_c13_5 + t_r5_c13_6;
  assign t_r5_c13_10 = t_r5_c13_7 + t_r5_c13_8;
  assign t_r5_c13_11 = t_r5_c13_9 + t_r5_c13_10;
  assign t_r5_c13_12 = t_r5_c13_11 + p_6_14;
  assign out_5_13 = t_r5_c13_12 >> 4;

  assign t_r5_c14_0 = p_4_14 << 1;
  assign t_r5_c14_1 = p_5_13 << 1;
  assign t_r5_c14_2 = p_5_14 << 2;
  assign t_r5_c14_3 = p_5_15 << 1;
  assign t_r5_c14_4 = p_6_14 << 1;
  assign t_r5_c14_5 = t_r5_c14_0 + p_4_13;
  assign t_r5_c14_6 = t_r5_c14_1 + p_4_15;
  assign t_r5_c14_7 = t_r5_c14_2 + t_r5_c14_3;
  assign t_r5_c14_8 = t_r5_c14_4 + p_6_13;
  assign t_r5_c14_9 = t_r5_c14_5 + t_r5_c14_6;
  assign t_r5_c14_10 = t_r5_c14_7 + t_r5_c14_8;
  assign t_r5_c14_11 = t_r5_c14_9 + t_r5_c14_10;
  assign t_r5_c14_12 = t_r5_c14_11 + p_6_15;
  assign out_5_14 = t_r5_c14_12 >> 4;

  assign t_r5_c15_0 = p_4_15 << 1;
  assign t_r5_c15_1 = p_5_14 << 1;
  assign t_r5_c15_2 = p_5_15 << 2;
  assign t_r5_c15_3 = p_5_16 << 1;
  assign t_r5_c15_4 = p_6_15 << 1;
  assign t_r5_c15_5 = t_r5_c15_0 + p_4_14;
  assign t_r5_c15_6 = t_r5_c15_1 + p_4_16;
  assign t_r5_c15_7 = t_r5_c15_2 + t_r5_c15_3;
  assign t_r5_c15_8 = t_r5_c15_4 + p_6_14;
  assign t_r5_c15_9 = t_r5_c15_5 + t_r5_c15_6;
  assign t_r5_c15_10 = t_r5_c15_7 + t_r5_c15_8;
  assign t_r5_c15_11 = t_r5_c15_9 + t_r5_c15_10;
  assign t_r5_c15_12 = t_r5_c15_11 + p_6_16;
  assign out_5_15 = t_r5_c15_12 >> 4;

  assign t_r5_c16_0 = p_4_16 << 1;
  assign t_r5_c16_1 = p_5_15 << 1;
  assign t_r5_c16_2 = p_5_16 << 2;
  assign t_r5_c16_3 = p_5_17 << 1;
  assign t_r5_c16_4 = p_6_16 << 1;
  assign t_r5_c16_5 = t_r5_c16_0 + p_4_15;
  assign t_r5_c16_6 = t_r5_c16_1 + p_4_17;
  assign t_r5_c16_7 = t_r5_c16_2 + t_r5_c16_3;
  assign t_r5_c16_8 = t_r5_c16_4 + p_6_15;
  assign t_r5_c16_9 = t_r5_c16_5 + t_r5_c16_6;
  assign t_r5_c16_10 = t_r5_c16_7 + t_r5_c16_8;
  assign t_r5_c16_11 = t_r5_c16_9 + t_r5_c16_10;
  assign t_r5_c16_12 = t_r5_c16_11 + p_6_17;
  assign out_5_16 = t_r5_c16_12 >> 4;

  assign t_r5_c17_0 = p_4_17 << 1;
  assign t_r5_c17_1 = p_5_16 << 1;
  assign t_r5_c17_2 = p_5_17 << 2;
  assign t_r5_c17_3 = p_5_18 << 1;
  assign t_r5_c17_4 = p_6_17 << 1;
  assign t_r5_c17_5 = t_r5_c17_0 + p_4_16;
  assign t_r5_c17_6 = t_r5_c17_1 + p_4_18;
  assign t_r5_c17_7 = t_r5_c17_2 + t_r5_c17_3;
  assign t_r5_c17_8 = t_r5_c17_4 + p_6_16;
  assign t_r5_c17_9 = t_r5_c17_5 + t_r5_c17_6;
  assign t_r5_c17_10 = t_r5_c17_7 + t_r5_c17_8;
  assign t_r5_c17_11 = t_r5_c17_9 + t_r5_c17_10;
  assign t_r5_c17_12 = t_r5_c17_11 + p_6_18;
  assign out_5_17 = t_r5_c17_12 >> 4;

  assign t_r5_c18_0 = p_4_18 << 1;
  assign t_r5_c18_1 = p_5_17 << 1;
  assign t_r5_c18_2 = p_5_18 << 2;
  assign t_r5_c18_3 = p_5_19 << 1;
  assign t_r5_c18_4 = p_6_18 << 1;
  assign t_r5_c18_5 = t_r5_c18_0 + p_4_17;
  assign t_r5_c18_6 = t_r5_c18_1 + p_4_19;
  assign t_r5_c18_7 = t_r5_c18_2 + t_r5_c18_3;
  assign t_r5_c18_8 = t_r5_c18_4 + p_6_17;
  assign t_r5_c18_9 = t_r5_c18_5 + t_r5_c18_6;
  assign t_r5_c18_10 = t_r5_c18_7 + t_r5_c18_8;
  assign t_r5_c18_11 = t_r5_c18_9 + t_r5_c18_10;
  assign t_r5_c18_12 = t_r5_c18_11 + p_6_19;
  assign out_5_18 = t_r5_c18_12 >> 4;

  assign t_r5_c19_0 = p_4_19 << 1;
  assign t_r5_c19_1 = p_5_18 << 1;
  assign t_r5_c19_2 = p_5_19 << 2;
  assign t_r5_c19_3 = p_5_20 << 1;
  assign t_r5_c19_4 = p_6_19 << 1;
  assign t_r5_c19_5 = t_r5_c19_0 + p_4_18;
  assign t_r5_c19_6 = t_r5_c19_1 + p_4_20;
  assign t_r5_c19_7 = t_r5_c19_2 + t_r5_c19_3;
  assign t_r5_c19_8 = t_r5_c19_4 + p_6_18;
  assign t_r5_c19_9 = t_r5_c19_5 + t_r5_c19_6;
  assign t_r5_c19_10 = t_r5_c19_7 + t_r5_c19_8;
  assign t_r5_c19_11 = t_r5_c19_9 + t_r5_c19_10;
  assign t_r5_c19_12 = t_r5_c19_11 + p_6_20;
  assign out_5_19 = t_r5_c19_12 >> 4;

  assign t_r5_c20_0 = p_4_20 << 1;
  assign t_r5_c20_1 = p_5_19 << 1;
  assign t_r5_c20_2 = p_5_20 << 2;
  assign t_r5_c20_3 = p_5_21 << 1;
  assign t_r5_c20_4 = p_6_20 << 1;
  assign t_r5_c20_5 = t_r5_c20_0 + p_4_19;
  assign t_r5_c20_6 = t_r5_c20_1 + p_4_21;
  assign t_r5_c20_7 = t_r5_c20_2 + t_r5_c20_3;
  assign t_r5_c20_8 = t_r5_c20_4 + p_6_19;
  assign t_r5_c20_9 = t_r5_c20_5 + t_r5_c20_6;
  assign t_r5_c20_10 = t_r5_c20_7 + t_r5_c20_8;
  assign t_r5_c20_11 = t_r5_c20_9 + t_r5_c20_10;
  assign t_r5_c20_12 = t_r5_c20_11 + p_6_21;
  assign out_5_20 = t_r5_c20_12 >> 4;

  assign t_r5_c21_0 = p_4_21 << 1;
  assign t_r5_c21_1 = p_5_20 << 1;
  assign t_r5_c21_2 = p_5_21 << 2;
  assign t_r5_c21_3 = p_5_22 << 1;
  assign t_r5_c21_4 = p_6_21 << 1;
  assign t_r5_c21_5 = t_r5_c21_0 + p_4_20;
  assign t_r5_c21_6 = t_r5_c21_1 + p_4_22;
  assign t_r5_c21_7 = t_r5_c21_2 + t_r5_c21_3;
  assign t_r5_c21_8 = t_r5_c21_4 + p_6_20;
  assign t_r5_c21_9 = t_r5_c21_5 + t_r5_c21_6;
  assign t_r5_c21_10 = t_r5_c21_7 + t_r5_c21_8;
  assign t_r5_c21_11 = t_r5_c21_9 + t_r5_c21_10;
  assign t_r5_c21_12 = t_r5_c21_11 + p_6_22;
  assign out_5_21 = t_r5_c21_12 >> 4;

  assign t_r5_c22_0 = p_4_22 << 1;
  assign t_r5_c22_1 = p_5_21 << 1;
  assign t_r5_c22_2 = p_5_22 << 2;
  assign t_r5_c22_3 = p_5_23 << 1;
  assign t_r5_c22_4 = p_6_22 << 1;
  assign t_r5_c22_5 = t_r5_c22_0 + p_4_21;
  assign t_r5_c22_6 = t_r5_c22_1 + p_4_23;
  assign t_r5_c22_7 = t_r5_c22_2 + t_r5_c22_3;
  assign t_r5_c22_8 = t_r5_c22_4 + p_6_21;
  assign t_r5_c22_9 = t_r5_c22_5 + t_r5_c22_6;
  assign t_r5_c22_10 = t_r5_c22_7 + t_r5_c22_8;
  assign t_r5_c22_11 = t_r5_c22_9 + t_r5_c22_10;
  assign t_r5_c22_12 = t_r5_c22_11 + p_6_23;
  assign out_5_22 = t_r5_c22_12 >> 4;

  assign t_r5_c23_0 = p_4_23 << 1;
  assign t_r5_c23_1 = p_5_22 << 1;
  assign t_r5_c23_2 = p_5_23 << 2;
  assign t_r5_c23_3 = p_5_24 << 1;
  assign t_r5_c23_4 = p_6_23 << 1;
  assign t_r5_c23_5 = t_r5_c23_0 + p_4_22;
  assign t_r5_c23_6 = t_r5_c23_1 + p_4_24;
  assign t_r5_c23_7 = t_r5_c23_2 + t_r5_c23_3;
  assign t_r5_c23_8 = t_r5_c23_4 + p_6_22;
  assign t_r5_c23_9 = t_r5_c23_5 + t_r5_c23_6;
  assign t_r5_c23_10 = t_r5_c23_7 + t_r5_c23_8;
  assign t_r5_c23_11 = t_r5_c23_9 + t_r5_c23_10;
  assign t_r5_c23_12 = t_r5_c23_11 + p_6_24;
  assign out_5_23 = t_r5_c23_12 >> 4;

  assign t_r5_c24_0 = p_4_24 << 1;
  assign t_r5_c24_1 = p_5_23 << 1;
  assign t_r5_c24_2 = p_5_24 << 2;
  assign t_r5_c24_3 = p_5_25 << 1;
  assign t_r5_c24_4 = p_6_24 << 1;
  assign t_r5_c24_5 = t_r5_c24_0 + p_4_23;
  assign t_r5_c24_6 = t_r5_c24_1 + p_4_25;
  assign t_r5_c24_7 = t_r5_c24_2 + t_r5_c24_3;
  assign t_r5_c24_8 = t_r5_c24_4 + p_6_23;
  assign t_r5_c24_9 = t_r5_c24_5 + t_r5_c24_6;
  assign t_r5_c24_10 = t_r5_c24_7 + t_r5_c24_8;
  assign t_r5_c24_11 = t_r5_c24_9 + t_r5_c24_10;
  assign t_r5_c24_12 = t_r5_c24_11 + p_6_25;
  assign out_5_24 = t_r5_c24_12 >> 4;

  assign t_r5_c25_0 = p_4_25 << 1;
  assign t_r5_c25_1 = p_5_24 << 1;
  assign t_r5_c25_2 = p_5_25 << 2;
  assign t_r5_c25_3 = p_5_26 << 1;
  assign t_r5_c25_4 = p_6_25 << 1;
  assign t_r5_c25_5 = t_r5_c25_0 + p_4_24;
  assign t_r5_c25_6 = t_r5_c25_1 + p_4_26;
  assign t_r5_c25_7 = t_r5_c25_2 + t_r5_c25_3;
  assign t_r5_c25_8 = t_r5_c25_4 + p_6_24;
  assign t_r5_c25_9 = t_r5_c25_5 + t_r5_c25_6;
  assign t_r5_c25_10 = t_r5_c25_7 + t_r5_c25_8;
  assign t_r5_c25_11 = t_r5_c25_9 + t_r5_c25_10;
  assign t_r5_c25_12 = t_r5_c25_11 + p_6_26;
  assign out_5_25 = t_r5_c25_12 >> 4;

  assign t_r5_c26_0 = p_4_26 << 1;
  assign t_r5_c26_1 = p_5_25 << 1;
  assign t_r5_c26_2 = p_5_26 << 2;
  assign t_r5_c26_3 = p_5_27 << 1;
  assign t_r5_c26_4 = p_6_26 << 1;
  assign t_r5_c26_5 = t_r5_c26_0 + p_4_25;
  assign t_r5_c26_6 = t_r5_c26_1 + p_4_27;
  assign t_r5_c26_7 = t_r5_c26_2 + t_r5_c26_3;
  assign t_r5_c26_8 = t_r5_c26_4 + p_6_25;
  assign t_r5_c26_9 = t_r5_c26_5 + t_r5_c26_6;
  assign t_r5_c26_10 = t_r5_c26_7 + t_r5_c26_8;
  assign t_r5_c26_11 = t_r5_c26_9 + t_r5_c26_10;
  assign t_r5_c26_12 = t_r5_c26_11 + p_6_27;
  assign out_5_26 = t_r5_c26_12 >> 4;

  assign t_r5_c27_0 = p_4_27 << 1;
  assign t_r5_c27_1 = p_5_26 << 1;
  assign t_r5_c27_2 = p_5_27 << 2;
  assign t_r5_c27_3 = p_5_28 << 1;
  assign t_r5_c27_4 = p_6_27 << 1;
  assign t_r5_c27_5 = t_r5_c27_0 + p_4_26;
  assign t_r5_c27_6 = t_r5_c27_1 + p_4_28;
  assign t_r5_c27_7 = t_r5_c27_2 + t_r5_c27_3;
  assign t_r5_c27_8 = t_r5_c27_4 + p_6_26;
  assign t_r5_c27_9 = t_r5_c27_5 + t_r5_c27_6;
  assign t_r5_c27_10 = t_r5_c27_7 + t_r5_c27_8;
  assign t_r5_c27_11 = t_r5_c27_9 + t_r5_c27_10;
  assign t_r5_c27_12 = t_r5_c27_11 + p_6_28;
  assign out_5_27 = t_r5_c27_12 >> 4;

  assign t_r5_c28_0 = p_4_28 << 1;
  assign t_r5_c28_1 = p_5_27 << 1;
  assign t_r5_c28_2 = p_5_28 << 2;
  assign t_r5_c28_3 = p_5_29 << 1;
  assign t_r5_c28_4 = p_6_28 << 1;
  assign t_r5_c28_5 = t_r5_c28_0 + p_4_27;
  assign t_r5_c28_6 = t_r5_c28_1 + p_4_29;
  assign t_r5_c28_7 = t_r5_c28_2 + t_r5_c28_3;
  assign t_r5_c28_8 = t_r5_c28_4 + p_6_27;
  assign t_r5_c28_9 = t_r5_c28_5 + t_r5_c28_6;
  assign t_r5_c28_10 = t_r5_c28_7 + t_r5_c28_8;
  assign t_r5_c28_11 = t_r5_c28_9 + t_r5_c28_10;
  assign t_r5_c28_12 = t_r5_c28_11 + p_6_29;
  assign out_5_28 = t_r5_c28_12 >> 4;

  assign t_r5_c29_0 = p_4_29 << 1;
  assign t_r5_c29_1 = p_5_28 << 1;
  assign t_r5_c29_2 = p_5_29 << 2;
  assign t_r5_c29_3 = p_5_30 << 1;
  assign t_r5_c29_4 = p_6_29 << 1;
  assign t_r5_c29_5 = t_r5_c29_0 + p_4_28;
  assign t_r5_c29_6 = t_r5_c29_1 + p_4_30;
  assign t_r5_c29_7 = t_r5_c29_2 + t_r5_c29_3;
  assign t_r5_c29_8 = t_r5_c29_4 + p_6_28;
  assign t_r5_c29_9 = t_r5_c29_5 + t_r5_c29_6;
  assign t_r5_c29_10 = t_r5_c29_7 + t_r5_c29_8;
  assign t_r5_c29_11 = t_r5_c29_9 + t_r5_c29_10;
  assign t_r5_c29_12 = t_r5_c29_11 + p_6_30;
  assign out_5_29 = t_r5_c29_12 >> 4;

  assign t_r5_c30_0 = p_4_30 << 1;
  assign t_r5_c30_1 = p_5_29 << 1;
  assign t_r5_c30_2 = p_5_30 << 2;
  assign t_r5_c30_3 = p_5_31 << 1;
  assign t_r5_c30_4 = p_6_30 << 1;
  assign t_r5_c30_5 = t_r5_c30_0 + p_4_29;
  assign t_r5_c30_6 = t_r5_c30_1 + p_4_31;
  assign t_r5_c30_7 = t_r5_c30_2 + t_r5_c30_3;
  assign t_r5_c30_8 = t_r5_c30_4 + p_6_29;
  assign t_r5_c30_9 = t_r5_c30_5 + t_r5_c30_6;
  assign t_r5_c30_10 = t_r5_c30_7 + t_r5_c30_8;
  assign t_r5_c30_11 = t_r5_c30_9 + t_r5_c30_10;
  assign t_r5_c30_12 = t_r5_c30_11 + p_6_31;
  assign out_5_30 = t_r5_c30_12 >> 4;

  assign t_r5_c31_0 = p_4_31 << 1;
  assign t_r5_c31_1 = p_5_30 << 1;
  assign t_r5_c31_2 = p_5_31 << 2;
  assign t_r5_c31_3 = p_5_32 << 1;
  assign t_r5_c31_4 = p_6_31 << 1;
  assign t_r5_c31_5 = t_r5_c31_0 + p_4_30;
  assign t_r5_c31_6 = t_r5_c31_1 + p_4_32;
  assign t_r5_c31_7 = t_r5_c31_2 + t_r5_c31_3;
  assign t_r5_c31_8 = t_r5_c31_4 + p_6_30;
  assign t_r5_c31_9 = t_r5_c31_5 + t_r5_c31_6;
  assign t_r5_c31_10 = t_r5_c31_7 + t_r5_c31_8;
  assign t_r5_c31_11 = t_r5_c31_9 + t_r5_c31_10;
  assign t_r5_c31_12 = t_r5_c31_11 + p_6_32;
  assign out_5_31 = t_r5_c31_12 >> 4;

  assign t_r5_c32_0 = p_4_32 << 1;
  assign t_r5_c32_1 = p_5_31 << 1;
  assign t_r5_c32_2 = p_5_32 << 2;
  assign t_r5_c32_3 = p_5_33 << 1;
  assign t_r5_c32_4 = p_6_32 << 1;
  assign t_r5_c32_5 = t_r5_c32_0 + p_4_31;
  assign t_r5_c32_6 = t_r5_c32_1 + p_4_33;
  assign t_r5_c32_7 = t_r5_c32_2 + t_r5_c32_3;
  assign t_r5_c32_8 = t_r5_c32_4 + p_6_31;
  assign t_r5_c32_9 = t_r5_c32_5 + t_r5_c32_6;
  assign t_r5_c32_10 = t_r5_c32_7 + t_r5_c32_8;
  assign t_r5_c32_11 = t_r5_c32_9 + t_r5_c32_10;
  assign t_r5_c32_12 = t_r5_c32_11 + p_6_33;
  assign out_5_32 = t_r5_c32_12 >> 4;

  assign t_r5_c33_0 = p_4_33 << 1;
  assign t_r5_c33_1 = p_5_32 << 1;
  assign t_r5_c33_2 = p_5_33 << 2;
  assign t_r5_c33_3 = p_5_34 << 1;
  assign t_r5_c33_4 = p_6_33 << 1;
  assign t_r5_c33_5 = t_r5_c33_0 + p_4_32;
  assign t_r5_c33_6 = t_r5_c33_1 + p_4_34;
  assign t_r5_c33_7 = t_r5_c33_2 + t_r5_c33_3;
  assign t_r5_c33_8 = t_r5_c33_4 + p_6_32;
  assign t_r5_c33_9 = t_r5_c33_5 + t_r5_c33_6;
  assign t_r5_c33_10 = t_r5_c33_7 + t_r5_c33_8;
  assign t_r5_c33_11 = t_r5_c33_9 + t_r5_c33_10;
  assign t_r5_c33_12 = t_r5_c33_11 + p_6_34;
  assign out_5_33 = t_r5_c33_12 >> 4;

  assign t_r5_c34_0 = p_4_34 << 1;
  assign t_r5_c34_1 = p_5_33 << 1;
  assign t_r5_c34_2 = p_5_34 << 2;
  assign t_r5_c34_3 = p_5_35 << 1;
  assign t_r5_c34_4 = p_6_34 << 1;
  assign t_r5_c34_5 = t_r5_c34_0 + p_4_33;
  assign t_r5_c34_6 = t_r5_c34_1 + p_4_35;
  assign t_r5_c34_7 = t_r5_c34_2 + t_r5_c34_3;
  assign t_r5_c34_8 = t_r5_c34_4 + p_6_33;
  assign t_r5_c34_9 = t_r5_c34_5 + t_r5_c34_6;
  assign t_r5_c34_10 = t_r5_c34_7 + t_r5_c34_8;
  assign t_r5_c34_11 = t_r5_c34_9 + t_r5_c34_10;
  assign t_r5_c34_12 = t_r5_c34_11 + p_6_35;
  assign out_5_34 = t_r5_c34_12 >> 4;

  assign t_r5_c35_0 = p_4_35 << 1;
  assign t_r5_c35_1 = p_5_34 << 1;
  assign t_r5_c35_2 = p_5_35 << 2;
  assign t_r5_c35_3 = p_5_36 << 1;
  assign t_r5_c35_4 = p_6_35 << 1;
  assign t_r5_c35_5 = t_r5_c35_0 + p_4_34;
  assign t_r5_c35_6 = t_r5_c35_1 + p_4_36;
  assign t_r5_c35_7 = t_r5_c35_2 + t_r5_c35_3;
  assign t_r5_c35_8 = t_r5_c35_4 + p_6_34;
  assign t_r5_c35_9 = t_r5_c35_5 + t_r5_c35_6;
  assign t_r5_c35_10 = t_r5_c35_7 + t_r5_c35_8;
  assign t_r5_c35_11 = t_r5_c35_9 + t_r5_c35_10;
  assign t_r5_c35_12 = t_r5_c35_11 + p_6_36;
  assign out_5_35 = t_r5_c35_12 >> 4;

  assign t_r5_c36_0 = p_4_36 << 1;
  assign t_r5_c36_1 = p_5_35 << 1;
  assign t_r5_c36_2 = p_5_36 << 2;
  assign t_r5_c36_3 = p_5_37 << 1;
  assign t_r5_c36_4 = p_6_36 << 1;
  assign t_r5_c36_5 = t_r5_c36_0 + p_4_35;
  assign t_r5_c36_6 = t_r5_c36_1 + p_4_37;
  assign t_r5_c36_7 = t_r5_c36_2 + t_r5_c36_3;
  assign t_r5_c36_8 = t_r5_c36_4 + p_6_35;
  assign t_r5_c36_9 = t_r5_c36_5 + t_r5_c36_6;
  assign t_r5_c36_10 = t_r5_c36_7 + t_r5_c36_8;
  assign t_r5_c36_11 = t_r5_c36_9 + t_r5_c36_10;
  assign t_r5_c36_12 = t_r5_c36_11 + p_6_37;
  assign out_5_36 = t_r5_c36_12 >> 4;

  assign t_r5_c37_0 = p_4_37 << 1;
  assign t_r5_c37_1 = p_5_36 << 1;
  assign t_r5_c37_2 = p_5_37 << 2;
  assign t_r5_c37_3 = p_5_38 << 1;
  assign t_r5_c37_4 = p_6_37 << 1;
  assign t_r5_c37_5 = t_r5_c37_0 + p_4_36;
  assign t_r5_c37_6 = t_r5_c37_1 + p_4_38;
  assign t_r5_c37_7 = t_r5_c37_2 + t_r5_c37_3;
  assign t_r5_c37_8 = t_r5_c37_4 + p_6_36;
  assign t_r5_c37_9 = t_r5_c37_5 + t_r5_c37_6;
  assign t_r5_c37_10 = t_r5_c37_7 + t_r5_c37_8;
  assign t_r5_c37_11 = t_r5_c37_9 + t_r5_c37_10;
  assign t_r5_c37_12 = t_r5_c37_11 + p_6_38;
  assign out_5_37 = t_r5_c37_12 >> 4;

  assign t_r5_c38_0 = p_4_38 << 1;
  assign t_r5_c38_1 = p_5_37 << 1;
  assign t_r5_c38_2 = p_5_38 << 2;
  assign t_r5_c38_3 = p_5_39 << 1;
  assign t_r5_c38_4 = p_6_38 << 1;
  assign t_r5_c38_5 = t_r5_c38_0 + p_4_37;
  assign t_r5_c38_6 = t_r5_c38_1 + p_4_39;
  assign t_r5_c38_7 = t_r5_c38_2 + t_r5_c38_3;
  assign t_r5_c38_8 = t_r5_c38_4 + p_6_37;
  assign t_r5_c38_9 = t_r5_c38_5 + t_r5_c38_6;
  assign t_r5_c38_10 = t_r5_c38_7 + t_r5_c38_8;
  assign t_r5_c38_11 = t_r5_c38_9 + t_r5_c38_10;
  assign t_r5_c38_12 = t_r5_c38_11 + p_6_39;
  assign out_5_38 = t_r5_c38_12 >> 4;

  assign t_r5_c39_0 = p_4_39 << 1;
  assign t_r5_c39_1 = p_5_38 << 1;
  assign t_r5_c39_2 = p_5_39 << 2;
  assign t_r5_c39_3 = p_5_40 << 1;
  assign t_r5_c39_4 = p_6_39 << 1;
  assign t_r5_c39_5 = t_r5_c39_0 + p_4_38;
  assign t_r5_c39_6 = t_r5_c39_1 + p_4_40;
  assign t_r5_c39_7 = t_r5_c39_2 + t_r5_c39_3;
  assign t_r5_c39_8 = t_r5_c39_4 + p_6_38;
  assign t_r5_c39_9 = t_r5_c39_5 + t_r5_c39_6;
  assign t_r5_c39_10 = t_r5_c39_7 + t_r5_c39_8;
  assign t_r5_c39_11 = t_r5_c39_9 + t_r5_c39_10;
  assign t_r5_c39_12 = t_r5_c39_11 + p_6_40;
  assign out_5_39 = t_r5_c39_12 >> 4;

  assign t_r5_c40_0 = p_4_40 << 1;
  assign t_r5_c40_1 = p_5_39 << 1;
  assign t_r5_c40_2 = p_5_40 << 2;
  assign t_r5_c40_3 = p_5_41 << 1;
  assign t_r5_c40_4 = p_6_40 << 1;
  assign t_r5_c40_5 = t_r5_c40_0 + p_4_39;
  assign t_r5_c40_6 = t_r5_c40_1 + p_4_41;
  assign t_r5_c40_7 = t_r5_c40_2 + t_r5_c40_3;
  assign t_r5_c40_8 = t_r5_c40_4 + p_6_39;
  assign t_r5_c40_9 = t_r5_c40_5 + t_r5_c40_6;
  assign t_r5_c40_10 = t_r5_c40_7 + t_r5_c40_8;
  assign t_r5_c40_11 = t_r5_c40_9 + t_r5_c40_10;
  assign t_r5_c40_12 = t_r5_c40_11 + p_6_41;
  assign out_5_40 = t_r5_c40_12 >> 4;

  assign t_r5_c41_0 = p_4_41 << 1;
  assign t_r5_c41_1 = p_5_40 << 1;
  assign t_r5_c41_2 = p_5_41 << 2;
  assign t_r5_c41_3 = p_5_42 << 1;
  assign t_r5_c41_4 = p_6_41 << 1;
  assign t_r5_c41_5 = t_r5_c41_0 + p_4_40;
  assign t_r5_c41_6 = t_r5_c41_1 + p_4_42;
  assign t_r5_c41_7 = t_r5_c41_2 + t_r5_c41_3;
  assign t_r5_c41_8 = t_r5_c41_4 + p_6_40;
  assign t_r5_c41_9 = t_r5_c41_5 + t_r5_c41_6;
  assign t_r5_c41_10 = t_r5_c41_7 + t_r5_c41_8;
  assign t_r5_c41_11 = t_r5_c41_9 + t_r5_c41_10;
  assign t_r5_c41_12 = t_r5_c41_11 + p_6_42;
  assign out_5_41 = t_r5_c41_12 >> 4;

  assign t_r5_c42_0 = p_4_42 << 1;
  assign t_r5_c42_1 = p_5_41 << 1;
  assign t_r5_c42_2 = p_5_42 << 2;
  assign t_r5_c42_3 = p_5_43 << 1;
  assign t_r5_c42_4 = p_6_42 << 1;
  assign t_r5_c42_5 = t_r5_c42_0 + p_4_41;
  assign t_r5_c42_6 = t_r5_c42_1 + p_4_43;
  assign t_r5_c42_7 = t_r5_c42_2 + t_r5_c42_3;
  assign t_r5_c42_8 = t_r5_c42_4 + p_6_41;
  assign t_r5_c42_9 = t_r5_c42_5 + t_r5_c42_6;
  assign t_r5_c42_10 = t_r5_c42_7 + t_r5_c42_8;
  assign t_r5_c42_11 = t_r5_c42_9 + t_r5_c42_10;
  assign t_r5_c42_12 = t_r5_c42_11 + p_6_43;
  assign out_5_42 = t_r5_c42_12 >> 4;

  assign t_r5_c43_0 = p_4_43 << 1;
  assign t_r5_c43_1 = p_5_42 << 1;
  assign t_r5_c43_2 = p_5_43 << 2;
  assign t_r5_c43_3 = p_5_44 << 1;
  assign t_r5_c43_4 = p_6_43 << 1;
  assign t_r5_c43_5 = t_r5_c43_0 + p_4_42;
  assign t_r5_c43_6 = t_r5_c43_1 + p_4_44;
  assign t_r5_c43_7 = t_r5_c43_2 + t_r5_c43_3;
  assign t_r5_c43_8 = t_r5_c43_4 + p_6_42;
  assign t_r5_c43_9 = t_r5_c43_5 + t_r5_c43_6;
  assign t_r5_c43_10 = t_r5_c43_7 + t_r5_c43_8;
  assign t_r5_c43_11 = t_r5_c43_9 + t_r5_c43_10;
  assign t_r5_c43_12 = t_r5_c43_11 + p_6_44;
  assign out_5_43 = t_r5_c43_12 >> 4;

  assign t_r5_c44_0 = p_4_44 << 1;
  assign t_r5_c44_1 = p_5_43 << 1;
  assign t_r5_c44_2 = p_5_44 << 2;
  assign t_r5_c44_3 = p_5_45 << 1;
  assign t_r5_c44_4 = p_6_44 << 1;
  assign t_r5_c44_5 = t_r5_c44_0 + p_4_43;
  assign t_r5_c44_6 = t_r5_c44_1 + p_4_45;
  assign t_r5_c44_7 = t_r5_c44_2 + t_r5_c44_3;
  assign t_r5_c44_8 = t_r5_c44_4 + p_6_43;
  assign t_r5_c44_9 = t_r5_c44_5 + t_r5_c44_6;
  assign t_r5_c44_10 = t_r5_c44_7 + t_r5_c44_8;
  assign t_r5_c44_11 = t_r5_c44_9 + t_r5_c44_10;
  assign t_r5_c44_12 = t_r5_c44_11 + p_6_45;
  assign out_5_44 = t_r5_c44_12 >> 4;

  assign t_r5_c45_0 = p_4_45 << 1;
  assign t_r5_c45_1 = p_5_44 << 1;
  assign t_r5_c45_2 = p_5_45 << 2;
  assign t_r5_c45_3 = p_5_46 << 1;
  assign t_r5_c45_4 = p_6_45 << 1;
  assign t_r5_c45_5 = t_r5_c45_0 + p_4_44;
  assign t_r5_c45_6 = t_r5_c45_1 + p_4_46;
  assign t_r5_c45_7 = t_r5_c45_2 + t_r5_c45_3;
  assign t_r5_c45_8 = t_r5_c45_4 + p_6_44;
  assign t_r5_c45_9 = t_r5_c45_5 + t_r5_c45_6;
  assign t_r5_c45_10 = t_r5_c45_7 + t_r5_c45_8;
  assign t_r5_c45_11 = t_r5_c45_9 + t_r5_c45_10;
  assign t_r5_c45_12 = t_r5_c45_11 + p_6_46;
  assign out_5_45 = t_r5_c45_12 >> 4;

  assign t_r5_c46_0 = p_4_46 << 1;
  assign t_r5_c46_1 = p_5_45 << 1;
  assign t_r5_c46_2 = p_5_46 << 2;
  assign t_r5_c46_3 = p_5_47 << 1;
  assign t_r5_c46_4 = p_6_46 << 1;
  assign t_r5_c46_5 = t_r5_c46_0 + p_4_45;
  assign t_r5_c46_6 = t_r5_c46_1 + p_4_47;
  assign t_r5_c46_7 = t_r5_c46_2 + t_r5_c46_3;
  assign t_r5_c46_8 = t_r5_c46_4 + p_6_45;
  assign t_r5_c46_9 = t_r5_c46_5 + t_r5_c46_6;
  assign t_r5_c46_10 = t_r5_c46_7 + t_r5_c46_8;
  assign t_r5_c46_11 = t_r5_c46_9 + t_r5_c46_10;
  assign t_r5_c46_12 = t_r5_c46_11 + p_6_47;
  assign out_5_46 = t_r5_c46_12 >> 4;

  assign t_r5_c47_0 = p_4_47 << 1;
  assign t_r5_c47_1 = p_5_46 << 1;
  assign t_r5_c47_2 = p_5_47 << 2;
  assign t_r5_c47_3 = p_5_48 << 1;
  assign t_r5_c47_4 = p_6_47 << 1;
  assign t_r5_c47_5 = t_r5_c47_0 + p_4_46;
  assign t_r5_c47_6 = t_r5_c47_1 + p_4_48;
  assign t_r5_c47_7 = t_r5_c47_2 + t_r5_c47_3;
  assign t_r5_c47_8 = t_r5_c47_4 + p_6_46;
  assign t_r5_c47_9 = t_r5_c47_5 + t_r5_c47_6;
  assign t_r5_c47_10 = t_r5_c47_7 + t_r5_c47_8;
  assign t_r5_c47_11 = t_r5_c47_9 + t_r5_c47_10;
  assign t_r5_c47_12 = t_r5_c47_11 + p_6_48;
  assign out_5_47 = t_r5_c47_12 >> 4;

  assign t_r5_c48_0 = p_4_48 << 1;
  assign t_r5_c48_1 = p_5_47 << 1;
  assign t_r5_c48_2 = p_5_48 << 2;
  assign t_r5_c48_3 = p_5_49 << 1;
  assign t_r5_c48_4 = p_6_48 << 1;
  assign t_r5_c48_5 = t_r5_c48_0 + p_4_47;
  assign t_r5_c48_6 = t_r5_c48_1 + p_4_49;
  assign t_r5_c48_7 = t_r5_c48_2 + t_r5_c48_3;
  assign t_r5_c48_8 = t_r5_c48_4 + p_6_47;
  assign t_r5_c48_9 = t_r5_c48_5 + t_r5_c48_6;
  assign t_r5_c48_10 = t_r5_c48_7 + t_r5_c48_8;
  assign t_r5_c48_11 = t_r5_c48_9 + t_r5_c48_10;
  assign t_r5_c48_12 = t_r5_c48_11 + p_6_49;
  assign out_5_48 = t_r5_c48_12 >> 4;

  assign t_r5_c49_0 = p_4_49 << 1;
  assign t_r5_c49_1 = p_5_48 << 1;
  assign t_r5_c49_2 = p_5_49 << 2;
  assign t_r5_c49_3 = p_5_50 << 1;
  assign t_r5_c49_4 = p_6_49 << 1;
  assign t_r5_c49_5 = t_r5_c49_0 + p_4_48;
  assign t_r5_c49_6 = t_r5_c49_1 + p_4_50;
  assign t_r5_c49_7 = t_r5_c49_2 + t_r5_c49_3;
  assign t_r5_c49_8 = t_r5_c49_4 + p_6_48;
  assign t_r5_c49_9 = t_r5_c49_5 + t_r5_c49_6;
  assign t_r5_c49_10 = t_r5_c49_7 + t_r5_c49_8;
  assign t_r5_c49_11 = t_r5_c49_9 + t_r5_c49_10;
  assign t_r5_c49_12 = t_r5_c49_11 + p_6_50;
  assign out_5_49 = t_r5_c49_12 >> 4;

  assign t_r5_c50_0 = p_4_50 << 1;
  assign t_r5_c50_1 = p_5_49 << 1;
  assign t_r5_c50_2 = p_5_50 << 2;
  assign t_r5_c50_3 = p_5_51 << 1;
  assign t_r5_c50_4 = p_6_50 << 1;
  assign t_r5_c50_5 = t_r5_c50_0 + p_4_49;
  assign t_r5_c50_6 = t_r5_c50_1 + p_4_51;
  assign t_r5_c50_7 = t_r5_c50_2 + t_r5_c50_3;
  assign t_r5_c50_8 = t_r5_c50_4 + p_6_49;
  assign t_r5_c50_9 = t_r5_c50_5 + t_r5_c50_6;
  assign t_r5_c50_10 = t_r5_c50_7 + t_r5_c50_8;
  assign t_r5_c50_11 = t_r5_c50_9 + t_r5_c50_10;
  assign t_r5_c50_12 = t_r5_c50_11 + p_6_51;
  assign out_5_50 = t_r5_c50_12 >> 4;

  assign t_r5_c51_0 = p_4_51 << 1;
  assign t_r5_c51_1 = p_5_50 << 1;
  assign t_r5_c51_2 = p_5_51 << 2;
  assign t_r5_c51_3 = p_5_52 << 1;
  assign t_r5_c51_4 = p_6_51 << 1;
  assign t_r5_c51_5 = t_r5_c51_0 + p_4_50;
  assign t_r5_c51_6 = t_r5_c51_1 + p_4_52;
  assign t_r5_c51_7 = t_r5_c51_2 + t_r5_c51_3;
  assign t_r5_c51_8 = t_r5_c51_4 + p_6_50;
  assign t_r5_c51_9 = t_r5_c51_5 + t_r5_c51_6;
  assign t_r5_c51_10 = t_r5_c51_7 + t_r5_c51_8;
  assign t_r5_c51_11 = t_r5_c51_9 + t_r5_c51_10;
  assign t_r5_c51_12 = t_r5_c51_11 + p_6_52;
  assign out_5_51 = t_r5_c51_12 >> 4;

  assign t_r5_c52_0 = p_4_52 << 1;
  assign t_r5_c52_1 = p_5_51 << 1;
  assign t_r5_c52_2 = p_5_52 << 2;
  assign t_r5_c52_3 = p_5_53 << 1;
  assign t_r5_c52_4 = p_6_52 << 1;
  assign t_r5_c52_5 = t_r5_c52_0 + p_4_51;
  assign t_r5_c52_6 = t_r5_c52_1 + p_4_53;
  assign t_r5_c52_7 = t_r5_c52_2 + t_r5_c52_3;
  assign t_r5_c52_8 = t_r5_c52_4 + p_6_51;
  assign t_r5_c52_9 = t_r5_c52_5 + t_r5_c52_6;
  assign t_r5_c52_10 = t_r5_c52_7 + t_r5_c52_8;
  assign t_r5_c52_11 = t_r5_c52_9 + t_r5_c52_10;
  assign t_r5_c52_12 = t_r5_c52_11 + p_6_53;
  assign out_5_52 = t_r5_c52_12 >> 4;

  assign t_r5_c53_0 = p_4_53 << 1;
  assign t_r5_c53_1 = p_5_52 << 1;
  assign t_r5_c53_2 = p_5_53 << 2;
  assign t_r5_c53_3 = p_5_54 << 1;
  assign t_r5_c53_4 = p_6_53 << 1;
  assign t_r5_c53_5 = t_r5_c53_0 + p_4_52;
  assign t_r5_c53_6 = t_r5_c53_1 + p_4_54;
  assign t_r5_c53_7 = t_r5_c53_2 + t_r5_c53_3;
  assign t_r5_c53_8 = t_r5_c53_4 + p_6_52;
  assign t_r5_c53_9 = t_r5_c53_5 + t_r5_c53_6;
  assign t_r5_c53_10 = t_r5_c53_7 + t_r5_c53_8;
  assign t_r5_c53_11 = t_r5_c53_9 + t_r5_c53_10;
  assign t_r5_c53_12 = t_r5_c53_11 + p_6_54;
  assign out_5_53 = t_r5_c53_12 >> 4;

  assign t_r5_c54_0 = p_4_54 << 1;
  assign t_r5_c54_1 = p_5_53 << 1;
  assign t_r5_c54_2 = p_5_54 << 2;
  assign t_r5_c54_3 = p_5_55 << 1;
  assign t_r5_c54_4 = p_6_54 << 1;
  assign t_r5_c54_5 = t_r5_c54_0 + p_4_53;
  assign t_r5_c54_6 = t_r5_c54_1 + p_4_55;
  assign t_r5_c54_7 = t_r5_c54_2 + t_r5_c54_3;
  assign t_r5_c54_8 = t_r5_c54_4 + p_6_53;
  assign t_r5_c54_9 = t_r5_c54_5 + t_r5_c54_6;
  assign t_r5_c54_10 = t_r5_c54_7 + t_r5_c54_8;
  assign t_r5_c54_11 = t_r5_c54_9 + t_r5_c54_10;
  assign t_r5_c54_12 = t_r5_c54_11 + p_6_55;
  assign out_5_54 = t_r5_c54_12 >> 4;

  assign t_r5_c55_0 = p_4_55 << 1;
  assign t_r5_c55_1 = p_5_54 << 1;
  assign t_r5_c55_2 = p_5_55 << 2;
  assign t_r5_c55_3 = p_5_56 << 1;
  assign t_r5_c55_4 = p_6_55 << 1;
  assign t_r5_c55_5 = t_r5_c55_0 + p_4_54;
  assign t_r5_c55_6 = t_r5_c55_1 + p_4_56;
  assign t_r5_c55_7 = t_r5_c55_2 + t_r5_c55_3;
  assign t_r5_c55_8 = t_r5_c55_4 + p_6_54;
  assign t_r5_c55_9 = t_r5_c55_5 + t_r5_c55_6;
  assign t_r5_c55_10 = t_r5_c55_7 + t_r5_c55_8;
  assign t_r5_c55_11 = t_r5_c55_9 + t_r5_c55_10;
  assign t_r5_c55_12 = t_r5_c55_11 + p_6_56;
  assign out_5_55 = t_r5_c55_12 >> 4;

  assign t_r5_c56_0 = p_4_56 << 1;
  assign t_r5_c56_1 = p_5_55 << 1;
  assign t_r5_c56_2 = p_5_56 << 2;
  assign t_r5_c56_3 = p_5_57 << 1;
  assign t_r5_c56_4 = p_6_56 << 1;
  assign t_r5_c56_5 = t_r5_c56_0 + p_4_55;
  assign t_r5_c56_6 = t_r5_c56_1 + p_4_57;
  assign t_r5_c56_7 = t_r5_c56_2 + t_r5_c56_3;
  assign t_r5_c56_8 = t_r5_c56_4 + p_6_55;
  assign t_r5_c56_9 = t_r5_c56_5 + t_r5_c56_6;
  assign t_r5_c56_10 = t_r5_c56_7 + t_r5_c56_8;
  assign t_r5_c56_11 = t_r5_c56_9 + t_r5_c56_10;
  assign t_r5_c56_12 = t_r5_c56_11 + p_6_57;
  assign out_5_56 = t_r5_c56_12 >> 4;

  assign t_r5_c57_0 = p_4_57 << 1;
  assign t_r5_c57_1 = p_5_56 << 1;
  assign t_r5_c57_2 = p_5_57 << 2;
  assign t_r5_c57_3 = p_5_58 << 1;
  assign t_r5_c57_4 = p_6_57 << 1;
  assign t_r5_c57_5 = t_r5_c57_0 + p_4_56;
  assign t_r5_c57_6 = t_r5_c57_1 + p_4_58;
  assign t_r5_c57_7 = t_r5_c57_2 + t_r5_c57_3;
  assign t_r5_c57_8 = t_r5_c57_4 + p_6_56;
  assign t_r5_c57_9 = t_r5_c57_5 + t_r5_c57_6;
  assign t_r5_c57_10 = t_r5_c57_7 + t_r5_c57_8;
  assign t_r5_c57_11 = t_r5_c57_9 + t_r5_c57_10;
  assign t_r5_c57_12 = t_r5_c57_11 + p_6_58;
  assign out_5_57 = t_r5_c57_12 >> 4;

  assign t_r5_c58_0 = p_4_58 << 1;
  assign t_r5_c58_1 = p_5_57 << 1;
  assign t_r5_c58_2 = p_5_58 << 2;
  assign t_r5_c58_3 = p_5_59 << 1;
  assign t_r5_c58_4 = p_6_58 << 1;
  assign t_r5_c58_5 = t_r5_c58_0 + p_4_57;
  assign t_r5_c58_6 = t_r5_c58_1 + p_4_59;
  assign t_r5_c58_7 = t_r5_c58_2 + t_r5_c58_3;
  assign t_r5_c58_8 = t_r5_c58_4 + p_6_57;
  assign t_r5_c58_9 = t_r5_c58_5 + t_r5_c58_6;
  assign t_r5_c58_10 = t_r5_c58_7 + t_r5_c58_8;
  assign t_r5_c58_11 = t_r5_c58_9 + t_r5_c58_10;
  assign t_r5_c58_12 = t_r5_c58_11 + p_6_59;
  assign out_5_58 = t_r5_c58_12 >> 4;

  assign t_r5_c59_0 = p_4_59 << 1;
  assign t_r5_c59_1 = p_5_58 << 1;
  assign t_r5_c59_2 = p_5_59 << 2;
  assign t_r5_c59_3 = p_5_60 << 1;
  assign t_r5_c59_4 = p_6_59 << 1;
  assign t_r5_c59_5 = t_r5_c59_0 + p_4_58;
  assign t_r5_c59_6 = t_r5_c59_1 + p_4_60;
  assign t_r5_c59_7 = t_r5_c59_2 + t_r5_c59_3;
  assign t_r5_c59_8 = t_r5_c59_4 + p_6_58;
  assign t_r5_c59_9 = t_r5_c59_5 + t_r5_c59_6;
  assign t_r5_c59_10 = t_r5_c59_7 + t_r5_c59_8;
  assign t_r5_c59_11 = t_r5_c59_9 + t_r5_c59_10;
  assign t_r5_c59_12 = t_r5_c59_11 + p_6_60;
  assign out_5_59 = t_r5_c59_12 >> 4;

  assign t_r5_c60_0 = p_4_60 << 1;
  assign t_r5_c60_1 = p_5_59 << 1;
  assign t_r5_c60_2 = p_5_60 << 2;
  assign t_r5_c60_3 = p_5_61 << 1;
  assign t_r5_c60_4 = p_6_60 << 1;
  assign t_r5_c60_5 = t_r5_c60_0 + p_4_59;
  assign t_r5_c60_6 = t_r5_c60_1 + p_4_61;
  assign t_r5_c60_7 = t_r5_c60_2 + t_r5_c60_3;
  assign t_r5_c60_8 = t_r5_c60_4 + p_6_59;
  assign t_r5_c60_9 = t_r5_c60_5 + t_r5_c60_6;
  assign t_r5_c60_10 = t_r5_c60_7 + t_r5_c60_8;
  assign t_r5_c60_11 = t_r5_c60_9 + t_r5_c60_10;
  assign t_r5_c60_12 = t_r5_c60_11 + p_6_61;
  assign out_5_60 = t_r5_c60_12 >> 4;

  assign t_r5_c61_0 = p_4_61 << 1;
  assign t_r5_c61_1 = p_5_60 << 1;
  assign t_r5_c61_2 = p_5_61 << 2;
  assign t_r5_c61_3 = p_5_62 << 1;
  assign t_r5_c61_4 = p_6_61 << 1;
  assign t_r5_c61_5 = t_r5_c61_0 + p_4_60;
  assign t_r5_c61_6 = t_r5_c61_1 + p_4_62;
  assign t_r5_c61_7 = t_r5_c61_2 + t_r5_c61_3;
  assign t_r5_c61_8 = t_r5_c61_4 + p_6_60;
  assign t_r5_c61_9 = t_r5_c61_5 + t_r5_c61_6;
  assign t_r5_c61_10 = t_r5_c61_7 + t_r5_c61_8;
  assign t_r5_c61_11 = t_r5_c61_9 + t_r5_c61_10;
  assign t_r5_c61_12 = t_r5_c61_11 + p_6_62;
  assign out_5_61 = t_r5_c61_12 >> 4;

  assign t_r5_c62_0 = p_4_62 << 1;
  assign t_r5_c62_1 = p_5_61 << 1;
  assign t_r5_c62_2 = p_5_62 << 2;
  assign t_r5_c62_3 = p_5_63 << 1;
  assign t_r5_c62_4 = p_6_62 << 1;
  assign t_r5_c62_5 = t_r5_c62_0 + p_4_61;
  assign t_r5_c62_6 = t_r5_c62_1 + p_4_63;
  assign t_r5_c62_7 = t_r5_c62_2 + t_r5_c62_3;
  assign t_r5_c62_8 = t_r5_c62_4 + p_6_61;
  assign t_r5_c62_9 = t_r5_c62_5 + t_r5_c62_6;
  assign t_r5_c62_10 = t_r5_c62_7 + t_r5_c62_8;
  assign t_r5_c62_11 = t_r5_c62_9 + t_r5_c62_10;
  assign t_r5_c62_12 = t_r5_c62_11 + p_6_63;
  assign out_5_62 = t_r5_c62_12 >> 4;

  assign t_r5_c63_0 = p_4_63 << 1;
  assign t_r5_c63_1 = p_5_62 << 1;
  assign t_r5_c63_2 = p_5_63 << 2;
  assign t_r5_c63_3 = p_5_64 << 1;
  assign t_r5_c63_4 = p_6_63 << 1;
  assign t_r5_c63_5 = t_r5_c63_0 + p_4_62;
  assign t_r5_c63_6 = t_r5_c63_1 + p_4_64;
  assign t_r5_c63_7 = t_r5_c63_2 + t_r5_c63_3;
  assign t_r5_c63_8 = t_r5_c63_4 + p_6_62;
  assign t_r5_c63_9 = t_r5_c63_5 + t_r5_c63_6;
  assign t_r5_c63_10 = t_r5_c63_7 + t_r5_c63_8;
  assign t_r5_c63_11 = t_r5_c63_9 + t_r5_c63_10;
  assign t_r5_c63_12 = t_r5_c63_11 + p_6_64;
  assign out_5_63 = t_r5_c63_12 >> 4;

  assign t_r5_c64_0 = p_4_64 << 1;
  assign t_r5_c64_1 = p_5_63 << 1;
  assign t_r5_c64_2 = p_5_64 << 2;
  assign t_r5_c64_3 = p_5_65 << 1;
  assign t_r5_c64_4 = p_6_64 << 1;
  assign t_r5_c64_5 = t_r5_c64_0 + p_4_63;
  assign t_r5_c64_6 = t_r5_c64_1 + p_4_65;
  assign t_r5_c64_7 = t_r5_c64_2 + t_r5_c64_3;
  assign t_r5_c64_8 = t_r5_c64_4 + p_6_63;
  assign t_r5_c64_9 = t_r5_c64_5 + t_r5_c64_6;
  assign t_r5_c64_10 = t_r5_c64_7 + t_r5_c64_8;
  assign t_r5_c64_11 = t_r5_c64_9 + t_r5_c64_10;
  assign t_r5_c64_12 = t_r5_c64_11 + p_6_65;
  assign out_5_64 = t_r5_c64_12 >> 4;

  assign t_r6_c1_0 = p_5_1 << 1;
  assign t_r6_c1_1 = p_6_0 << 1;
  assign t_r6_c1_2 = p_6_1 << 2;
  assign t_r6_c1_3 = p_6_2 << 1;
  assign t_r6_c1_4 = p_7_1 << 1;
  assign t_r6_c1_5 = t_r6_c1_0 + p_5_0;
  assign t_r6_c1_6 = t_r6_c1_1 + p_5_2;
  assign t_r6_c1_7 = t_r6_c1_2 + t_r6_c1_3;
  assign t_r6_c1_8 = t_r6_c1_4 + p_7_0;
  assign t_r6_c1_9 = t_r6_c1_5 + t_r6_c1_6;
  assign t_r6_c1_10 = t_r6_c1_7 + t_r6_c1_8;
  assign t_r6_c1_11 = t_r6_c1_9 + t_r6_c1_10;
  assign t_r6_c1_12 = t_r6_c1_11 + p_7_2;
  assign out_6_1 = t_r6_c1_12 >> 4;

  assign t_r6_c2_0 = p_5_2 << 1;
  assign t_r6_c2_1 = p_6_1 << 1;
  assign t_r6_c2_2 = p_6_2 << 2;
  assign t_r6_c2_3 = p_6_3 << 1;
  assign t_r6_c2_4 = p_7_2 << 1;
  assign t_r6_c2_5 = t_r6_c2_0 + p_5_1;
  assign t_r6_c2_6 = t_r6_c2_1 + p_5_3;
  assign t_r6_c2_7 = t_r6_c2_2 + t_r6_c2_3;
  assign t_r6_c2_8 = t_r6_c2_4 + p_7_1;
  assign t_r6_c2_9 = t_r6_c2_5 + t_r6_c2_6;
  assign t_r6_c2_10 = t_r6_c2_7 + t_r6_c2_8;
  assign t_r6_c2_11 = t_r6_c2_9 + t_r6_c2_10;
  assign t_r6_c2_12 = t_r6_c2_11 + p_7_3;
  assign out_6_2 = t_r6_c2_12 >> 4;

  assign t_r6_c3_0 = p_5_3 << 1;
  assign t_r6_c3_1 = p_6_2 << 1;
  assign t_r6_c3_2 = p_6_3 << 2;
  assign t_r6_c3_3 = p_6_4 << 1;
  assign t_r6_c3_4 = p_7_3 << 1;
  assign t_r6_c3_5 = t_r6_c3_0 + p_5_2;
  assign t_r6_c3_6 = t_r6_c3_1 + p_5_4;
  assign t_r6_c3_7 = t_r6_c3_2 + t_r6_c3_3;
  assign t_r6_c3_8 = t_r6_c3_4 + p_7_2;
  assign t_r6_c3_9 = t_r6_c3_5 + t_r6_c3_6;
  assign t_r6_c3_10 = t_r6_c3_7 + t_r6_c3_8;
  assign t_r6_c3_11 = t_r6_c3_9 + t_r6_c3_10;
  assign t_r6_c3_12 = t_r6_c3_11 + p_7_4;
  assign out_6_3 = t_r6_c3_12 >> 4;

  assign t_r6_c4_0 = p_5_4 << 1;
  assign t_r6_c4_1 = p_6_3 << 1;
  assign t_r6_c4_2 = p_6_4 << 2;
  assign t_r6_c4_3 = p_6_5 << 1;
  assign t_r6_c4_4 = p_7_4 << 1;
  assign t_r6_c4_5 = t_r6_c4_0 + p_5_3;
  assign t_r6_c4_6 = t_r6_c4_1 + p_5_5;
  assign t_r6_c4_7 = t_r6_c4_2 + t_r6_c4_3;
  assign t_r6_c4_8 = t_r6_c4_4 + p_7_3;
  assign t_r6_c4_9 = t_r6_c4_5 + t_r6_c4_6;
  assign t_r6_c4_10 = t_r6_c4_7 + t_r6_c4_8;
  assign t_r6_c4_11 = t_r6_c4_9 + t_r6_c4_10;
  assign t_r6_c4_12 = t_r6_c4_11 + p_7_5;
  assign out_6_4 = t_r6_c4_12 >> 4;

  assign t_r6_c5_0 = p_5_5 << 1;
  assign t_r6_c5_1 = p_6_4 << 1;
  assign t_r6_c5_2 = p_6_5 << 2;
  assign t_r6_c5_3 = p_6_6 << 1;
  assign t_r6_c5_4 = p_7_5 << 1;
  assign t_r6_c5_5 = t_r6_c5_0 + p_5_4;
  assign t_r6_c5_6 = t_r6_c5_1 + p_5_6;
  assign t_r6_c5_7 = t_r6_c5_2 + t_r6_c5_3;
  assign t_r6_c5_8 = t_r6_c5_4 + p_7_4;
  assign t_r6_c5_9 = t_r6_c5_5 + t_r6_c5_6;
  assign t_r6_c5_10 = t_r6_c5_7 + t_r6_c5_8;
  assign t_r6_c5_11 = t_r6_c5_9 + t_r6_c5_10;
  assign t_r6_c5_12 = t_r6_c5_11 + p_7_6;
  assign out_6_5 = t_r6_c5_12 >> 4;

  assign t_r6_c6_0 = p_5_6 << 1;
  assign t_r6_c6_1 = p_6_5 << 1;
  assign t_r6_c6_2 = p_6_6 << 2;
  assign t_r6_c6_3 = p_6_7 << 1;
  assign t_r6_c6_4 = p_7_6 << 1;
  assign t_r6_c6_5 = t_r6_c6_0 + p_5_5;
  assign t_r6_c6_6 = t_r6_c6_1 + p_5_7;
  assign t_r6_c6_7 = t_r6_c6_2 + t_r6_c6_3;
  assign t_r6_c6_8 = t_r6_c6_4 + p_7_5;
  assign t_r6_c6_9 = t_r6_c6_5 + t_r6_c6_6;
  assign t_r6_c6_10 = t_r6_c6_7 + t_r6_c6_8;
  assign t_r6_c6_11 = t_r6_c6_9 + t_r6_c6_10;
  assign t_r6_c6_12 = t_r6_c6_11 + p_7_7;
  assign out_6_6 = t_r6_c6_12 >> 4;

  assign t_r6_c7_0 = p_5_7 << 1;
  assign t_r6_c7_1 = p_6_6 << 1;
  assign t_r6_c7_2 = p_6_7 << 2;
  assign t_r6_c7_3 = p_6_8 << 1;
  assign t_r6_c7_4 = p_7_7 << 1;
  assign t_r6_c7_5 = t_r6_c7_0 + p_5_6;
  assign t_r6_c7_6 = t_r6_c7_1 + p_5_8;
  assign t_r6_c7_7 = t_r6_c7_2 + t_r6_c7_3;
  assign t_r6_c7_8 = t_r6_c7_4 + p_7_6;
  assign t_r6_c7_9 = t_r6_c7_5 + t_r6_c7_6;
  assign t_r6_c7_10 = t_r6_c7_7 + t_r6_c7_8;
  assign t_r6_c7_11 = t_r6_c7_9 + t_r6_c7_10;
  assign t_r6_c7_12 = t_r6_c7_11 + p_7_8;
  assign out_6_7 = t_r6_c7_12 >> 4;

  assign t_r6_c8_0 = p_5_8 << 1;
  assign t_r6_c8_1 = p_6_7 << 1;
  assign t_r6_c8_2 = p_6_8 << 2;
  assign t_r6_c8_3 = p_6_9 << 1;
  assign t_r6_c8_4 = p_7_8 << 1;
  assign t_r6_c8_5 = t_r6_c8_0 + p_5_7;
  assign t_r6_c8_6 = t_r6_c8_1 + p_5_9;
  assign t_r6_c8_7 = t_r6_c8_2 + t_r6_c8_3;
  assign t_r6_c8_8 = t_r6_c8_4 + p_7_7;
  assign t_r6_c8_9 = t_r6_c8_5 + t_r6_c8_6;
  assign t_r6_c8_10 = t_r6_c8_7 + t_r6_c8_8;
  assign t_r6_c8_11 = t_r6_c8_9 + t_r6_c8_10;
  assign t_r6_c8_12 = t_r6_c8_11 + p_7_9;
  assign out_6_8 = t_r6_c8_12 >> 4;

  assign t_r6_c9_0 = p_5_9 << 1;
  assign t_r6_c9_1 = p_6_8 << 1;
  assign t_r6_c9_2 = p_6_9 << 2;
  assign t_r6_c9_3 = p_6_10 << 1;
  assign t_r6_c9_4 = p_7_9 << 1;
  assign t_r6_c9_5 = t_r6_c9_0 + p_5_8;
  assign t_r6_c9_6 = t_r6_c9_1 + p_5_10;
  assign t_r6_c9_7 = t_r6_c9_2 + t_r6_c9_3;
  assign t_r6_c9_8 = t_r6_c9_4 + p_7_8;
  assign t_r6_c9_9 = t_r6_c9_5 + t_r6_c9_6;
  assign t_r6_c9_10 = t_r6_c9_7 + t_r6_c9_8;
  assign t_r6_c9_11 = t_r6_c9_9 + t_r6_c9_10;
  assign t_r6_c9_12 = t_r6_c9_11 + p_7_10;
  assign out_6_9 = t_r6_c9_12 >> 4;

  assign t_r6_c10_0 = p_5_10 << 1;
  assign t_r6_c10_1 = p_6_9 << 1;
  assign t_r6_c10_2 = p_6_10 << 2;
  assign t_r6_c10_3 = p_6_11 << 1;
  assign t_r6_c10_4 = p_7_10 << 1;
  assign t_r6_c10_5 = t_r6_c10_0 + p_5_9;
  assign t_r6_c10_6 = t_r6_c10_1 + p_5_11;
  assign t_r6_c10_7 = t_r6_c10_2 + t_r6_c10_3;
  assign t_r6_c10_8 = t_r6_c10_4 + p_7_9;
  assign t_r6_c10_9 = t_r6_c10_5 + t_r6_c10_6;
  assign t_r6_c10_10 = t_r6_c10_7 + t_r6_c10_8;
  assign t_r6_c10_11 = t_r6_c10_9 + t_r6_c10_10;
  assign t_r6_c10_12 = t_r6_c10_11 + p_7_11;
  assign out_6_10 = t_r6_c10_12 >> 4;

  assign t_r6_c11_0 = p_5_11 << 1;
  assign t_r6_c11_1 = p_6_10 << 1;
  assign t_r6_c11_2 = p_6_11 << 2;
  assign t_r6_c11_3 = p_6_12 << 1;
  assign t_r6_c11_4 = p_7_11 << 1;
  assign t_r6_c11_5 = t_r6_c11_0 + p_5_10;
  assign t_r6_c11_6 = t_r6_c11_1 + p_5_12;
  assign t_r6_c11_7 = t_r6_c11_2 + t_r6_c11_3;
  assign t_r6_c11_8 = t_r6_c11_4 + p_7_10;
  assign t_r6_c11_9 = t_r6_c11_5 + t_r6_c11_6;
  assign t_r6_c11_10 = t_r6_c11_7 + t_r6_c11_8;
  assign t_r6_c11_11 = t_r6_c11_9 + t_r6_c11_10;
  assign t_r6_c11_12 = t_r6_c11_11 + p_7_12;
  assign out_6_11 = t_r6_c11_12 >> 4;

  assign t_r6_c12_0 = p_5_12 << 1;
  assign t_r6_c12_1 = p_6_11 << 1;
  assign t_r6_c12_2 = p_6_12 << 2;
  assign t_r6_c12_3 = p_6_13 << 1;
  assign t_r6_c12_4 = p_7_12 << 1;
  assign t_r6_c12_5 = t_r6_c12_0 + p_5_11;
  assign t_r6_c12_6 = t_r6_c12_1 + p_5_13;
  assign t_r6_c12_7 = t_r6_c12_2 + t_r6_c12_3;
  assign t_r6_c12_8 = t_r6_c12_4 + p_7_11;
  assign t_r6_c12_9 = t_r6_c12_5 + t_r6_c12_6;
  assign t_r6_c12_10 = t_r6_c12_7 + t_r6_c12_8;
  assign t_r6_c12_11 = t_r6_c12_9 + t_r6_c12_10;
  assign t_r6_c12_12 = t_r6_c12_11 + p_7_13;
  assign out_6_12 = t_r6_c12_12 >> 4;

  assign t_r6_c13_0 = p_5_13 << 1;
  assign t_r6_c13_1 = p_6_12 << 1;
  assign t_r6_c13_2 = p_6_13 << 2;
  assign t_r6_c13_3 = p_6_14 << 1;
  assign t_r6_c13_4 = p_7_13 << 1;
  assign t_r6_c13_5 = t_r6_c13_0 + p_5_12;
  assign t_r6_c13_6 = t_r6_c13_1 + p_5_14;
  assign t_r6_c13_7 = t_r6_c13_2 + t_r6_c13_3;
  assign t_r6_c13_8 = t_r6_c13_4 + p_7_12;
  assign t_r6_c13_9 = t_r6_c13_5 + t_r6_c13_6;
  assign t_r6_c13_10 = t_r6_c13_7 + t_r6_c13_8;
  assign t_r6_c13_11 = t_r6_c13_9 + t_r6_c13_10;
  assign t_r6_c13_12 = t_r6_c13_11 + p_7_14;
  assign out_6_13 = t_r6_c13_12 >> 4;

  assign t_r6_c14_0 = p_5_14 << 1;
  assign t_r6_c14_1 = p_6_13 << 1;
  assign t_r6_c14_2 = p_6_14 << 2;
  assign t_r6_c14_3 = p_6_15 << 1;
  assign t_r6_c14_4 = p_7_14 << 1;
  assign t_r6_c14_5 = t_r6_c14_0 + p_5_13;
  assign t_r6_c14_6 = t_r6_c14_1 + p_5_15;
  assign t_r6_c14_7 = t_r6_c14_2 + t_r6_c14_3;
  assign t_r6_c14_8 = t_r6_c14_4 + p_7_13;
  assign t_r6_c14_9 = t_r6_c14_5 + t_r6_c14_6;
  assign t_r6_c14_10 = t_r6_c14_7 + t_r6_c14_8;
  assign t_r6_c14_11 = t_r6_c14_9 + t_r6_c14_10;
  assign t_r6_c14_12 = t_r6_c14_11 + p_7_15;
  assign out_6_14 = t_r6_c14_12 >> 4;

  assign t_r6_c15_0 = p_5_15 << 1;
  assign t_r6_c15_1 = p_6_14 << 1;
  assign t_r6_c15_2 = p_6_15 << 2;
  assign t_r6_c15_3 = p_6_16 << 1;
  assign t_r6_c15_4 = p_7_15 << 1;
  assign t_r6_c15_5 = t_r6_c15_0 + p_5_14;
  assign t_r6_c15_6 = t_r6_c15_1 + p_5_16;
  assign t_r6_c15_7 = t_r6_c15_2 + t_r6_c15_3;
  assign t_r6_c15_8 = t_r6_c15_4 + p_7_14;
  assign t_r6_c15_9 = t_r6_c15_5 + t_r6_c15_6;
  assign t_r6_c15_10 = t_r6_c15_7 + t_r6_c15_8;
  assign t_r6_c15_11 = t_r6_c15_9 + t_r6_c15_10;
  assign t_r6_c15_12 = t_r6_c15_11 + p_7_16;
  assign out_6_15 = t_r6_c15_12 >> 4;

  assign t_r6_c16_0 = p_5_16 << 1;
  assign t_r6_c16_1 = p_6_15 << 1;
  assign t_r6_c16_2 = p_6_16 << 2;
  assign t_r6_c16_3 = p_6_17 << 1;
  assign t_r6_c16_4 = p_7_16 << 1;
  assign t_r6_c16_5 = t_r6_c16_0 + p_5_15;
  assign t_r6_c16_6 = t_r6_c16_1 + p_5_17;
  assign t_r6_c16_7 = t_r6_c16_2 + t_r6_c16_3;
  assign t_r6_c16_8 = t_r6_c16_4 + p_7_15;
  assign t_r6_c16_9 = t_r6_c16_5 + t_r6_c16_6;
  assign t_r6_c16_10 = t_r6_c16_7 + t_r6_c16_8;
  assign t_r6_c16_11 = t_r6_c16_9 + t_r6_c16_10;
  assign t_r6_c16_12 = t_r6_c16_11 + p_7_17;
  assign out_6_16 = t_r6_c16_12 >> 4;

  assign t_r6_c17_0 = p_5_17 << 1;
  assign t_r6_c17_1 = p_6_16 << 1;
  assign t_r6_c17_2 = p_6_17 << 2;
  assign t_r6_c17_3 = p_6_18 << 1;
  assign t_r6_c17_4 = p_7_17 << 1;
  assign t_r6_c17_5 = t_r6_c17_0 + p_5_16;
  assign t_r6_c17_6 = t_r6_c17_1 + p_5_18;
  assign t_r6_c17_7 = t_r6_c17_2 + t_r6_c17_3;
  assign t_r6_c17_8 = t_r6_c17_4 + p_7_16;
  assign t_r6_c17_9 = t_r6_c17_5 + t_r6_c17_6;
  assign t_r6_c17_10 = t_r6_c17_7 + t_r6_c17_8;
  assign t_r6_c17_11 = t_r6_c17_9 + t_r6_c17_10;
  assign t_r6_c17_12 = t_r6_c17_11 + p_7_18;
  assign out_6_17 = t_r6_c17_12 >> 4;

  assign t_r6_c18_0 = p_5_18 << 1;
  assign t_r6_c18_1 = p_6_17 << 1;
  assign t_r6_c18_2 = p_6_18 << 2;
  assign t_r6_c18_3 = p_6_19 << 1;
  assign t_r6_c18_4 = p_7_18 << 1;
  assign t_r6_c18_5 = t_r6_c18_0 + p_5_17;
  assign t_r6_c18_6 = t_r6_c18_1 + p_5_19;
  assign t_r6_c18_7 = t_r6_c18_2 + t_r6_c18_3;
  assign t_r6_c18_8 = t_r6_c18_4 + p_7_17;
  assign t_r6_c18_9 = t_r6_c18_5 + t_r6_c18_6;
  assign t_r6_c18_10 = t_r6_c18_7 + t_r6_c18_8;
  assign t_r6_c18_11 = t_r6_c18_9 + t_r6_c18_10;
  assign t_r6_c18_12 = t_r6_c18_11 + p_7_19;
  assign out_6_18 = t_r6_c18_12 >> 4;

  assign t_r6_c19_0 = p_5_19 << 1;
  assign t_r6_c19_1 = p_6_18 << 1;
  assign t_r6_c19_2 = p_6_19 << 2;
  assign t_r6_c19_3 = p_6_20 << 1;
  assign t_r6_c19_4 = p_7_19 << 1;
  assign t_r6_c19_5 = t_r6_c19_0 + p_5_18;
  assign t_r6_c19_6 = t_r6_c19_1 + p_5_20;
  assign t_r6_c19_7 = t_r6_c19_2 + t_r6_c19_3;
  assign t_r6_c19_8 = t_r6_c19_4 + p_7_18;
  assign t_r6_c19_9 = t_r6_c19_5 + t_r6_c19_6;
  assign t_r6_c19_10 = t_r6_c19_7 + t_r6_c19_8;
  assign t_r6_c19_11 = t_r6_c19_9 + t_r6_c19_10;
  assign t_r6_c19_12 = t_r6_c19_11 + p_7_20;
  assign out_6_19 = t_r6_c19_12 >> 4;

  assign t_r6_c20_0 = p_5_20 << 1;
  assign t_r6_c20_1 = p_6_19 << 1;
  assign t_r6_c20_2 = p_6_20 << 2;
  assign t_r6_c20_3 = p_6_21 << 1;
  assign t_r6_c20_4 = p_7_20 << 1;
  assign t_r6_c20_5 = t_r6_c20_0 + p_5_19;
  assign t_r6_c20_6 = t_r6_c20_1 + p_5_21;
  assign t_r6_c20_7 = t_r6_c20_2 + t_r6_c20_3;
  assign t_r6_c20_8 = t_r6_c20_4 + p_7_19;
  assign t_r6_c20_9 = t_r6_c20_5 + t_r6_c20_6;
  assign t_r6_c20_10 = t_r6_c20_7 + t_r6_c20_8;
  assign t_r6_c20_11 = t_r6_c20_9 + t_r6_c20_10;
  assign t_r6_c20_12 = t_r6_c20_11 + p_7_21;
  assign out_6_20 = t_r6_c20_12 >> 4;

  assign t_r6_c21_0 = p_5_21 << 1;
  assign t_r6_c21_1 = p_6_20 << 1;
  assign t_r6_c21_2 = p_6_21 << 2;
  assign t_r6_c21_3 = p_6_22 << 1;
  assign t_r6_c21_4 = p_7_21 << 1;
  assign t_r6_c21_5 = t_r6_c21_0 + p_5_20;
  assign t_r6_c21_6 = t_r6_c21_1 + p_5_22;
  assign t_r6_c21_7 = t_r6_c21_2 + t_r6_c21_3;
  assign t_r6_c21_8 = t_r6_c21_4 + p_7_20;
  assign t_r6_c21_9 = t_r6_c21_5 + t_r6_c21_6;
  assign t_r6_c21_10 = t_r6_c21_7 + t_r6_c21_8;
  assign t_r6_c21_11 = t_r6_c21_9 + t_r6_c21_10;
  assign t_r6_c21_12 = t_r6_c21_11 + p_7_22;
  assign out_6_21 = t_r6_c21_12 >> 4;

  assign t_r6_c22_0 = p_5_22 << 1;
  assign t_r6_c22_1 = p_6_21 << 1;
  assign t_r6_c22_2 = p_6_22 << 2;
  assign t_r6_c22_3 = p_6_23 << 1;
  assign t_r6_c22_4 = p_7_22 << 1;
  assign t_r6_c22_5 = t_r6_c22_0 + p_5_21;
  assign t_r6_c22_6 = t_r6_c22_1 + p_5_23;
  assign t_r6_c22_7 = t_r6_c22_2 + t_r6_c22_3;
  assign t_r6_c22_8 = t_r6_c22_4 + p_7_21;
  assign t_r6_c22_9 = t_r6_c22_5 + t_r6_c22_6;
  assign t_r6_c22_10 = t_r6_c22_7 + t_r6_c22_8;
  assign t_r6_c22_11 = t_r6_c22_9 + t_r6_c22_10;
  assign t_r6_c22_12 = t_r6_c22_11 + p_7_23;
  assign out_6_22 = t_r6_c22_12 >> 4;

  assign t_r6_c23_0 = p_5_23 << 1;
  assign t_r6_c23_1 = p_6_22 << 1;
  assign t_r6_c23_2 = p_6_23 << 2;
  assign t_r6_c23_3 = p_6_24 << 1;
  assign t_r6_c23_4 = p_7_23 << 1;
  assign t_r6_c23_5 = t_r6_c23_0 + p_5_22;
  assign t_r6_c23_6 = t_r6_c23_1 + p_5_24;
  assign t_r6_c23_7 = t_r6_c23_2 + t_r6_c23_3;
  assign t_r6_c23_8 = t_r6_c23_4 + p_7_22;
  assign t_r6_c23_9 = t_r6_c23_5 + t_r6_c23_6;
  assign t_r6_c23_10 = t_r6_c23_7 + t_r6_c23_8;
  assign t_r6_c23_11 = t_r6_c23_9 + t_r6_c23_10;
  assign t_r6_c23_12 = t_r6_c23_11 + p_7_24;
  assign out_6_23 = t_r6_c23_12 >> 4;

  assign t_r6_c24_0 = p_5_24 << 1;
  assign t_r6_c24_1 = p_6_23 << 1;
  assign t_r6_c24_2 = p_6_24 << 2;
  assign t_r6_c24_3 = p_6_25 << 1;
  assign t_r6_c24_4 = p_7_24 << 1;
  assign t_r6_c24_5 = t_r6_c24_0 + p_5_23;
  assign t_r6_c24_6 = t_r6_c24_1 + p_5_25;
  assign t_r6_c24_7 = t_r6_c24_2 + t_r6_c24_3;
  assign t_r6_c24_8 = t_r6_c24_4 + p_7_23;
  assign t_r6_c24_9 = t_r6_c24_5 + t_r6_c24_6;
  assign t_r6_c24_10 = t_r6_c24_7 + t_r6_c24_8;
  assign t_r6_c24_11 = t_r6_c24_9 + t_r6_c24_10;
  assign t_r6_c24_12 = t_r6_c24_11 + p_7_25;
  assign out_6_24 = t_r6_c24_12 >> 4;

  assign t_r6_c25_0 = p_5_25 << 1;
  assign t_r6_c25_1 = p_6_24 << 1;
  assign t_r6_c25_2 = p_6_25 << 2;
  assign t_r6_c25_3 = p_6_26 << 1;
  assign t_r6_c25_4 = p_7_25 << 1;
  assign t_r6_c25_5 = t_r6_c25_0 + p_5_24;
  assign t_r6_c25_6 = t_r6_c25_1 + p_5_26;
  assign t_r6_c25_7 = t_r6_c25_2 + t_r6_c25_3;
  assign t_r6_c25_8 = t_r6_c25_4 + p_7_24;
  assign t_r6_c25_9 = t_r6_c25_5 + t_r6_c25_6;
  assign t_r6_c25_10 = t_r6_c25_7 + t_r6_c25_8;
  assign t_r6_c25_11 = t_r6_c25_9 + t_r6_c25_10;
  assign t_r6_c25_12 = t_r6_c25_11 + p_7_26;
  assign out_6_25 = t_r6_c25_12 >> 4;

  assign t_r6_c26_0 = p_5_26 << 1;
  assign t_r6_c26_1 = p_6_25 << 1;
  assign t_r6_c26_2 = p_6_26 << 2;
  assign t_r6_c26_3 = p_6_27 << 1;
  assign t_r6_c26_4 = p_7_26 << 1;
  assign t_r6_c26_5 = t_r6_c26_0 + p_5_25;
  assign t_r6_c26_6 = t_r6_c26_1 + p_5_27;
  assign t_r6_c26_7 = t_r6_c26_2 + t_r6_c26_3;
  assign t_r6_c26_8 = t_r6_c26_4 + p_7_25;
  assign t_r6_c26_9 = t_r6_c26_5 + t_r6_c26_6;
  assign t_r6_c26_10 = t_r6_c26_7 + t_r6_c26_8;
  assign t_r6_c26_11 = t_r6_c26_9 + t_r6_c26_10;
  assign t_r6_c26_12 = t_r6_c26_11 + p_7_27;
  assign out_6_26 = t_r6_c26_12 >> 4;

  assign t_r6_c27_0 = p_5_27 << 1;
  assign t_r6_c27_1 = p_6_26 << 1;
  assign t_r6_c27_2 = p_6_27 << 2;
  assign t_r6_c27_3 = p_6_28 << 1;
  assign t_r6_c27_4 = p_7_27 << 1;
  assign t_r6_c27_5 = t_r6_c27_0 + p_5_26;
  assign t_r6_c27_6 = t_r6_c27_1 + p_5_28;
  assign t_r6_c27_7 = t_r6_c27_2 + t_r6_c27_3;
  assign t_r6_c27_8 = t_r6_c27_4 + p_7_26;
  assign t_r6_c27_9 = t_r6_c27_5 + t_r6_c27_6;
  assign t_r6_c27_10 = t_r6_c27_7 + t_r6_c27_8;
  assign t_r6_c27_11 = t_r6_c27_9 + t_r6_c27_10;
  assign t_r6_c27_12 = t_r6_c27_11 + p_7_28;
  assign out_6_27 = t_r6_c27_12 >> 4;

  assign t_r6_c28_0 = p_5_28 << 1;
  assign t_r6_c28_1 = p_6_27 << 1;
  assign t_r6_c28_2 = p_6_28 << 2;
  assign t_r6_c28_3 = p_6_29 << 1;
  assign t_r6_c28_4 = p_7_28 << 1;
  assign t_r6_c28_5 = t_r6_c28_0 + p_5_27;
  assign t_r6_c28_6 = t_r6_c28_1 + p_5_29;
  assign t_r6_c28_7 = t_r6_c28_2 + t_r6_c28_3;
  assign t_r6_c28_8 = t_r6_c28_4 + p_7_27;
  assign t_r6_c28_9 = t_r6_c28_5 + t_r6_c28_6;
  assign t_r6_c28_10 = t_r6_c28_7 + t_r6_c28_8;
  assign t_r6_c28_11 = t_r6_c28_9 + t_r6_c28_10;
  assign t_r6_c28_12 = t_r6_c28_11 + p_7_29;
  assign out_6_28 = t_r6_c28_12 >> 4;

  assign t_r6_c29_0 = p_5_29 << 1;
  assign t_r6_c29_1 = p_6_28 << 1;
  assign t_r6_c29_2 = p_6_29 << 2;
  assign t_r6_c29_3 = p_6_30 << 1;
  assign t_r6_c29_4 = p_7_29 << 1;
  assign t_r6_c29_5 = t_r6_c29_0 + p_5_28;
  assign t_r6_c29_6 = t_r6_c29_1 + p_5_30;
  assign t_r6_c29_7 = t_r6_c29_2 + t_r6_c29_3;
  assign t_r6_c29_8 = t_r6_c29_4 + p_7_28;
  assign t_r6_c29_9 = t_r6_c29_5 + t_r6_c29_6;
  assign t_r6_c29_10 = t_r6_c29_7 + t_r6_c29_8;
  assign t_r6_c29_11 = t_r6_c29_9 + t_r6_c29_10;
  assign t_r6_c29_12 = t_r6_c29_11 + p_7_30;
  assign out_6_29 = t_r6_c29_12 >> 4;

  assign t_r6_c30_0 = p_5_30 << 1;
  assign t_r6_c30_1 = p_6_29 << 1;
  assign t_r6_c30_2 = p_6_30 << 2;
  assign t_r6_c30_3 = p_6_31 << 1;
  assign t_r6_c30_4 = p_7_30 << 1;
  assign t_r6_c30_5 = t_r6_c30_0 + p_5_29;
  assign t_r6_c30_6 = t_r6_c30_1 + p_5_31;
  assign t_r6_c30_7 = t_r6_c30_2 + t_r6_c30_3;
  assign t_r6_c30_8 = t_r6_c30_4 + p_7_29;
  assign t_r6_c30_9 = t_r6_c30_5 + t_r6_c30_6;
  assign t_r6_c30_10 = t_r6_c30_7 + t_r6_c30_8;
  assign t_r6_c30_11 = t_r6_c30_9 + t_r6_c30_10;
  assign t_r6_c30_12 = t_r6_c30_11 + p_7_31;
  assign out_6_30 = t_r6_c30_12 >> 4;

  assign t_r6_c31_0 = p_5_31 << 1;
  assign t_r6_c31_1 = p_6_30 << 1;
  assign t_r6_c31_2 = p_6_31 << 2;
  assign t_r6_c31_3 = p_6_32 << 1;
  assign t_r6_c31_4 = p_7_31 << 1;
  assign t_r6_c31_5 = t_r6_c31_0 + p_5_30;
  assign t_r6_c31_6 = t_r6_c31_1 + p_5_32;
  assign t_r6_c31_7 = t_r6_c31_2 + t_r6_c31_3;
  assign t_r6_c31_8 = t_r6_c31_4 + p_7_30;
  assign t_r6_c31_9 = t_r6_c31_5 + t_r6_c31_6;
  assign t_r6_c31_10 = t_r6_c31_7 + t_r6_c31_8;
  assign t_r6_c31_11 = t_r6_c31_9 + t_r6_c31_10;
  assign t_r6_c31_12 = t_r6_c31_11 + p_7_32;
  assign out_6_31 = t_r6_c31_12 >> 4;

  assign t_r6_c32_0 = p_5_32 << 1;
  assign t_r6_c32_1 = p_6_31 << 1;
  assign t_r6_c32_2 = p_6_32 << 2;
  assign t_r6_c32_3 = p_6_33 << 1;
  assign t_r6_c32_4 = p_7_32 << 1;
  assign t_r6_c32_5 = t_r6_c32_0 + p_5_31;
  assign t_r6_c32_6 = t_r6_c32_1 + p_5_33;
  assign t_r6_c32_7 = t_r6_c32_2 + t_r6_c32_3;
  assign t_r6_c32_8 = t_r6_c32_4 + p_7_31;
  assign t_r6_c32_9 = t_r6_c32_5 + t_r6_c32_6;
  assign t_r6_c32_10 = t_r6_c32_7 + t_r6_c32_8;
  assign t_r6_c32_11 = t_r6_c32_9 + t_r6_c32_10;
  assign t_r6_c32_12 = t_r6_c32_11 + p_7_33;
  assign out_6_32 = t_r6_c32_12 >> 4;

  assign t_r6_c33_0 = p_5_33 << 1;
  assign t_r6_c33_1 = p_6_32 << 1;
  assign t_r6_c33_2 = p_6_33 << 2;
  assign t_r6_c33_3 = p_6_34 << 1;
  assign t_r6_c33_4 = p_7_33 << 1;
  assign t_r6_c33_5 = t_r6_c33_0 + p_5_32;
  assign t_r6_c33_6 = t_r6_c33_1 + p_5_34;
  assign t_r6_c33_7 = t_r6_c33_2 + t_r6_c33_3;
  assign t_r6_c33_8 = t_r6_c33_4 + p_7_32;
  assign t_r6_c33_9 = t_r6_c33_5 + t_r6_c33_6;
  assign t_r6_c33_10 = t_r6_c33_7 + t_r6_c33_8;
  assign t_r6_c33_11 = t_r6_c33_9 + t_r6_c33_10;
  assign t_r6_c33_12 = t_r6_c33_11 + p_7_34;
  assign out_6_33 = t_r6_c33_12 >> 4;

  assign t_r6_c34_0 = p_5_34 << 1;
  assign t_r6_c34_1 = p_6_33 << 1;
  assign t_r6_c34_2 = p_6_34 << 2;
  assign t_r6_c34_3 = p_6_35 << 1;
  assign t_r6_c34_4 = p_7_34 << 1;
  assign t_r6_c34_5 = t_r6_c34_0 + p_5_33;
  assign t_r6_c34_6 = t_r6_c34_1 + p_5_35;
  assign t_r6_c34_7 = t_r6_c34_2 + t_r6_c34_3;
  assign t_r6_c34_8 = t_r6_c34_4 + p_7_33;
  assign t_r6_c34_9 = t_r6_c34_5 + t_r6_c34_6;
  assign t_r6_c34_10 = t_r6_c34_7 + t_r6_c34_8;
  assign t_r6_c34_11 = t_r6_c34_9 + t_r6_c34_10;
  assign t_r6_c34_12 = t_r6_c34_11 + p_7_35;
  assign out_6_34 = t_r6_c34_12 >> 4;

  assign t_r6_c35_0 = p_5_35 << 1;
  assign t_r6_c35_1 = p_6_34 << 1;
  assign t_r6_c35_2 = p_6_35 << 2;
  assign t_r6_c35_3 = p_6_36 << 1;
  assign t_r6_c35_4 = p_7_35 << 1;
  assign t_r6_c35_5 = t_r6_c35_0 + p_5_34;
  assign t_r6_c35_6 = t_r6_c35_1 + p_5_36;
  assign t_r6_c35_7 = t_r6_c35_2 + t_r6_c35_3;
  assign t_r6_c35_8 = t_r6_c35_4 + p_7_34;
  assign t_r6_c35_9 = t_r6_c35_5 + t_r6_c35_6;
  assign t_r6_c35_10 = t_r6_c35_7 + t_r6_c35_8;
  assign t_r6_c35_11 = t_r6_c35_9 + t_r6_c35_10;
  assign t_r6_c35_12 = t_r6_c35_11 + p_7_36;
  assign out_6_35 = t_r6_c35_12 >> 4;

  assign t_r6_c36_0 = p_5_36 << 1;
  assign t_r6_c36_1 = p_6_35 << 1;
  assign t_r6_c36_2 = p_6_36 << 2;
  assign t_r6_c36_3 = p_6_37 << 1;
  assign t_r6_c36_4 = p_7_36 << 1;
  assign t_r6_c36_5 = t_r6_c36_0 + p_5_35;
  assign t_r6_c36_6 = t_r6_c36_1 + p_5_37;
  assign t_r6_c36_7 = t_r6_c36_2 + t_r6_c36_3;
  assign t_r6_c36_8 = t_r6_c36_4 + p_7_35;
  assign t_r6_c36_9 = t_r6_c36_5 + t_r6_c36_6;
  assign t_r6_c36_10 = t_r6_c36_7 + t_r6_c36_8;
  assign t_r6_c36_11 = t_r6_c36_9 + t_r6_c36_10;
  assign t_r6_c36_12 = t_r6_c36_11 + p_7_37;
  assign out_6_36 = t_r6_c36_12 >> 4;

  assign t_r6_c37_0 = p_5_37 << 1;
  assign t_r6_c37_1 = p_6_36 << 1;
  assign t_r6_c37_2 = p_6_37 << 2;
  assign t_r6_c37_3 = p_6_38 << 1;
  assign t_r6_c37_4 = p_7_37 << 1;
  assign t_r6_c37_5 = t_r6_c37_0 + p_5_36;
  assign t_r6_c37_6 = t_r6_c37_1 + p_5_38;
  assign t_r6_c37_7 = t_r6_c37_2 + t_r6_c37_3;
  assign t_r6_c37_8 = t_r6_c37_4 + p_7_36;
  assign t_r6_c37_9 = t_r6_c37_5 + t_r6_c37_6;
  assign t_r6_c37_10 = t_r6_c37_7 + t_r6_c37_8;
  assign t_r6_c37_11 = t_r6_c37_9 + t_r6_c37_10;
  assign t_r6_c37_12 = t_r6_c37_11 + p_7_38;
  assign out_6_37 = t_r6_c37_12 >> 4;

  assign t_r6_c38_0 = p_5_38 << 1;
  assign t_r6_c38_1 = p_6_37 << 1;
  assign t_r6_c38_2 = p_6_38 << 2;
  assign t_r6_c38_3 = p_6_39 << 1;
  assign t_r6_c38_4 = p_7_38 << 1;
  assign t_r6_c38_5 = t_r6_c38_0 + p_5_37;
  assign t_r6_c38_6 = t_r6_c38_1 + p_5_39;
  assign t_r6_c38_7 = t_r6_c38_2 + t_r6_c38_3;
  assign t_r6_c38_8 = t_r6_c38_4 + p_7_37;
  assign t_r6_c38_9 = t_r6_c38_5 + t_r6_c38_6;
  assign t_r6_c38_10 = t_r6_c38_7 + t_r6_c38_8;
  assign t_r6_c38_11 = t_r6_c38_9 + t_r6_c38_10;
  assign t_r6_c38_12 = t_r6_c38_11 + p_7_39;
  assign out_6_38 = t_r6_c38_12 >> 4;

  assign t_r6_c39_0 = p_5_39 << 1;
  assign t_r6_c39_1 = p_6_38 << 1;
  assign t_r6_c39_2 = p_6_39 << 2;
  assign t_r6_c39_3 = p_6_40 << 1;
  assign t_r6_c39_4 = p_7_39 << 1;
  assign t_r6_c39_5 = t_r6_c39_0 + p_5_38;
  assign t_r6_c39_6 = t_r6_c39_1 + p_5_40;
  assign t_r6_c39_7 = t_r6_c39_2 + t_r6_c39_3;
  assign t_r6_c39_8 = t_r6_c39_4 + p_7_38;
  assign t_r6_c39_9 = t_r6_c39_5 + t_r6_c39_6;
  assign t_r6_c39_10 = t_r6_c39_7 + t_r6_c39_8;
  assign t_r6_c39_11 = t_r6_c39_9 + t_r6_c39_10;
  assign t_r6_c39_12 = t_r6_c39_11 + p_7_40;
  assign out_6_39 = t_r6_c39_12 >> 4;

  assign t_r6_c40_0 = p_5_40 << 1;
  assign t_r6_c40_1 = p_6_39 << 1;
  assign t_r6_c40_2 = p_6_40 << 2;
  assign t_r6_c40_3 = p_6_41 << 1;
  assign t_r6_c40_4 = p_7_40 << 1;
  assign t_r6_c40_5 = t_r6_c40_0 + p_5_39;
  assign t_r6_c40_6 = t_r6_c40_1 + p_5_41;
  assign t_r6_c40_7 = t_r6_c40_2 + t_r6_c40_3;
  assign t_r6_c40_8 = t_r6_c40_4 + p_7_39;
  assign t_r6_c40_9 = t_r6_c40_5 + t_r6_c40_6;
  assign t_r6_c40_10 = t_r6_c40_7 + t_r6_c40_8;
  assign t_r6_c40_11 = t_r6_c40_9 + t_r6_c40_10;
  assign t_r6_c40_12 = t_r6_c40_11 + p_7_41;
  assign out_6_40 = t_r6_c40_12 >> 4;

  assign t_r6_c41_0 = p_5_41 << 1;
  assign t_r6_c41_1 = p_6_40 << 1;
  assign t_r6_c41_2 = p_6_41 << 2;
  assign t_r6_c41_3 = p_6_42 << 1;
  assign t_r6_c41_4 = p_7_41 << 1;
  assign t_r6_c41_5 = t_r6_c41_0 + p_5_40;
  assign t_r6_c41_6 = t_r6_c41_1 + p_5_42;
  assign t_r6_c41_7 = t_r6_c41_2 + t_r6_c41_3;
  assign t_r6_c41_8 = t_r6_c41_4 + p_7_40;
  assign t_r6_c41_9 = t_r6_c41_5 + t_r6_c41_6;
  assign t_r6_c41_10 = t_r6_c41_7 + t_r6_c41_8;
  assign t_r6_c41_11 = t_r6_c41_9 + t_r6_c41_10;
  assign t_r6_c41_12 = t_r6_c41_11 + p_7_42;
  assign out_6_41 = t_r6_c41_12 >> 4;

  assign t_r6_c42_0 = p_5_42 << 1;
  assign t_r6_c42_1 = p_6_41 << 1;
  assign t_r6_c42_2 = p_6_42 << 2;
  assign t_r6_c42_3 = p_6_43 << 1;
  assign t_r6_c42_4 = p_7_42 << 1;
  assign t_r6_c42_5 = t_r6_c42_0 + p_5_41;
  assign t_r6_c42_6 = t_r6_c42_1 + p_5_43;
  assign t_r6_c42_7 = t_r6_c42_2 + t_r6_c42_3;
  assign t_r6_c42_8 = t_r6_c42_4 + p_7_41;
  assign t_r6_c42_9 = t_r6_c42_5 + t_r6_c42_6;
  assign t_r6_c42_10 = t_r6_c42_7 + t_r6_c42_8;
  assign t_r6_c42_11 = t_r6_c42_9 + t_r6_c42_10;
  assign t_r6_c42_12 = t_r6_c42_11 + p_7_43;
  assign out_6_42 = t_r6_c42_12 >> 4;

  assign t_r6_c43_0 = p_5_43 << 1;
  assign t_r6_c43_1 = p_6_42 << 1;
  assign t_r6_c43_2 = p_6_43 << 2;
  assign t_r6_c43_3 = p_6_44 << 1;
  assign t_r6_c43_4 = p_7_43 << 1;
  assign t_r6_c43_5 = t_r6_c43_0 + p_5_42;
  assign t_r6_c43_6 = t_r6_c43_1 + p_5_44;
  assign t_r6_c43_7 = t_r6_c43_2 + t_r6_c43_3;
  assign t_r6_c43_8 = t_r6_c43_4 + p_7_42;
  assign t_r6_c43_9 = t_r6_c43_5 + t_r6_c43_6;
  assign t_r6_c43_10 = t_r6_c43_7 + t_r6_c43_8;
  assign t_r6_c43_11 = t_r6_c43_9 + t_r6_c43_10;
  assign t_r6_c43_12 = t_r6_c43_11 + p_7_44;
  assign out_6_43 = t_r6_c43_12 >> 4;

  assign t_r6_c44_0 = p_5_44 << 1;
  assign t_r6_c44_1 = p_6_43 << 1;
  assign t_r6_c44_2 = p_6_44 << 2;
  assign t_r6_c44_3 = p_6_45 << 1;
  assign t_r6_c44_4 = p_7_44 << 1;
  assign t_r6_c44_5 = t_r6_c44_0 + p_5_43;
  assign t_r6_c44_6 = t_r6_c44_1 + p_5_45;
  assign t_r6_c44_7 = t_r6_c44_2 + t_r6_c44_3;
  assign t_r6_c44_8 = t_r6_c44_4 + p_7_43;
  assign t_r6_c44_9 = t_r6_c44_5 + t_r6_c44_6;
  assign t_r6_c44_10 = t_r6_c44_7 + t_r6_c44_8;
  assign t_r6_c44_11 = t_r6_c44_9 + t_r6_c44_10;
  assign t_r6_c44_12 = t_r6_c44_11 + p_7_45;
  assign out_6_44 = t_r6_c44_12 >> 4;

  assign t_r6_c45_0 = p_5_45 << 1;
  assign t_r6_c45_1 = p_6_44 << 1;
  assign t_r6_c45_2 = p_6_45 << 2;
  assign t_r6_c45_3 = p_6_46 << 1;
  assign t_r6_c45_4 = p_7_45 << 1;
  assign t_r6_c45_5 = t_r6_c45_0 + p_5_44;
  assign t_r6_c45_6 = t_r6_c45_1 + p_5_46;
  assign t_r6_c45_7 = t_r6_c45_2 + t_r6_c45_3;
  assign t_r6_c45_8 = t_r6_c45_4 + p_7_44;
  assign t_r6_c45_9 = t_r6_c45_5 + t_r6_c45_6;
  assign t_r6_c45_10 = t_r6_c45_7 + t_r6_c45_8;
  assign t_r6_c45_11 = t_r6_c45_9 + t_r6_c45_10;
  assign t_r6_c45_12 = t_r6_c45_11 + p_7_46;
  assign out_6_45 = t_r6_c45_12 >> 4;

  assign t_r6_c46_0 = p_5_46 << 1;
  assign t_r6_c46_1 = p_6_45 << 1;
  assign t_r6_c46_2 = p_6_46 << 2;
  assign t_r6_c46_3 = p_6_47 << 1;
  assign t_r6_c46_4 = p_7_46 << 1;
  assign t_r6_c46_5 = t_r6_c46_0 + p_5_45;
  assign t_r6_c46_6 = t_r6_c46_1 + p_5_47;
  assign t_r6_c46_7 = t_r6_c46_2 + t_r6_c46_3;
  assign t_r6_c46_8 = t_r6_c46_4 + p_7_45;
  assign t_r6_c46_9 = t_r6_c46_5 + t_r6_c46_6;
  assign t_r6_c46_10 = t_r6_c46_7 + t_r6_c46_8;
  assign t_r6_c46_11 = t_r6_c46_9 + t_r6_c46_10;
  assign t_r6_c46_12 = t_r6_c46_11 + p_7_47;
  assign out_6_46 = t_r6_c46_12 >> 4;

  assign t_r6_c47_0 = p_5_47 << 1;
  assign t_r6_c47_1 = p_6_46 << 1;
  assign t_r6_c47_2 = p_6_47 << 2;
  assign t_r6_c47_3 = p_6_48 << 1;
  assign t_r6_c47_4 = p_7_47 << 1;
  assign t_r6_c47_5 = t_r6_c47_0 + p_5_46;
  assign t_r6_c47_6 = t_r6_c47_1 + p_5_48;
  assign t_r6_c47_7 = t_r6_c47_2 + t_r6_c47_3;
  assign t_r6_c47_8 = t_r6_c47_4 + p_7_46;
  assign t_r6_c47_9 = t_r6_c47_5 + t_r6_c47_6;
  assign t_r6_c47_10 = t_r6_c47_7 + t_r6_c47_8;
  assign t_r6_c47_11 = t_r6_c47_9 + t_r6_c47_10;
  assign t_r6_c47_12 = t_r6_c47_11 + p_7_48;
  assign out_6_47 = t_r6_c47_12 >> 4;

  assign t_r6_c48_0 = p_5_48 << 1;
  assign t_r6_c48_1 = p_6_47 << 1;
  assign t_r6_c48_2 = p_6_48 << 2;
  assign t_r6_c48_3 = p_6_49 << 1;
  assign t_r6_c48_4 = p_7_48 << 1;
  assign t_r6_c48_5 = t_r6_c48_0 + p_5_47;
  assign t_r6_c48_6 = t_r6_c48_1 + p_5_49;
  assign t_r6_c48_7 = t_r6_c48_2 + t_r6_c48_3;
  assign t_r6_c48_8 = t_r6_c48_4 + p_7_47;
  assign t_r6_c48_9 = t_r6_c48_5 + t_r6_c48_6;
  assign t_r6_c48_10 = t_r6_c48_7 + t_r6_c48_8;
  assign t_r6_c48_11 = t_r6_c48_9 + t_r6_c48_10;
  assign t_r6_c48_12 = t_r6_c48_11 + p_7_49;
  assign out_6_48 = t_r6_c48_12 >> 4;

  assign t_r6_c49_0 = p_5_49 << 1;
  assign t_r6_c49_1 = p_6_48 << 1;
  assign t_r6_c49_2 = p_6_49 << 2;
  assign t_r6_c49_3 = p_6_50 << 1;
  assign t_r6_c49_4 = p_7_49 << 1;
  assign t_r6_c49_5 = t_r6_c49_0 + p_5_48;
  assign t_r6_c49_6 = t_r6_c49_1 + p_5_50;
  assign t_r6_c49_7 = t_r6_c49_2 + t_r6_c49_3;
  assign t_r6_c49_8 = t_r6_c49_4 + p_7_48;
  assign t_r6_c49_9 = t_r6_c49_5 + t_r6_c49_6;
  assign t_r6_c49_10 = t_r6_c49_7 + t_r6_c49_8;
  assign t_r6_c49_11 = t_r6_c49_9 + t_r6_c49_10;
  assign t_r6_c49_12 = t_r6_c49_11 + p_7_50;
  assign out_6_49 = t_r6_c49_12 >> 4;

  assign t_r6_c50_0 = p_5_50 << 1;
  assign t_r6_c50_1 = p_6_49 << 1;
  assign t_r6_c50_2 = p_6_50 << 2;
  assign t_r6_c50_3 = p_6_51 << 1;
  assign t_r6_c50_4 = p_7_50 << 1;
  assign t_r6_c50_5 = t_r6_c50_0 + p_5_49;
  assign t_r6_c50_6 = t_r6_c50_1 + p_5_51;
  assign t_r6_c50_7 = t_r6_c50_2 + t_r6_c50_3;
  assign t_r6_c50_8 = t_r6_c50_4 + p_7_49;
  assign t_r6_c50_9 = t_r6_c50_5 + t_r6_c50_6;
  assign t_r6_c50_10 = t_r6_c50_7 + t_r6_c50_8;
  assign t_r6_c50_11 = t_r6_c50_9 + t_r6_c50_10;
  assign t_r6_c50_12 = t_r6_c50_11 + p_7_51;
  assign out_6_50 = t_r6_c50_12 >> 4;

  assign t_r6_c51_0 = p_5_51 << 1;
  assign t_r6_c51_1 = p_6_50 << 1;
  assign t_r6_c51_2 = p_6_51 << 2;
  assign t_r6_c51_3 = p_6_52 << 1;
  assign t_r6_c51_4 = p_7_51 << 1;
  assign t_r6_c51_5 = t_r6_c51_0 + p_5_50;
  assign t_r6_c51_6 = t_r6_c51_1 + p_5_52;
  assign t_r6_c51_7 = t_r6_c51_2 + t_r6_c51_3;
  assign t_r6_c51_8 = t_r6_c51_4 + p_7_50;
  assign t_r6_c51_9 = t_r6_c51_5 + t_r6_c51_6;
  assign t_r6_c51_10 = t_r6_c51_7 + t_r6_c51_8;
  assign t_r6_c51_11 = t_r6_c51_9 + t_r6_c51_10;
  assign t_r6_c51_12 = t_r6_c51_11 + p_7_52;
  assign out_6_51 = t_r6_c51_12 >> 4;

  assign t_r6_c52_0 = p_5_52 << 1;
  assign t_r6_c52_1 = p_6_51 << 1;
  assign t_r6_c52_2 = p_6_52 << 2;
  assign t_r6_c52_3 = p_6_53 << 1;
  assign t_r6_c52_4 = p_7_52 << 1;
  assign t_r6_c52_5 = t_r6_c52_0 + p_5_51;
  assign t_r6_c52_6 = t_r6_c52_1 + p_5_53;
  assign t_r6_c52_7 = t_r6_c52_2 + t_r6_c52_3;
  assign t_r6_c52_8 = t_r6_c52_4 + p_7_51;
  assign t_r6_c52_9 = t_r6_c52_5 + t_r6_c52_6;
  assign t_r6_c52_10 = t_r6_c52_7 + t_r6_c52_8;
  assign t_r6_c52_11 = t_r6_c52_9 + t_r6_c52_10;
  assign t_r6_c52_12 = t_r6_c52_11 + p_7_53;
  assign out_6_52 = t_r6_c52_12 >> 4;

  assign t_r6_c53_0 = p_5_53 << 1;
  assign t_r6_c53_1 = p_6_52 << 1;
  assign t_r6_c53_2 = p_6_53 << 2;
  assign t_r6_c53_3 = p_6_54 << 1;
  assign t_r6_c53_4 = p_7_53 << 1;
  assign t_r6_c53_5 = t_r6_c53_0 + p_5_52;
  assign t_r6_c53_6 = t_r6_c53_1 + p_5_54;
  assign t_r6_c53_7 = t_r6_c53_2 + t_r6_c53_3;
  assign t_r6_c53_8 = t_r6_c53_4 + p_7_52;
  assign t_r6_c53_9 = t_r6_c53_5 + t_r6_c53_6;
  assign t_r6_c53_10 = t_r6_c53_7 + t_r6_c53_8;
  assign t_r6_c53_11 = t_r6_c53_9 + t_r6_c53_10;
  assign t_r6_c53_12 = t_r6_c53_11 + p_7_54;
  assign out_6_53 = t_r6_c53_12 >> 4;

  assign t_r6_c54_0 = p_5_54 << 1;
  assign t_r6_c54_1 = p_6_53 << 1;
  assign t_r6_c54_2 = p_6_54 << 2;
  assign t_r6_c54_3 = p_6_55 << 1;
  assign t_r6_c54_4 = p_7_54 << 1;
  assign t_r6_c54_5 = t_r6_c54_0 + p_5_53;
  assign t_r6_c54_6 = t_r6_c54_1 + p_5_55;
  assign t_r6_c54_7 = t_r6_c54_2 + t_r6_c54_3;
  assign t_r6_c54_8 = t_r6_c54_4 + p_7_53;
  assign t_r6_c54_9 = t_r6_c54_5 + t_r6_c54_6;
  assign t_r6_c54_10 = t_r6_c54_7 + t_r6_c54_8;
  assign t_r6_c54_11 = t_r6_c54_9 + t_r6_c54_10;
  assign t_r6_c54_12 = t_r6_c54_11 + p_7_55;
  assign out_6_54 = t_r6_c54_12 >> 4;

  assign t_r6_c55_0 = p_5_55 << 1;
  assign t_r6_c55_1 = p_6_54 << 1;
  assign t_r6_c55_2 = p_6_55 << 2;
  assign t_r6_c55_3 = p_6_56 << 1;
  assign t_r6_c55_4 = p_7_55 << 1;
  assign t_r6_c55_5 = t_r6_c55_0 + p_5_54;
  assign t_r6_c55_6 = t_r6_c55_1 + p_5_56;
  assign t_r6_c55_7 = t_r6_c55_2 + t_r6_c55_3;
  assign t_r6_c55_8 = t_r6_c55_4 + p_7_54;
  assign t_r6_c55_9 = t_r6_c55_5 + t_r6_c55_6;
  assign t_r6_c55_10 = t_r6_c55_7 + t_r6_c55_8;
  assign t_r6_c55_11 = t_r6_c55_9 + t_r6_c55_10;
  assign t_r6_c55_12 = t_r6_c55_11 + p_7_56;
  assign out_6_55 = t_r6_c55_12 >> 4;

  assign t_r6_c56_0 = p_5_56 << 1;
  assign t_r6_c56_1 = p_6_55 << 1;
  assign t_r6_c56_2 = p_6_56 << 2;
  assign t_r6_c56_3 = p_6_57 << 1;
  assign t_r6_c56_4 = p_7_56 << 1;
  assign t_r6_c56_5 = t_r6_c56_0 + p_5_55;
  assign t_r6_c56_6 = t_r6_c56_1 + p_5_57;
  assign t_r6_c56_7 = t_r6_c56_2 + t_r6_c56_3;
  assign t_r6_c56_8 = t_r6_c56_4 + p_7_55;
  assign t_r6_c56_9 = t_r6_c56_5 + t_r6_c56_6;
  assign t_r6_c56_10 = t_r6_c56_7 + t_r6_c56_8;
  assign t_r6_c56_11 = t_r6_c56_9 + t_r6_c56_10;
  assign t_r6_c56_12 = t_r6_c56_11 + p_7_57;
  assign out_6_56 = t_r6_c56_12 >> 4;

  assign t_r6_c57_0 = p_5_57 << 1;
  assign t_r6_c57_1 = p_6_56 << 1;
  assign t_r6_c57_2 = p_6_57 << 2;
  assign t_r6_c57_3 = p_6_58 << 1;
  assign t_r6_c57_4 = p_7_57 << 1;
  assign t_r6_c57_5 = t_r6_c57_0 + p_5_56;
  assign t_r6_c57_6 = t_r6_c57_1 + p_5_58;
  assign t_r6_c57_7 = t_r6_c57_2 + t_r6_c57_3;
  assign t_r6_c57_8 = t_r6_c57_4 + p_7_56;
  assign t_r6_c57_9 = t_r6_c57_5 + t_r6_c57_6;
  assign t_r6_c57_10 = t_r6_c57_7 + t_r6_c57_8;
  assign t_r6_c57_11 = t_r6_c57_9 + t_r6_c57_10;
  assign t_r6_c57_12 = t_r6_c57_11 + p_7_58;
  assign out_6_57 = t_r6_c57_12 >> 4;

  assign t_r6_c58_0 = p_5_58 << 1;
  assign t_r6_c58_1 = p_6_57 << 1;
  assign t_r6_c58_2 = p_6_58 << 2;
  assign t_r6_c58_3 = p_6_59 << 1;
  assign t_r6_c58_4 = p_7_58 << 1;
  assign t_r6_c58_5 = t_r6_c58_0 + p_5_57;
  assign t_r6_c58_6 = t_r6_c58_1 + p_5_59;
  assign t_r6_c58_7 = t_r6_c58_2 + t_r6_c58_3;
  assign t_r6_c58_8 = t_r6_c58_4 + p_7_57;
  assign t_r6_c58_9 = t_r6_c58_5 + t_r6_c58_6;
  assign t_r6_c58_10 = t_r6_c58_7 + t_r6_c58_8;
  assign t_r6_c58_11 = t_r6_c58_9 + t_r6_c58_10;
  assign t_r6_c58_12 = t_r6_c58_11 + p_7_59;
  assign out_6_58 = t_r6_c58_12 >> 4;

  assign t_r6_c59_0 = p_5_59 << 1;
  assign t_r6_c59_1 = p_6_58 << 1;
  assign t_r6_c59_2 = p_6_59 << 2;
  assign t_r6_c59_3 = p_6_60 << 1;
  assign t_r6_c59_4 = p_7_59 << 1;
  assign t_r6_c59_5 = t_r6_c59_0 + p_5_58;
  assign t_r6_c59_6 = t_r6_c59_1 + p_5_60;
  assign t_r6_c59_7 = t_r6_c59_2 + t_r6_c59_3;
  assign t_r6_c59_8 = t_r6_c59_4 + p_7_58;
  assign t_r6_c59_9 = t_r6_c59_5 + t_r6_c59_6;
  assign t_r6_c59_10 = t_r6_c59_7 + t_r6_c59_8;
  assign t_r6_c59_11 = t_r6_c59_9 + t_r6_c59_10;
  assign t_r6_c59_12 = t_r6_c59_11 + p_7_60;
  assign out_6_59 = t_r6_c59_12 >> 4;

  assign t_r6_c60_0 = p_5_60 << 1;
  assign t_r6_c60_1 = p_6_59 << 1;
  assign t_r6_c60_2 = p_6_60 << 2;
  assign t_r6_c60_3 = p_6_61 << 1;
  assign t_r6_c60_4 = p_7_60 << 1;
  assign t_r6_c60_5 = t_r6_c60_0 + p_5_59;
  assign t_r6_c60_6 = t_r6_c60_1 + p_5_61;
  assign t_r6_c60_7 = t_r6_c60_2 + t_r6_c60_3;
  assign t_r6_c60_8 = t_r6_c60_4 + p_7_59;
  assign t_r6_c60_9 = t_r6_c60_5 + t_r6_c60_6;
  assign t_r6_c60_10 = t_r6_c60_7 + t_r6_c60_8;
  assign t_r6_c60_11 = t_r6_c60_9 + t_r6_c60_10;
  assign t_r6_c60_12 = t_r6_c60_11 + p_7_61;
  assign out_6_60 = t_r6_c60_12 >> 4;

  assign t_r6_c61_0 = p_5_61 << 1;
  assign t_r6_c61_1 = p_6_60 << 1;
  assign t_r6_c61_2 = p_6_61 << 2;
  assign t_r6_c61_3 = p_6_62 << 1;
  assign t_r6_c61_4 = p_7_61 << 1;
  assign t_r6_c61_5 = t_r6_c61_0 + p_5_60;
  assign t_r6_c61_6 = t_r6_c61_1 + p_5_62;
  assign t_r6_c61_7 = t_r6_c61_2 + t_r6_c61_3;
  assign t_r6_c61_8 = t_r6_c61_4 + p_7_60;
  assign t_r6_c61_9 = t_r6_c61_5 + t_r6_c61_6;
  assign t_r6_c61_10 = t_r6_c61_7 + t_r6_c61_8;
  assign t_r6_c61_11 = t_r6_c61_9 + t_r6_c61_10;
  assign t_r6_c61_12 = t_r6_c61_11 + p_7_62;
  assign out_6_61 = t_r6_c61_12 >> 4;

  assign t_r6_c62_0 = p_5_62 << 1;
  assign t_r6_c62_1 = p_6_61 << 1;
  assign t_r6_c62_2 = p_6_62 << 2;
  assign t_r6_c62_3 = p_6_63 << 1;
  assign t_r6_c62_4 = p_7_62 << 1;
  assign t_r6_c62_5 = t_r6_c62_0 + p_5_61;
  assign t_r6_c62_6 = t_r6_c62_1 + p_5_63;
  assign t_r6_c62_7 = t_r6_c62_2 + t_r6_c62_3;
  assign t_r6_c62_8 = t_r6_c62_4 + p_7_61;
  assign t_r6_c62_9 = t_r6_c62_5 + t_r6_c62_6;
  assign t_r6_c62_10 = t_r6_c62_7 + t_r6_c62_8;
  assign t_r6_c62_11 = t_r6_c62_9 + t_r6_c62_10;
  assign t_r6_c62_12 = t_r6_c62_11 + p_7_63;
  assign out_6_62 = t_r6_c62_12 >> 4;

  assign t_r6_c63_0 = p_5_63 << 1;
  assign t_r6_c63_1 = p_6_62 << 1;
  assign t_r6_c63_2 = p_6_63 << 2;
  assign t_r6_c63_3 = p_6_64 << 1;
  assign t_r6_c63_4 = p_7_63 << 1;
  assign t_r6_c63_5 = t_r6_c63_0 + p_5_62;
  assign t_r6_c63_6 = t_r6_c63_1 + p_5_64;
  assign t_r6_c63_7 = t_r6_c63_2 + t_r6_c63_3;
  assign t_r6_c63_8 = t_r6_c63_4 + p_7_62;
  assign t_r6_c63_9 = t_r6_c63_5 + t_r6_c63_6;
  assign t_r6_c63_10 = t_r6_c63_7 + t_r6_c63_8;
  assign t_r6_c63_11 = t_r6_c63_9 + t_r6_c63_10;
  assign t_r6_c63_12 = t_r6_c63_11 + p_7_64;
  assign out_6_63 = t_r6_c63_12 >> 4;

  assign t_r6_c64_0 = p_5_64 << 1;
  assign t_r6_c64_1 = p_6_63 << 1;
  assign t_r6_c64_2 = p_6_64 << 2;
  assign t_r6_c64_3 = p_6_65 << 1;
  assign t_r6_c64_4 = p_7_64 << 1;
  assign t_r6_c64_5 = t_r6_c64_0 + p_5_63;
  assign t_r6_c64_6 = t_r6_c64_1 + p_5_65;
  assign t_r6_c64_7 = t_r6_c64_2 + t_r6_c64_3;
  assign t_r6_c64_8 = t_r6_c64_4 + p_7_63;
  assign t_r6_c64_9 = t_r6_c64_5 + t_r6_c64_6;
  assign t_r6_c64_10 = t_r6_c64_7 + t_r6_c64_8;
  assign t_r6_c64_11 = t_r6_c64_9 + t_r6_c64_10;
  assign t_r6_c64_12 = t_r6_c64_11 + p_7_65;
  assign out_6_64 = t_r6_c64_12 >> 4;

  assign t_r7_c1_0 = p_6_1 << 1;
  assign t_r7_c1_1 = p_7_0 << 1;
  assign t_r7_c1_2 = p_7_1 << 2;
  assign t_r7_c1_3 = p_7_2 << 1;
  assign t_r7_c1_4 = p_8_1 << 1;
  assign t_r7_c1_5 = t_r7_c1_0 + p_6_0;
  assign t_r7_c1_6 = t_r7_c1_1 + p_6_2;
  assign t_r7_c1_7 = t_r7_c1_2 + t_r7_c1_3;
  assign t_r7_c1_8 = t_r7_c1_4 + p_8_0;
  assign t_r7_c1_9 = t_r7_c1_5 + t_r7_c1_6;
  assign t_r7_c1_10 = t_r7_c1_7 + t_r7_c1_8;
  assign t_r7_c1_11 = t_r7_c1_9 + t_r7_c1_10;
  assign t_r7_c1_12 = t_r7_c1_11 + p_8_2;
  assign out_7_1 = t_r7_c1_12 >> 4;

  assign t_r7_c2_0 = p_6_2 << 1;
  assign t_r7_c2_1 = p_7_1 << 1;
  assign t_r7_c2_2 = p_7_2 << 2;
  assign t_r7_c2_3 = p_7_3 << 1;
  assign t_r7_c2_4 = p_8_2 << 1;
  assign t_r7_c2_5 = t_r7_c2_0 + p_6_1;
  assign t_r7_c2_6 = t_r7_c2_1 + p_6_3;
  assign t_r7_c2_7 = t_r7_c2_2 + t_r7_c2_3;
  assign t_r7_c2_8 = t_r7_c2_4 + p_8_1;
  assign t_r7_c2_9 = t_r7_c2_5 + t_r7_c2_6;
  assign t_r7_c2_10 = t_r7_c2_7 + t_r7_c2_8;
  assign t_r7_c2_11 = t_r7_c2_9 + t_r7_c2_10;
  assign t_r7_c2_12 = t_r7_c2_11 + p_8_3;
  assign out_7_2 = t_r7_c2_12 >> 4;

  assign t_r7_c3_0 = p_6_3 << 1;
  assign t_r7_c3_1 = p_7_2 << 1;
  assign t_r7_c3_2 = p_7_3 << 2;
  assign t_r7_c3_3 = p_7_4 << 1;
  assign t_r7_c3_4 = p_8_3 << 1;
  assign t_r7_c3_5 = t_r7_c3_0 + p_6_2;
  assign t_r7_c3_6 = t_r7_c3_1 + p_6_4;
  assign t_r7_c3_7 = t_r7_c3_2 + t_r7_c3_3;
  assign t_r7_c3_8 = t_r7_c3_4 + p_8_2;
  assign t_r7_c3_9 = t_r7_c3_5 + t_r7_c3_6;
  assign t_r7_c3_10 = t_r7_c3_7 + t_r7_c3_8;
  assign t_r7_c3_11 = t_r7_c3_9 + t_r7_c3_10;
  assign t_r7_c3_12 = t_r7_c3_11 + p_8_4;
  assign out_7_3 = t_r7_c3_12 >> 4;

  assign t_r7_c4_0 = p_6_4 << 1;
  assign t_r7_c4_1 = p_7_3 << 1;
  assign t_r7_c4_2 = p_7_4 << 2;
  assign t_r7_c4_3 = p_7_5 << 1;
  assign t_r7_c4_4 = p_8_4 << 1;
  assign t_r7_c4_5 = t_r7_c4_0 + p_6_3;
  assign t_r7_c4_6 = t_r7_c4_1 + p_6_5;
  assign t_r7_c4_7 = t_r7_c4_2 + t_r7_c4_3;
  assign t_r7_c4_8 = t_r7_c4_4 + p_8_3;
  assign t_r7_c4_9 = t_r7_c4_5 + t_r7_c4_6;
  assign t_r7_c4_10 = t_r7_c4_7 + t_r7_c4_8;
  assign t_r7_c4_11 = t_r7_c4_9 + t_r7_c4_10;
  assign t_r7_c4_12 = t_r7_c4_11 + p_8_5;
  assign out_7_4 = t_r7_c4_12 >> 4;

  assign t_r7_c5_0 = p_6_5 << 1;
  assign t_r7_c5_1 = p_7_4 << 1;
  assign t_r7_c5_2 = p_7_5 << 2;
  assign t_r7_c5_3 = p_7_6 << 1;
  assign t_r7_c5_4 = p_8_5 << 1;
  assign t_r7_c5_5 = t_r7_c5_0 + p_6_4;
  assign t_r7_c5_6 = t_r7_c5_1 + p_6_6;
  assign t_r7_c5_7 = t_r7_c5_2 + t_r7_c5_3;
  assign t_r7_c5_8 = t_r7_c5_4 + p_8_4;
  assign t_r7_c5_9 = t_r7_c5_5 + t_r7_c5_6;
  assign t_r7_c5_10 = t_r7_c5_7 + t_r7_c5_8;
  assign t_r7_c5_11 = t_r7_c5_9 + t_r7_c5_10;
  assign t_r7_c5_12 = t_r7_c5_11 + p_8_6;
  assign out_7_5 = t_r7_c5_12 >> 4;

  assign t_r7_c6_0 = p_6_6 << 1;
  assign t_r7_c6_1 = p_7_5 << 1;
  assign t_r7_c6_2 = p_7_6 << 2;
  assign t_r7_c6_3 = p_7_7 << 1;
  assign t_r7_c6_4 = p_8_6 << 1;
  assign t_r7_c6_5 = t_r7_c6_0 + p_6_5;
  assign t_r7_c6_6 = t_r7_c6_1 + p_6_7;
  assign t_r7_c6_7 = t_r7_c6_2 + t_r7_c6_3;
  assign t_r7_c6_8 = t_r7_c6_4 + p_8_5;
  assign t_r7_c6_9 = t_r7_c6_5 + t_r7_c6_6;
  assign t_r7_c6_10 = t_r7_c6_7 + t_r7_c6_8;
  assign t_r7_c6_11 = t_r7_c6_9 + t_r7_c6_10;
  assign t_r7_c6_12 = t_r7_c6_11 + p_8_7;
  assign out_7_6 = t_r7_c6_12 >> 4;

  assign t_r7_c7_0 = p_6_7 << 1;
  assign t_r7_c7_1 = p_7_6 << 1;
  assign t_r7_c7_2 = p_7_7 << 2;
  assign t_r7_c7_3 = p_7_8 << 1;
  assign t_r7_c7_4 = p_8_7 << 1;
  assign t_r7_c7_5 = t_r7_c7_0 + p_6_6;
  assign t_r7_c7_6 = t_r7_c7_1 + p_6_8;
  assign t_r7_c7_7 = t_r7_c7_2 + t_r7_c7_3;
  assign t_r7_c7_8 = t_r7_c7_4 + p_8_6;
  assign t_r7_c7_9 = t_r7_c7_5 + t_r7_c7_6;
  assign t_r7_c7_10 = t_r7_c7_7 + t_r7_c7_8;
  assign t_r7_c7_11 = t_r7_c7_9 + t_r7_c7_10;
  assign t_r7_c7_12 = t_r7_c7_11 + p_8_8;
  assign out_7_7 = t_r7_c7_12 >> 4;

  assign t_r7_c8_0 = p_6_8 << 1;
  assign t_r7_c8_1 = p_7_7 << 1;
  assign t_r7_c8_2 = p_7_8 << 2;
  assign t_r7_c8_3 = p_7_9 << 1;
  assign t_r7_c8_4 = p_8_8 << 1;
  assign t_r7_c8_5 = t_r7_c8_0 + p_6_7;
  assign t_r7_c8_6 = t_r7_c8_1 + p_6_9;
  assign t_r7_c8_7 = t_r7_c8_2 + t_r7_c8_3;
  assign t_r7_c8_8 = t_r7_c8_4 + p_8_7;
  assign t_r7_c8_9 = t_r7_c8_5 + t_r7_c8_6;
  assign t_r7_c8_10 = t_r7_c8_7 + t_r7_c8_8;
  assign t_r7_c8_11 = t_r7_c8_9 + t_r7_c8_10;
  assign t_r7_c8_12 = t_r7_c8_11 + p_8_9;
  assign out_7_8 = t_r7_c8_12 >> 4;

  assign t_r7_c9_0 = p_6_9 << 1;
  assign t_r7_c9_1 = p_7_8 << 1;
  assign t_r7_c9_2 = p_7_9 << 2;
  assign t_r7_c9_3 = p_7_10 << 1;
  assign t_r7_c9_4 = p_8_9 << 1;
  assign t_r7_c9_5 = t_r7_c9_0 + p_6_8;
  assign t_r7_c9_6 = t_r7_c9_1 + p_6_10;
  assign t_r7_c9_7 = t_r7_c9_2 + t_r7_c9_3;
  assign t_r7_c9_8 = t_r7_c9_4 + p_8_8;
  assign t_r7_c9_9 = t_r7_c9_5 + t_r7_c9_6;
  assign t_r7_c9_10 = t_r7_c9_7 + t_r7_c9_8;
  assign t_r7_c9_11 = t_r7_c9_9 + t_r7_c9_10;
  assign t_r7_c9_12 = t_r7_c9_11 + p_8_10;
  assign out_7_9 = t_r7_c9_12 >> 4;

  assign t_r7_c10_0 = p_6_10 << 1;
  assign t_r7_c10_1 = p_7_9 << 1;
  assign t_r7_c10_2 = p_7_10 << 2;
  assign t_r7_c10_3 = p_7_11 << 1;
  assign t_r7_c10_4 = p_8_10 << 1;
  assign t_r7_c10_5 = t_r7_c10_0 + p_6_9;
  assign t_r7_c10_6 = t_r7_c10_1 + p_6_11;
  assign t_r7_c10_7 = t_r7_c10_2 + t_r7_c10_3;
  assign t_r7_c10_8 = t_r7_c10_4 + p_8_9;
  assign t_r7_c10_9 = t_r7_c10_5 + t_r7_c10_6;
  assign t_r7_c10_10 = t_r7_c10_7 + t_r7_c10_8;
  assign t_r7_c10_11 = t_r7_c10_9 + t_r7_c10_10;
  assign t_r7_c10_12 = t_r7_c10_11 + p_8_11;
  assign out_7_10 = t_r7_c10_12 >> 4;

  assign t_r7_c11_0 = p_6_11 << 1;
  assign t_r7_c11_1 = p_7_10 << 1;
  assign t_r7_c11_2 = p_7_11 << 2;
  assign t_r7_c11_3 = p_7_12 << 1;
  assign t_r7_c11_4 = p_8_11 << 1;
  assign t_r7_c11_5 = t_r7_c11_0 + p_6_10;
  assign t_r7_c11_6 = t_r7_c11_1 + p_6_12;
  assign t_r7_c11_7 = t_r7_c11_2 + t_r7_c11_3;
  assign t_r7_c11_8 = t_r7_c11_4 + p_8_10;
  assign t_r7_c11_9 = t_r7_c11_5 + t_r7_c11_6;
  assign t_r7_c11_10 = t_r7_c11_7 + t_r7_c11_8;
  assign t_r7_c11_11 = t_r7_c11_9 + t_r7_c11_10;
  assign t_r7_c11_12 = t_r7_c11_11 + p_8_12;
  assign out_7_11 = t_r7_c11_12 >> 4;

  assign t_r7_c12_0 = p_6_12 << 1;
  assign t_r7_c12_1 = p_7_11 << 1;
  assign t_r7_c12_2 = p_7_12 << 2;
  assign t_r7_c12_3 = p_7_13 << 1;
  assign t_r7_c12_4 = p_8_12 << 1;
  assign t_r7_c12_5 = t_r7_c12_0 + p_6_11;
  assign t_r7_c12_6 = t_r7_c12_1 + p_6_13;
  assign t_r7_c12_7 = t_r7_c12_2 + t_r7_c12_3;
  assign t_r7_c12_8 = t_r7_c12_4 + p_8_11;
  assign t_r7_c12_9 = t_r7_c12_5 + t_r7_c12_6;
  assign t_r7_c12_10 = t_r7_c12_7 + t_r7_c12_8;
  assign t_r7_c12_11 = t_r7_c12_9 + t_r7_c12_10;
  assign t_r7_c12_12 = t_r7_c12_11 + p_8_13;
  assign out_7_12 = t_r7_c12_12 >> 4;

  assign t_r7_c13_0 = p_6_13 << 1;
  assign t_r7_c13_1 = p_7_12 << 1;
  assign t_r7_c13_2 = p_7_13 << 2;
  assign t_r7_c13_3 = p_7_14 << 1;
  assign t_r7_c13_4 = p_8_13 << 1;
  assign t_r7_c13_5 = t_r7_c13_0 + p_6_12;
  assign t_r7_c13_6 = t_r7_c13_1 + p_6_14;
  assign t_r7_c13_7 = t_r7_c13_2 + t_r7_c13_3;
  assign t_r7_c13_8 = t_r7_c13_4 + p_8_12;
  assign t_r7_c13_9 = t_r7_c13_5 + t_r7_c13_6;
  assign t_r7_c13_10 = t_r7_c13_7 + t_r7_c13_8;
  assign t_r7_c13_11 = t_r7_c13_9 + t_r7_c13_10;
  assign t_r7_c13_12 = t_r7_c13_11 + p_8_14;
  assign out_7_13 = t_r7_c13_12 >> 4;

  assign t_r7_c14_0 = p_6_14 << 1;
  assign t_r7_c14_1 = p_7_13 << 1;
  assign t_r7_c14_2 = p_7_14 << 2;
  assign t_r7_c14_3 = p_7_15 << 1;
  assign t_r7_c14_4 = p_8_14 << 1;
  assign t_r7_c14_5 = t_r7_c14_0 + p_6_13;
  assign t_r7_c14_6 = t_r7_c14_1 + p_6_15;
  assign t_r7_c14_7 = t_r7_c14_2 + t_r7_c14_3;
  assign t_r7_c14_8 = t_r7_c14_4 + p_8_13;
  assign t_r7_c14_9 = t_r7_c14_5 + t_r7_c14_6;
  assign t_r7_c14_10 = t_r7_c14_7 + t_r7_c14_8;
  assign t_r7_c14_11 = t_r7_c14_9 + t_r7_c14_10;
  assign t_r7_c14_12 = t_r7_c14_11 + p_8_15;
  assign out_7_14 = t_r7_c14_12 >> 4;

  assign t_r7_c15_0 = p_6_15 << 1;
  assign t_r7_c15_1 = p_7_14 << 1;
  assign t_r7_c15_2 = p_7_15 << 2;
  assign t_r7_c15_3 = p_7_16 << 1;
  assign t_r7_c15_4 = p_8_15 << 1;
  assign t_r7_c15_5 = t_r7_c15_0 + p_6_14;
  assign t_r7_c15_6 = t_r7_c15_1 + p_6_16;
  assign t_r7_c15_7 = t_r7_c15_2 + t_r7_c15_3;
  assign t_r7_c15_8 = t_r7_c15_4 + p_8_14;
  assign t_r7_c15_9 = t_r7_c15_5 + t_r7_c15_6;
  assign t_r7_c15_10 = t_r7_c15_7 + t_r7_c15_8;
  assign t_r7_c15_11 = t_r7_c15_9 + t_r7_c15_10;
  assign t_r7_c15_12 = t_r7_c15_11 + p_8_16;
  assign out_7_15 = t_r7_c15_12 >> 4;

  assign t_r7_c16_0 = p_6_16 << 1;
  assign t_r7_c16_1 = p_7_15 << 1;
  assign t_r7_c16_2 = p_7_16 << 2;
  assign t_r7_c16_3 = p_7_17 << 1;
  assign t_r7_c16_4 = p_8_16 << 1;
  assign t_r7_c16_5 = t_r7_c16_0 + p_6_15;
  assign t_r7_c16_6 = t_r7_c16_1 + p_6_17;
  assign t_r7_c16_7 = t_r7_c16_2 + t_r7_c16_3;
  assign t_r7_c16_8 = t_r7_c16_4 + p_8_15;
  assign t_r7_c16_9 = t_r7_c16_5 + t_r7_c16_6;
  assign t_r7_c16_10 = t_r7_c16_7 + t_r7_c16_8;
  assign t_r7_c16_11 = t_r7_c16_9 + t_r7_c16_10;
  assign t_r7_c16_12 = t_r7_c16_11 + p_8_17;
  assign out_7_16 = t_r7_c16_12 >> 4;

  assign t_r7_c17_0 = p_6_17 << 1;
  assign t_r7_c17_1 = p_7_16 << 1;
  assign t_r7_c17_2 = p_7_17 << 2;
  assign t_r7_c17_3 = p_7_18 << 1;
  assign t_r7_c17_4 = p_8_17 << 1;
  assign t_r7_c17_5 = t_r7_c17_0 + p_6_16;
  assign t_r7_c17_6 = t_r7_c17_1 + p_6_18;
  assign t_r7_c17_7 = t_r7_c17_2 + t_r7_c17_3;
  assign t_r7_c17_8 = t_r7_c17_4 + p_8_16;
  assign t_r7_c17_9 = t_r7_c17_5 + t_r7_c17_6;
  assign t_r7_c17_10 = t_r7_c17_7 + t_r7_c17_8;
  assign t_r7_c17_11 = t_r7_c17_9 + t_r7_c17_10;
  assign t_r7_c17_12 = t_r7_c17_11 + p_8_18;
  assign out_7_17 = t_r7_c17_12 >> 4;

  assign t_r7_c18_0 = p_6_18 << 1;
  assign t_r7_c18_1 = p_7_17 << 1;
  assign t_r7_c18_2 = p_7_18 << 2;
  assign t_r7_c18_3 = p_7_19 << 1;
  assign t_r7_c18_4 = p_8_18 << 1;
  assign t_r7_c18_5 = t_r7_c18_0 + p_6_17;
  assign t_r7_c18_6 = t_r7_c18_1 + p_6_19;
  assign t_r7_c18_7 = t_r7_c18_2 + t_r7_c18_3;
  assign t_r7_c18_8 = t_r7_c18_4 + p_8_17;
  assign t_r7_c18_9 = t_r7_c18_5 + t_r7_c18_6;
  assign t_r7_c18_10 = t_r7_c18_7 + t_r7_c18_8;
  assign t_r7_c18_11 = t_r7_c18_9 + t_r7_c18_10;
  assign t_r7_c18_12 = t_r7_c18_11 + p_8_19;
  assign out_7_18 = t_r7_c18_12 >> 4;

  assign t_r7_c19_0 = p_6_19 << 1;
  assign t_r7_c19_1 = p_7_18 << 1;
  assign t_r7_c19_2 = p_7_19 << 2;
  assign t_r7_c19_3 = p_7_20 << 1;
  assign t_r7_c19_4 = p_8_19 << 1;
  assign t_r7_c19_5 = t_r7_c19_0 + p_6_18;
  assign t_r7_c19_6 = t_r7_c19_1 + p_6_20;
  assign t_r7_c19_7 = t_r7_c19_2 + t_r7_c19_3;
  assign t_r7_c19_8 = t_r7_c19_4 + p_8_18;
  assign t_r7_c19_9 = t_r7_c19_5 + t_r7_c19_6;
  assign t_r7_c19_10 = t_r7_c19_7 + t_r7_c19_8;
  assign t_r7_c19_11 = t_r7_c19_9 + t_r7_c19_10;
  assign t_r7_c19_12 = t_r7_c19_11 + p_8_20;
  assign out_7_19 = t_r7_c19_12 >> 4;

  assign t_r7_c20_0 = p_6_20 << 1;
  assign t_r7_c20_1 = p_7_19 << 1;
  assign t_r7_c20_2 = p_7_20 << 2;
  assign t_r7_c20_3 = p_7_21 << 1;
  assign t_r7_c20_4 = p_8_20 << 1;
  assign t_r7_c20_5 = t_r7_c20_0 + p_6_19;
  assign t_r7_c20_6 = t_r7_c20_1 + p_6_21;
  assign t_r7_c20_7 = t_r7_c20_2 + t_r7_c20_3;
  assign t_r7_c20_8 = t_r7_c20_4 + p_8_19;
  assign t_r7_c20_9 = t_r7_c20_5 + t_r7_c20_6;
  assign t_r7_c20_10 = t_r7_c20_7 + t_r7_c20_8;
  assign t_r7_c20_11 = t_r7_c20_9 + t_r7_c20_10;
  assign t_r7_c20_12 = t_r7_c20_11 + p_8_21;
  assign out_7_20 = t_r7_c20_12 >> 4;

  assign t_r7_c21_0 = p_6_21 << 1;
  assign t_r7_c21_1 = p_7_20 << 1;
  assign t_r7_c21_2 = p_7_21 << 2;
  assign t_r7_c21_3 = p_7_22 << 1;
  assign t_r7_c21_4 = p_8_21 << 1;
  assign t_r7_c21_5 = t_r7_c21_0 + p_6_20;
  assign t_r7_c21_6 = t_r7_c21_1 + p_6_22;
  assign t_r7_c21_7 = t_r7_c21_2 + t_r7_c21_3;
  assign t_r7_c21_8 = t_r7_c21_4 + p_8_20;
  assign t_r7_c21_9 = t_r7_c21_5 + t_r7_c21_6;
  assign t_r7_c21_10 = t_r7_c21_7 + t_r7_c21_8;
  assign t_r7_c21_11 = t_r7_c21_9 + t_r7_c21_10;
  assign t_r7_c21_12 = t_r7_c21_11 + p_8_22;
  assign out_7_21 = t_r7_c21_12 >> 4;

  assign t_r7_c22_0 = p_6_22 << 1;
  assign t_r7_c22_1 = p_7_21 << 1;
  assign t_r7_c22_2 = p_7_22 << 2;
  assign t_r7_c22_3 = p_7_23 << 1;
  assign t_r7_c22_4 = p_8_22 << 1;
  assign t_r7_c22_5 = t_r7_c22_0 + p_6_21;
  assign t_r7_c22_6 = t_r7_c22_1 + p_6_23;
  assign t_r7_c22_7 = t_r7_c22_2 + t_r7_c22_3;
  assign t_r7_c22_8 = t_r7_c22_4 + p_8_21;
  assign t_r7_c22_9 = t_r7_c22_5 + t_r7_c22_6;
  assign t_r7_c22_10 = t_r7_c22_7 + t_r7_c22_8;
  assign t_r7_c22_11 = t_r7_c22_9 + t_r7_c22_10;
  assign t_r7_c22_12 = t_r7_c22_11 + p_8_23;
  assign out_7_22 = t_r7_c22_12 >> 4;

  assign t_r7_c23_0 = p_6_23 << 1;
  assign t_r7_c23_1 = p_7_22 << 1;
  assign t_r7_c23_2 = p_7_23 << 2;
  assign t_r7_c23_3 = p_7_24 << 1;
  assign t_r7_c23_4 = p_8_23 << 1;
  assign t_r7_c23_5 = t_r7_c23_0 + p_6_22;
  assign t_r7_c23_6 = t_r7_c23_1 + p_6_24;
  assign t_r7_c23_7 = t_r7_c23_2 + t_r7_c23_3;
  assign t_r7_c23_8 = t_r7_c23_4 + p_8_22;
  assign t_r7_c23_9 = t_r7_c23_5 + t_r7_c23_6;
  assign t_r7_c23_10 = t_r7_c23_7 + t_r7_c23_8;
  assign t_r7_c23_11 = t_r7_c23_9 + t_r7_c23_10;
  assign t_r7_c23_12 = t_r7_c23_11 + p_8_24;
  assign out_7_23 = t_r7_c23_12 >> 4;

  assign t_r7_c24_0 = p_6_24 << 1;
  assign t_r7_c24_1 = p_7_23 << 1;
  assign t_r7_c24_2 = p_7_24 << 2;
  assign t_r7_c24_3 = p_7_25 << 1;
  assign t_r7_c24_4 = p_8_24 << 1;
  assign t_r7_c24_5 = t_r7_c24_0 + p_6_23;
  assign t_r7_c24_6 = t_r7_c24_1 + p_6_25;
  assign t_r7_c24_7 = t_r7_c24_2 + t_r7_c24_3;
  assign t_r7_c24_8 = t_r7_c24_4 + p_8_23;
  assign t_r7_c24_9 = t_r7_c24_5 + t_r7_c24_6;
  assign t_r7_c24_10 = t_r7_c24_7 + t_r7_c24_8;
  assign t_r7_c24_11 = t_r7_c24_9 + t_r7_c24_10;
  assign t_r7_c24_12 = t_r7_c24_11 + p_8_25;
  assign out_7_24 = t_r7_c24_12 >> 4;

  assign t_r7_c25_0 = p_6_25 << 1;
  assign t_r7_c25_1 = p_7_24 << 1;
  assign t_r7_c25_2 = p_7_25 << 2;
  assign t_r7_c25_3 = p_7_26 << 1;
  assign t_r7_c25_4 = p_8_25 << 1;
  assign t_r7_c25_5 = t_r7_c25_0 + p_6_24;
  assign t_r7_c25_6 = t_r7_c25_1 + p_6_26;
  assign t_r7_c25_7 = t_r7_c25_2 + t_r7_c25_3;
  assign t_r7_c25_8 = t_r7_c25_4 + p_8_24;
  assign t_r7_c25_9 = t_r7_c25_5 + t_r7_c25_6;
  assign t_r7_c25_10 = t_r7_c25_7 + t_r7_c25_8;
  assign t_r7_c25_11 = t_r7_c25_9 + t_r7_c25_10;
  assign t_r7_c25_12 = t_r7_c25_11 + p_8_26;
  assign out_7_25 = t_r7_c25_12 >> 4;

  assign t_r7_c26_0 = p_6_26 << 1;
  assign t_r7_c26_1 = p_7_25 << 1;
  assign t_r7_c26_2 = p_7_26 << 2;
  assign t_r7_c26_3 = p_7_27 << 1;
  assign t_r7_c26_4 = p_8_26 << 1;
  assign t_r7_c26_5 = t_r7_c26_0 + p_6_25;
  assign t_r7_c26_6 = t_r7_c26_1 + p_6_27;
  assign t_r7_c26_7 = t_r7_c26_2 + t_r7_c26_3;
  assign t_r7_c26_8 = t_r7_c26_4 + p_8_25;
  assign t_r7_c26_9 = t_r7_c26_5 + t_r7_c26_6;
  assign t_r7_c26_10 = t_r7_c26_7 + t_r7_c26_8;
  assign t_r7_c26_11 = t_r7_c26_9 + t_r7_c26_10;
  assign t_r7_c26_12 = t_r7_c26_11 + p_8_27;
  assign out_7_26 = t_r7_c26_12 >> 4;

  assign t_r7_c27_0 = p_6_27 << 1;
  assign t_r7_c27_1 = p_7_26 << 1;
  assign t_r7_c27_2 = p_7_27 << 2;
  assign t_r7_c27_3 = p_7_28 << 1;
  assign t_r7_c27_4 = p_8_27 << 1;
  assign t_r7_c27_5 = t_r7_c27_0 + p_6_26;
  assign t_r7_c27_6 = t_r7_c27_1 + p_6_28;
  assign t_r7_c27_7 = t_r7_c27_2 + t_r7_c27_3;
  assign t_r7_c27_8 = t_r7_c27_4 + p_8_26;
  assign t_r7_c27_9 = t_r7_c27_5 + t_r7_c27_6;
  assign t_r7_c27_10 = t_r7_c27_7 + t_r7_c27_8;
  assign t_r7_c27_11 = t_r7_c27_9 + t_r7_c27_10;
  assign t_r7_c27_12 = t_r7_c27_11 + p_8_28;
  assign out_7_27 = t_r7_c27_12 >> 4;

  assign t_r7_c28_0 = p_6_28 << 1;
  assign t_r7_c28_1 = p_7_27 << 1;
  assign t_r7_c28_2 = p_7_28 << 2;
  assign t_r7_c28_3 = p_7_29 << 1;
  assign t_r7_c28_4 = p_8_28 << 1;
  assign t_r7_c28_5 = t_r7_c28_0 + p_6_27;
  assign t_r7_c28_6 = t_r7_c28_1 + p_6_29;
  assign t_r7_c28_7 = t_r7_c28_2 + t_r7_c28_3;
  assign t_r7_c28_8 = t_r7_c28_4 + p_8_27;
  assign t_r7_c28_9 = t_r7_c28_5 + t_r7_c28_6;
  assign t_r7_c28_10 = t_r7_c28_7 + t_r7_c28_8;
  assign t_r7_c28_11 = t_r7_c28_9 + t_r7_c28_10;
  assign t_r7_c28_12 = t_r7_c28_11 + p_8_29;
  assign out_7_28 = t_r7_c28_12 >> 4;

  assign t_r7_c29_0 = p_6_29 << 1;
  assign t_r7_c29_1 = p_7_28 << 1;
  assign t_r7_c29_2 = p_7_29 << 2;
  assign t_r7_c29_3 = p_7_30 << 1;
  assign t_r7_c29_4 = p_8_29 << 1;
  assign t_r7_c29_5 = t_r7_c29_0 + p_6_28;
  assign t_r7_c29_6 = t_r7_c29_1 + p_6_30;
  assign t_r7_c29_7 = t_r7_c29_2 + t_r7_c29_3;
  assign t_r7_c29_8 = t_r7_c29_4 + p_8_28;
  assign t_r7_c29_9 = t_r7_c29_5 + t_r7_c29_6;
  assign t_r7_c29_10 = t_r7_c29_7 + t_r7_c29_8;
  assign t_r7_c29_11 = t_r7_c29_9 + t_r7_c29_10;
  assign t_r7_c29_12 = t_r7_c29_11 + p_8_30;
  assign out_7_29 = t_r7_c29_12 >> 4;

  assign t_r7_c30_0 = p_6_30 << 1;
  assign t_r7_c30_1 = p_7_29 << 1;
  assign t_r7_c30_2 = p_7_30 << 2;
  assign t_r7_c30_3 = p_7_31 << 1;
  assign t_r7_c30_4 = p_8_30 << 1;
  assign t_r7_c30_5 = t_r7_c30_0 + p_6_29;
  assign t_r7_c30_6 = t_r7_c30_1 + p_6_31;
  assign t_r7_c30_7 = t_r7_c30_2 + t_r7_c30_3;
  assign t_r7_c30_8 = t_r7_c30_4 + p_8_29;
  assign t_r7_c30_9 = t_r7_c30_5 + t_r7_c30_6;
  assign t_r7_c30_10 = t_r7_c30_7 + t_r7_c30_8;
  assign t_r7_c30_11 = t_r7_c30_9 + t_r7_c30_10;
  assign t_r7_c30_12 = t_r7_c30_11 + p_8_31;
  assign out_7_30 = t_r7_c30_12 >> 4;

  assign t_r7_c31_0 = p_6_31 << 1;
  assign t_r7_c31_1 = p_7_30 << 1;
  assign t_r7_c31_2 = p_7_31 << 2;
  assign t_r7_c31_3 = p_7_32 << 1;
  assign t_r7_c31_4 = p_8_31 << 1;
  assign t_r7_c31_5 = t_r7_c31_0 + p_6_30;
  assign t_r7_c31_6 = t_r7_c31_1 + p_6_32;
  assign t_r7_c31_7 = t_r7_c31_2 + t_r7_c31_3;
  assign t_r7_c31_8 = t_r7_c31_4 + p_8_30;
  assign t_r7_c31_9 = t_r7_c31_5 + t_r7_c31_6;
  assign t_r7_c31_10 = t_r7_c31_7 + t_r7_c31_8;
  assign t_r7_c31_11 = t_r7_c31_9 + t_r7_c31_10;
  assign t_r7_c31_12 = t_r7_c31_11 + p_8_32;
  assign out_7_31 = t_r7_c31_12 >> 4;

  assign t_r7_c32_0 = p_6_32 << 1;
  assign t_r7_c32_1 = p_7_31 << 1;
  assign t_r7_c32_2 = p_7_32 << 2;
  assign t_r7_c32_3 = p_7_33 << 1;
  assign t_r7_c32_4 = p_8_32 << 1;
  assign t_r7_c32_5 = t_r7_c32_0 + p_6_31;
  assign t_r7_c32_6 = t_r7_c32_1 + p_6_33;
  assign t_r7_c32_7 = t_r7_c32_2 + t_r7_c32_3;
  assign t_r7_c32_8 = t_r7_c32_4 + p_8_31;
  assign t_r7_c32_9 = t_r7_c32_5 + t_r7_c32_6;
  assign t_r7_c32_10 = t_r7_c32_7 + t_r7_c32_8;
  assign t_r7_c32_11 = t_r7_c32_9 + t_r7_c32_10;
  assign t_r7_c32_12 = t_r7_c32_11 + p_8_33;
  assign out_7_32 = t_r7_c32_12 >> 4;

  assign t_r7_c33_0 = p_6_33 << 1;
  assign t_r7_c33_1 = p_7_32 << 1;
  assign t_r7_c33_2 = p_7_33 << 2;
  assign t_r7_c33_3 = p_7_34 << 1;
  assign t_r7_c33_4 = p_8_33 << 1;
  assign t_r7_c33_5 = t_r7_c33_0 + p_6_32;
  assign t_r7_c33_6 = t_r7_c33_1 + p_6_34;
  assign t_r7_c33_7 = t_r7_c33_2 + t_r7_c33_3;
  assign t_r7_c33_8 = t_r7_c33_4 + p_8_32;
  assign t_r7_c33_9 = t_r7_c33_5 + t_r7_c33_6;
  assign t_r7_c33_10 = t_r7_c33_7 + t_r7_c33_8;
  assign t_r7_c33_11 = t_r7_c33_9 + t_r7_c33_10;
  assign t_r7_c33_12 = t_r7_c33_11 + p_8_34;
  assign out_7_33 = t_r7_c33_12 >> 4;

  assign t_r7_c34_0 = p_6_34 << 1;
  assign t_r7_c34_1 = p_7_33 << 1;
  assign t_r7_c34_2 = p_7_34 << 2;
  assign t_r7_c34_3 = p_7_35 << 1;
  assign t_r7_c34_4 = p_8_34 << 1;
  assign t_r7_c34_5 = t_r7_c34_0 + p_6_33;
  assign t_r7_c34_6 = t_r7_c34_1 + p_6_35;
  assign t_r7_c34_7 = t_r7_c34_2 + t_r7_c34_3;
  assign t_r7_c34_8 = t_r7_c34_4 + p_8_33;
  assign t_r7_c34_9 = t_r7_c34_5 + t_r7_c34_6;
  assign t_r7_c34_10 = t_r7_c34_7 + t_r7_c34_8;
  assign t_r7_c34_11 = t_r7_c34_9 + t_r7_c34_10;
  assign t_r7_c34_12 = t_r7_c34_11 + p_8_35;
  assign out_7_34 = t_r7_c34_12 >> 4;

  assign t_r7_c35_0 = p_6_35 << 1;
  assign t_r7_c35_1 = p_7_34 << 1;
  assign t_r7_c35_2 = p_7_35 << 2;
  assign t_r7_c35_3 = p_7_36 << 1;
  assign t_r7_c35_4 = p_8_35 << 1;
  assign t_r7_c35_5 = t_r7_c35_0 + p_6_34;
  assign t_r7_c35_6 = t_r7_c35_1 + p_6_36;
  assign t_r7_c35_7 = t_r7_c35_2 + t_r7_c35_3;
  assign t_r7_c35_8 = t_r7_c35_4 + p_8_34;
  assign t_r7_c35_9 = t_r7_c35_5 + t_r7_c35_6;
  assign t_r7_c35_10 = t_r7_c35_7 + t_r7_c35_8;
  assign t_r7_c35_11 = t_r7_c35_9 + t_r7_c35_10;
  assign t_r7_c35_12 = t_r7_c35_11 + p_8_36;
  assign out_7_35 = t_r7_c35_12 >> 4;

  assign t_r7_c36_0 = p_6_36 << 1;
  assign t_r7_c36_1 = p_7_35 << 1;
  assign t_r7_c36_2 = p_7_36 << 2;
  assign t_r7_c36_3 = p_7_37 << 1;
  assign t_r7_c36_4 = p_8_36 << 1;
  assign t_r7_c36_5 = t_r7_c36_0 + p_6_35;
  assign t_r7_c36_6 = t_r7_c36_1 + p_6_37;
  assign t_r7_c36_7 = t_r7_c36_2 + t_r7_c36_3;
  assign t_r7_c36_8 = t_r7_c36_4 + p_8_35;
  assign t_r7_c36_9 = t_r7_c36_5 + t_r7_c36_6;
  assign t_r7_c36_10 = t_r7_c36_7 + t_r7_c36_8;
  assign t_r7_c36_11 = t_r7_c36_9 + t_r7_c36_10;
  assign t_r7_c36_12 = t_r7_c36_11 + p_8_37;
  assign out_7_36 = t_r7_c36_12 >> 4;

  assign t_r7_c37_0 = p_6_37 << 1;
  assign t_r7_c37_1 = p_7_36 << 1;
  assign t_r7_c37_2 = p_7_37 << 2;
  assign t_r7_c37_3 = p_7_38 << 1;
  assign t_r7_c37_4 = p_8_37 << 1;
  assign t_r7_c37_5 = t_r7_c37_0 + p_6_36;
  assign t_r7_c37_6 = t_r7_c37_1 + p_6_38;
  assign t_r7_c37_7 = t_r7_c37_2 + t_r7_c37_3;
  assign t_r7_c37_8 = t_r7_c37_4 + p_8_36;
  assign t_r7_c37_9 = t_r7_c37_5 + t_r7_c37_6;
  assign t_r7_c37_10 = t_r7_c37_7 + t_r7_c37_8;
  assign t_r7_c37_11 = t_r7_c37_9 + t_r7_c37_10;
  assign t_r7_c37_12 = t_r7_c37_11 + p_8_38;
  assign out_7_37 = t_r7_c37_12 >> 4;

  assign t_r7_c38_0 = p_6_38 << 1;
  assign t_r7_c38_1 = p_7_37 << 1;
  assign t_r7_c38_2 = p_7_38 << 2;
  assign t_r7_c38_3 = p_7_39 << 1;
  assign t_r7_c38_4 = p_8_38 << 1;
  assign t_r7_c38_5 = t_r7_c38_0 + p_6_37;
  assign t_r7_c38_6 = t_r7_c38_1 + p_6_39;
  assign t_r7_c38_7 = t_r7_c38_2 + t_r7_c38_3;
  assign t_r7_c38_8 = t_r7_c38_4 + p_8_37;
  assign t_r7_c38_9 = t_r7_c38_5 + t_r7_c38_6;
  assign t_r7_c38_10 = t_r7_c38_7 + t_r7_c38_8;
  assign t_r7_c38_11 = t_r7_c38_9 + t_r7_c38_10;
  assign t_r7_c38_12 = t_r7_c38_11 + p_8_39;
  assign out_7_38 = t_r7_c38_12 >> 4;

  assign t_r7_c39_0 = p_6_39 << 1;
  assign t_r7_c39_1 = p_7_38 << 1;
  assign t_r7_c39_2 = p_7_39 << 2;
  assign t_r7_c39_3 = p_7_40 << 1;
  assign t_r7_c39_4 = p_8_39 << 1;
  assign t_r7_c39_5 = t_r7_c39_0 + p_6_38;
  assign t_r7_c39_6 = t_r7_c39_1 + p_6_40;
  assign t_r7_c39_7 = t_r7_c39_2 + t_r7_c39_3;
  assign t_r7_c39_8 = t_r7_c39_4 + p_8_38;
  assign t_r7_c39_9 = t_r7_c39_5 + t_r7_c39_6;
  assign t_r7_c39_10 = t_r7_c39_7 + t_r7_c39_8;
  assign t_r7_c39_11 = t_r7_c39_9 + t_r7_c39_10;
  assign t_r7_c39_12 = t_r7_c39_11 + p_8_40;
  assign out_7_39 = t_r7_c39_12 >> 4;

  assign t_r7_c40_0 = p_6_40 << 1;
  assign t_r7_c40_1 = p_7_39 << 1;
  assign t_r7_c40_2 = p_7_40 << 2;
  assign t_r7_c40_3 = p_7_41 << 1;
  assign t_r7_c40_4 = p_8_40 << 1;
  assign t_r7_c40_5 = t_r7_c40_0 + p_6_39;
  assign t_r7_c40_6 = t_r7_c40_1 + p_6_41;
  assign t_r7_c40_7 = t_r7_c40_2 + t_r7_c40_3;
  assign t_r7_c40_8 = t_r7_c40_4 + p_8_39;
  assign t_r7_c40_9 = t_r7_c40_5 + t_r7_c40_6;
  assign t_r7_c40_10 = t_r7_c40_7 + t_r7_c40_8;
  assign t_r7_c40_11 = t_r7_c40_9 + t_r7_c40_10;
  assign t_r7_c40_12 = t_r7_c40_11 + p_8_41;
  assign out_7_40 = t_r7_c40_12 >> 4;

  assign t_r7_c41_0 = p_6_41 << 1;
  assign t_r7_c41_1 = p_7_40 << 1;
  assign t_r7_c41_2 = p_7_41 << 2;
  assign t_r7_c41_3 = p_7_42 << 1;
  assign t_r7_c41_4 = p_8_41 << 1;
  assign t_r7_c41_5 = t_r7_c41_0 + p_6_40;
  assign t_r7_c41_6 = t_r7_c41_1 + p_6_42;
  assign t_r7_c41_7 = t_r7_c41_2 + t_r7_c41_3;
  assign t_r7_c41_8 = t_r7_c41_4 + p_8_40;
  assign t_r7_c41_9 = t_r7_c41_5 + t_r7_c41_6;
  assign t_r7_c41_10 = t_r7_c41_7 + t_r7_c41_8;
  assign t_r7_c41_11 = t_r7_c41_9 + t_r7_c41_10;
  assign t_r7_c41_12 = t_r7_c41_11 + p_8_42;
  assign out_7_41 = t_r7_c41_12 >> 4;

  assign t_r7_c42_0 = p_6_42 << 1;
  assign t_r7_c42_1 = p_7_41 << 1;
  assign t_r7_c42_2 = p_7_42 << 2;
  assign t_r7_c42_3 = p_7_43 << 1;
  assign t_r7_c42_4 = p_8_42 << 1;
  assign t_r7_c42_5 = t_r7_c42_0 + p_6_41;
  assign t_r7_c42_6 = t_r7_c42_1 + p_6_43;
  assign t_r7_c42_7 = t_r7_c42_2 + t_r7_c42_3;
  assign t_r7_c42_8 = t_r7_c42_4 + p_8_41;
  assign t_r7_c42_9 = t_r7_c42_5 + t_r7_c42_6;
  assign t_r7_c42_10 = t_r7_c42_7 + t_r7_c42_8;
  assign t_r7_c42_11 = t_r7_c42_9 + t_r7_c42_10;
  assign t_r7_c42_12 = t_r7_c42_11 + p_8_43;
  assign out_7_42 = t_r7_c42_12 >> 4;

  assign t_r7_c43_0 = p_6_43 << 1;
  assign t_r7_c43_1 = p_7_42 << 1;
  assign t_r7_c43_2 = p_7_43 << 2;
  assign t_r7_c43_3 = p_7_44 << 1;
  assign t_r7_c43_4 = p_8_43 << 1;
  assign t_r7_c43_5 = t_r7_c43_0 + p_6_42;
  assign t_r7_c43_6 = t_r7_c43_1 + p_6_44;
  assign t_r7_c43_7 = t_r7_c43_2 + t_r7_c43_3;
  assign t_r7_c43_8 = t_r7_c43_4 + p_8_42;
  assign t_r7_c43_9 = t_r7_c43_5 + t_r7_c43_6;
  assign t_r7_c43_10 = t_r7_c43_7 + t_r7_c43_8;
  assign t_r7_c43_11 = t_r7_c43_9 + t_r7_c43_10;
  assign t_r7_c43_12 = t_r7_c43_11 + p_8_44;
  assign out_7_43 = t_r7_c43_12 >> 4;

  assign t_r7_c44_0 = p_6_44 << 1;
  assign t_r7_c44_1 = p_7_43 << 1;
  assign t_r7_c44_2 = p_7_44 << 2;
  assign t_r7_c44_3 = p_7_45 << 1;
  assign t_r7_c44_4 = p_8_44 << 1;
  assign t_r7_c44_5 = t_r7_c44_0 + p_6_43;
  assign t_r7_c44_6 = t_r7_c44_1 + p_6_45;
  assign t_r7_c44_7 = t_r7_c44_2 + t_r7_c44_3;
  assign t_r7_c44_8 = t_r7_c44_4 + p_8_43;
  assign t_r7_c44_9 = t_r7_c44_5 + t_r7_c44_6;
  assign t_r7_c44_10 = t_r7_c44_7 + t_r7_c44_8;
  assign t_r7_c44_11 = t_r7_c44_9 + t_r7_c44_10;
  assign t_r7_c44_12 = t_r7_c44_11 + p_8_45;
  assign out_7_44 = t_r7_c44_12 >> 4;

  assign t_r7_c45_0 = p_6_45 << 1;
  assign t_r7_c45_1 = p_7_44 << 1;
  assign t_r7_c45_2 = p_7_45 << 2;
  assign t_r7_c45_3 = p_7_46 << 1;
  assign t_r7_c45_4 = p_8_45 << 1;
  assign t_r7_c45_5 = t_r7_c45_0 + p_6_44;
  assign t_r7_c45_6 = t_r7_c45_1 + p_6_46;
  assign t_r7_c45_7 = t_r7_c45_2 + t_r7_c45_3;
  assign t_r7_c45_8 = t_r7_c45_4 + p_8_44;
  assign t_r7_c45_9 = t_r7_c45_5 + t_r7_c45_6;
  assign t_r7_c45_10 = t_r7_c45_7 + t_r7_c45_8;
  assign t_r7_c45_11 = t_r7_c45_9 + t_r7_c45_10;
  assign t_r7_c45_12 = t_r7_c45_11 + p_8_46;
  assign out_7_45 = t_r7_c45_12 >> 4;

  assign t_r7_c46_0 = p_6_46 << 1;
  assign t_r7_c46_1 = p_7_45 << 1;
  assign t_r7_c46_2 = p_7_46 << 2;
  assign t_r7_c46_3 = p_7_47 << 1;
  assign t_r7_c46_4 = p_8_46 << 1;
  assign t_r7_c46_5 = t_r7_c46_0 + p_6_45;
  assign t_r7_c46_6 = t_r7_c46_1 + p_6_47;
  assign t_r7_c46_7 = t_r7_c46_2 + t_r7_c46_3;
  assign t_r7_c46_8 = t_r7_c46_4 + p_8_45;
  assign t_r7_c46_9 = t_r7_c46_5 + t_r7_c46_6;
  assign t_r7_c46_10 = t_r7_c46_7 + t_r7_c46_8;
  assign t_r7_c46_11 = t_r7_c46_9 + t_r7_c46_10;
  assign t_r7_c46_12 = t_r7_c46_11 + p_8_47;
  assign out_7_46 = t_r7_c46_12 >> 4;

  assign t_r7_c47_0 = p_6_47 << 1;
  assign t_r7_c47_1 = p_7_46 << 1;
  assign t_r7_c47_2 = p_7_47 << 2;
  assign t_r7_c47_3 = p_7_48 << 1;
  assign t_r7_c47_4 = p_8_47 << 1;
  assign t_r7_c47_5 = t_r7_c47_0 + p_6_46;
  assign t_r7_c47_6 = t_r7_c47_1 + p_6_48;
  assign t_r7_c47_7 = t_r7_c47_2 + t_r7_c47_3;
  assign t_r7_c47_8 = t_r7_c47_4 + p_8_46;
  assign t_r7_c47_9 = t_r7_c47_5 + t_r7_c47_6;
  assign t_r7_c47_10 = t_r7_c47_7 + t_r7_c47_8;
  assign t_r7_c47_11 = t_r7_c47_9 + t_r7_c47_10;
  assign t_r7_c47_12 = t_r7_c47_11 + p_8_48;
  assign out_7_47 = t_r7_c47_12 >> 4;

  assign t_r7_c48_0 = p_6_48 << 1;
  assign t_r7_c48_1 = p_7_47 << 1;
  assign t_r7_c48_2 = p_7_48 << 2;
  assign t_r7_c48_3 = p_7_49 << 1;
  assign t_r7_c48_4 = p_8_48 << 1;
  assign t_r7_c48_5 = t_r7_c48_0 + p_6_47;
  assign t_r7_c48_6 = t_r7_c48_1 + p_6_49;
  assign t_r7_c48_7 = t_r7_c48_2 + t_r7_c48_3;
  assign t_r7_c48_8 = t_r7_c48_4 + p_8_47;
  assign t_r7_c48_9 = t_r7_c48_5 + t_r7_c48_6;
  assign t_r7_c48_10 = t_r7_c48_7 + t_r7_c48_8;
  assign t_r7_c48_11 = t_r7_c48_9 + t_r7_c48_10;
  assign t_r7_c48_12 = t_r7_c48_11 + p_8_49;
  assign out_7_48 = t_r7_c48_12 >> 4;

  assign t_r7_c49_0 = p_6_49 << 1;
  assign t_r7_c49_1 = p_7_48 << 1;
  assign t_r7_c49_2 = p_7_49 << 2;
  assign t_r7_c49_3 = p_7_50 << 1;
  assign t_r7_c49_4 = p_8_49 << 1;
  assign t_r7_c49_5 = t_r7_c49_0 + p_6_48;
  assign t_r7_c49_6 = t_r7_c49_1 + p_6_50;
  assign t_r7_c49_7 = t_r7_c49_2 + t_r7_c49_3;
  assign t_r7_c49_8 = t_r7_c49_4 + p_8_48;
  assign t_r7_c49_9 = t_r7_c49_5 + t_r7_c49_6;
  assign t_r7_c49_10 = t_r7_c49_7 + t_r7_c49_8;
  assign t_r7_c49_11 = t_r7_c49_9 + t_r7_c49_10;
  assign t_r7_c49_12 = t_r7_c49_11 + p_8_50;
  assign out_7_49 = t_r7_c49_12 >> 4;

  assign t_r7_c50_0 = p_6_50 << 1;
  assign t_r7_c50_1 = p_7_49 << 1;
  assign t_r7_c50_2 = p_7_50 << 2;
  assign t_r7_c50_3 = p_7_51 << 1;
  assign t_r7_c50_4 = p_8_50 << 1;
  assign t_r7_c50_5 = t_r7_c50_0 + p_6_49;
  assign t_r7_c50_6 = t_r7_c50_1 + p_6_51;
  assign t_r7_c50_7 = t_r7_c50_2 + t_r7_c50_3;
  assign t_r7_c50_8 = t_r7_c50_4 + p_8_49;
  assign t_r7_c50_9 = t_r7_c50_5 + t_r7_c50_6;
  assign t_r7_c50_10 = t_r7_c50_7 + t_r7_c50_8;
  assign t_r7_c50_11 = t_r7_c50_9 + t_r7_c50_10;
  assign t_r7_c50_12 = t_r7_c50_11 + p_8_51;
  assign out_7_50 = t_r7_c50_12 >> 4;

  assign t_r7_c51_0 = p_6_51 << 1;
  assign t_r7_c51_1 = p_7_50 << 1;
  assign t_r7_c51_2 = p_7_51 << 2;
  assign t_r7_c51_3 = p_7_52 << 1;
  assign t_r7_c51_4 = p_8_51 << 1;
  assign t_r7_c51_5 = t_r7_c51_0 + p_6_50;
  assign t_r7_c51_6 = t_r7_c51_1 + p_6_52;
  assign t_r7_c51_7 = t_r7_c51_2 + t_r7_c51_3;
  assign t_r7_c51_8 = t_r7_c51_4 + p_8_50;
  assign t_r7_c51_9 = t_r7_c51_5 + t_r7_c51_6;
  assign t_r7_c51_10 = t_r7_c51_7 + t_r7_c51_8;
  assign t_r7_c51_11 = t_r7_c51_9 + t_r7_c51_10;
  assign t_r7_c51_12 = t_r7_c51_11 + p_8_52;
  assign out_7_51 = t_r7_c51_12 >> 4;

  assign t_r7_c52_0 = p_6_52 << 1;
  assign t_r7_c52_1 = p_7_51 << 1;
  assign t_r7_c52_2 = p_7_52 << 2;
  assign t_r7_c52_3 = p_7_53 << 1;
  assign t_r7_c52_4 = p_8_52 << 1;
  assign t_r7_c52_5 = t_r7_c52_0 + p_6_51;
  assign t_r7_c52_6 = t_r7_c52_1 + p_6_53;
  assign t_r7_c52_7 = t_r7_c52_2 + t_r7_c52_3;
  assign t_r7_c52_8 = t_r7_c52_4 + p_8_51;
  assign t_r7_c52_9 = t_r7_c52_5 + t_r7_c52_6;
  assign t_r7_c52_10 = t_r7_c52_7 + t_r7_c52_8;
  assign t_r7_c52_11 = t_r7_c52_9 + t_r7_c52_10;
  assign t_r7_c52_12 = t_r7_c52_11 + p_8_53;
  assign out_7_52 = t_r7_c52_12 >> 4;

  assign t_r7_c53_0 = p_6_53 << 1;
  assign t_r7_c53_1 = p_7_52 << 1;
  assign t_r7_c53_2 = p_7_53 << 2;
  assign t_r7_c53_3 = p_7_54 << 1;
  assign t_r7_c53_4 = p_8_53 << 1;
  assign t_r7_c53_5 = t_r7_c53_0 + p_6_52;
  assign t_r7_c53_6 = t_r7_c53_1 + p_6_54;
  assign t_r7_c53_7 = t_r7_c53_2 + t_r7_c53_3;
  assign t_r7_c53_8 = t_r7_c53_4 + p_8_52;
  assign t_r7_c53_9 = t_r7_c53_5 + t_r7_c53_6;
  assign t_r7_c53_10 = t_r7_c53_7 + t_r7_c53_8;
  assign t_r7_c53_11 = t_r7_c53_9 + t_r7_c53_10;
  assign t_r7_c53_12 = t_r7_c53_11 + p_8_54;
  assign out_7_53 = t_r7_c53_12 >> 4;

  assign t_r7_c54_0 = p_6_54 << 1;
  assign t_r7_c54_1 = p_7_53 << 1;
  assign t_r7_c54_2 = p_7_54 << 2;
  assign t_r7_c54_3 = p_7_55 << 1;
  assign t_r7_c54_4 = p_8_54 << 1;
  assign t_r7_c54_5 = t_r7_c54_0 + p_6_53;
  assign t_r7_c54_6 = t_r7_c54_1 + p_6_55;
  assign t_r7_c54_7 = t_r7_c54_2 + t_r7_c54_3;
  assign t_r7_c54_8 = t_r7_c54_4 + p_8_53;
  assign t_r7_c54_9 = t_r7_c54_5 + t_r7_c54_6;
  assign t_r7_c54_10 = t_r7_c54_7 + t_r7_c54_8;
  assign t_r7_c54_11 = t_r7_c54_9 + t_r7_c54_10;
  assign t_r7_c54_12 = t_r7_c54_11 + p_8_55;
  assign out_7_54 = t_r7_c54_12 >> 4;

  assign t_r7_c55_0 = p_6_55 << 1;
  assign t_r7_c55_1 = p_7_54 << 1;
  assign t_r7_c55_2 = p_7_55 << 2;
  assign t_r7_c55_3 = p_7_56 << 1;
  assign t_r7_c55_4 = p_8_55 << 1;
  assign t_r7_c55_5 = t_r7_c55_0 + p_6_54;
  assign t_r7_c55_6 = t_r7_c55_1 + p_6_56;
  assign t_r7_c55_7 = t_r7_c55_2 + t_r7_c55_3;
  assign t_r7_c55_8 = t_r7_c55_4 + p_8_54;
  assign t_r7_c55_9 = t_r7_c55_5 + t_r7_c55_6;
  assign t_r7_c55_10 = t_r7_c55_7 + t_r7_c55_8;
  assign t_r7_c55_11 = t_r7_c55_9 + t_r7_c55_10;
  assign t_r7_c55_12 = t_r7_c55_11 + p_8_56;
  assign out_7_55 = t_r7_c55_12 >> 4;

  assign t_r7_c56_0 = p_6_56 << 1;
  assign t_r7_c56_1 = p_7_55 << 1;
  assign t_r7_c56_2 = p_7_56 << 2;
  assign t_r7_c56_3 = p_7_57 << 1;
  assign t_r7_c56_4 = p_8_56 << 1;
  assign t_r7_c56_5 = t_r7_c56_0 + p_6_55;
  assign t_r7_c56_6 = t_r7_c56_1 + p_6_57;
  assign t_r7_c56_7 = t_r7_c56_2 + t_r7_c56_3;
  assign t_r7_c56_8 = t_r7_c56_4 + p_8_55;
  assign t_r7_c56_9 = t_r7_c56_5 + t_r7_c56_6;
  assign t_r7_c56_10 = t_r7_c56_7 + t_r7_c56_8;
  assign t_r7_c56_11 = t_r7_c56_9 + t_r7_c56_10;
  assign t_r7_c56_12 = t_r7_c56_11 + p_8_57;
  assign out_7_56 = t_r7_c56_12 >> 4;

  assign t_r7_c57_0 = p_6_57 << 1;
  assign t_r7_c57_1 = p_7_56 << 1;
  assign t_r7_c57_2 = p_7_57 << 2;
  assign t_r7_c57_3 = p_7_58 << 1;
  assign t_r7_c57_4 = p_8_57 << 1;
  assign t_r7_c57_5 = t_r7_c57_0 + p_6_56;
  assign t_r7_c57_6 = t_r7_c57_1 + p_6_58;
  assign t_r7_c57_7 = t_r7_c57_2 + t_r7_c57_3;
  assign t_r7_c57_8 = t_r7_c57_4 + p_8_56;
  assign t_r7_c57_9 = t_r7_c57_5 + t_r7_c57_6;
  assign t_r7_c57_10 = t_r7_c57_7 + t_r7_c57_8;
  assign t_r7_c57_11 = t_r7_c57_9 + t_r7_c57_10;
  assign t_r7_c57_12 = t_r7_c57_11 + p_8_58;
  assign out_7_57 = t_r7_c57_12 >> 4;

  assign t_r7_c58_0 = p_6_58 << 1;
  assign t_r7_c58_1 = p_7_57 << 1;
  assign t_r7_c58_2 = p_7_58 << 2;
  assign t_r7_c58_3 = p_7_59 << 1;
  assign t_r7_c58_4 = p_8_58 << 1;
  assign t_r7_c58_5 = t_r7_c58_0 + p_6_57;
  assign t_r7_c58_6 = t_r7_c58_1 + p_6_59;
  assign t_r7_c58_7 = t_r7_c58_2 + t_r7_c58_3;
  assign t_r7_c58_8 = t_r7_c58_4 + p_8_57;
  assign t_r7_c58_9 = t_r7_c58_5 + t_r7_c58_6;
  assign t_r7_c58_10 = t_r7_c58_7 + t_r7_c58_8;
  assign t_r7_c58_11 = t_r7_c58_9 + t_r7_c58_10;
  assign t_r7_c58_12 = t_r7_c58_11 + p_8_59;
  assign out_7_58 = t_r7_c58_12 >> 4;

  assign t_r7_c59_0 = p_6_59 << 1;
  assign t_r7_c59_1 = p_7_58 << 1;
  assign t_r7_c59_2 = p_7_59 << 2;
  assign t_r7_c59_3 = p_7_60 << 1;
  assign t_r7_c59_4 = p_8_59 << 1;
  assign t_r7_c59_5 = t_r7_c59_0 + p_6_58;
  assign t_r7_c59_6 = t_r7_c59_1 + p_6_60;
  assign t_r7_c59_7 = t_r7_c59_2 + t_r7_c59_3;
  assign t_r7_c59_8 = t_r7_c59_4 + p_8_58;
  assign t_r7_c59_9 = t_r7_c59_5 + t_r7_c59_6;
  assign t_r7_c59_10 = t_r7_c59_7 + t_r7_c59_8;
  assign t_r7_c59_11 = t_r7_c59_9 + t_r7_c59_10;
  assign t_r7_c59_12 = t_r7_c59_11 + p_8_60;
  assign out_7_59 = t_r7_c59_12 >> 4;

  assign t_r7_c60_0 = p_6_60 << 1;
  assign t_r7_c60_1 = p_7_59 << 1;
  assign t_r7_c60_2 = p_7_60 << 2;
  assign t_r7_c60_3 = p_7_61 << 1;
  assign t_r7_c60_4 = p_8_60 << 1;
  assign t_r7_c60_5 = t_r7_c60_0 + p_6_59;
  assign t_r7_c60_6 = t_r7_c60_1 + p_6_61;
  assign t_r7_c60_7 = t_r7_c60_2 + t_r7_c60_3;
  assign t_r7_c60_8 = t_r7_c60_4 + p_8_59;
  assign t_r7_c60_9 = t_r7_c60_5 + t_r7_c60_6;
  assign t_r7_c60_10 = t_r7_c60_7 + t_r7_c60_8;
  assign t_r7_c60_11 = t_r7_c60_9 + t_r7_c60_10;
  assign t_r7_c60_12 = t_r7_c60_11 + p_8_61;
  assign out_7_60 = t_r7_c60_12 >> 4;

  assign t_r7_c61_0 = p_6_61 << 1;
  assign t_r7_c61_1 = p_7_60 << 1;
  assign t_r7_c61_2 = p_7_61 << 2;
  assign t_r7_c61_3 = p_7_62 << 1;
  assign t_r7_c61_4 = p_8_61 << 1;
  assign t_r7_c61_5 = t_r7_c61_0 + p_6_60;
  assign t_r7_c61_6 = t_r7_c61_1 + p_6_62;
  assign t_r7_c61_7 = t_r7_c61_2 + t_r7_c61_3;
  assign t_r7_c61_8 = t_r7_c61_4 + p_8_60;
  assign t_r7_c61_9 = t_r7_c61_5 + t_r7_c61_6;
  assign t_r7_c61_10 = t_r7_c61_7 + t_r7_c61_8;
  assign t_r7_c61_11 = t_r7_c61_9 + t_r7_c61_10;
  assign t_r7_c61_12 = t_r7_c61_11 + p_8_62;
  assign out_7_61 = t_r7_c61_12 >> 4;

  assign t_r7_c62_0 = p_6_62 << 1;
  assign t_r7_c62_1 = p_7_61 << 1;
  assign t_r7_c62_2 = p_7_62 << 2;
  assign t_r7_c62_3 = p_7_63 << 1;
  assign t_r7_c62_4 = p_8_62 << 1;
  assign t_r7_c62_5 = t_r7_c62_0 + p_6_61;
  assign t_r7_c62_6 = t_r7_c62_1 + p_6_63;
  assign t_r7_c62_7 = t_r7_c62_2 + t_r7_c62_3;
  assign t_r7_c62_8 = t_r7_c62_4 + p_8_61;
  assign t_r7_c62_9 = t_r7_c62_5 + t_r7_c62_6;
  assign t_r7_c62_10 = t_r7_c62_7 + t_r7_c62_8;
  assign t_r7_c62_11 = t_r7_c62_9 + t_r7_c62_10;
  assign t_r7_c62_12 = t_r7_c62_11 + p_8_63;
  assign out_7_62 = t_r7_c62_12 >> 4;

  assign t_r7_c63_0 = p_6_63 << 1;
  assign t_r7_c63_1 = p_7_62 << 1;
  assign t_r7_c63_2 = p_7_63 << 2;
  assign t_r7_c63_3 = p_7_64 << 1;
  assign t_r7_c63_4 = p_8_63 << 1;
  assign t_r7_c63_5 = t_r7_c63_0 + p_6_62;
  assign t_r7_c63_6 = t_r7_c63_1 + p_6_64;
  assign t_r7_c63_7 = t_r7_c63_2 + t_r7_c63_3;
  assign t_r7_c63_8 = t_r7_c63_4 + p_8_62;
  assign t_r7_c63_9 = t_r7_c63_5 + t_r7_c63_6;
  assign t_r7_c63_10 = t_r7_c63_7 + t_r7_c63_8;
  assign t_r7_c63_11 = t_r7_c63_9 + t_r7_c63_10;
  assign t_r7_c63_12 = t_r7_c63_11 + p_8_64;
  assign out_7_63 = t_r7_c63_12 >> 4;

  assign t_r7_c64_0 = p_6_64 << 1;
  assign t_r7_c64_1 = p_7_63 << 1;
  assign t_r7_c64_2 = p_7_64 << 2;
  assign t_r7_c64_3 = p_7_65 << 1;
  assign t_r7_c64_4 = p_8_64 << 1;
  assign t_r7_c64_5 = t_r7_c64_0 + p_6_63;
  assign t_r7_c64_6 = t_r7_c64_1 + p_6_65;
  assign t_r7_c64_7 = t_r7_c64_2 + t_r7_c64_3;
  assign t_r7_c64_8 = t_r7_c64_4 + p_8_63;
  assign t_r7_c64_9 = t_r7_c64_5 + t_r7_c64_6;
  assign t_r7_c64_10 = t_r7_c64_7 + t_r7_c64_8;
  assign t_r7_c64_11 = t_r7_c64_9 + t_r7_c64_10;
  assign t_r7_c64_12 = t_r7_c64_11 + p_8_65;
  assign out_7_64 = t_r7_c64_12 >> 4;

  assign t_r8_c1_0 = p_7_1 << 1;
  assign t_r8_c1_1 = p_8_0 << 1;
  assign t_r8_c1_2 = p_8_1 << 2;
  assign t_r8_c1_3 = p_8_2 << 1;
  assign t_r8_c1_4 = p_9_1 << 1;
  assign t_r8_c1_5 = t_r8_c1_0 + p_7_0;
  assign t_r8_c1_6 = t_r8_c1_1 + p_7_2;
  assign t_r8_c1_7 = t_r8_c1_2 + t_r8_c1_3;
  assign t_r8_c1_8 = t_r8_c1_4 + p_9_0;
  assign t_r8_c1_9 = t_r8_c1_5 + t_r8_c1_6;
  assign t_r8_c1_10 = t_r8_c1_7 + t_r8_c1_8;
  assign t_r8_c1_11 = t_r8_c1_9 + t_r8_c1_10;
  assign t_r8_c1_12 = t_r8_c1_11 + p_9_2;
  assign out_8_1 = t_r8_c1_12 >> 4;

  assign t_r8_c2_0 = p_7_2 << 1;
  assign t_r8_c2_1 = p_8_1 << 1;
  assign t_r8_c2_2 = p_8_2 << 2;
  assign t_r8_c2_3 = p_8_3 << 1;
  assign t_r8_c2_4 = p_9_2 << 1;
  assign t_r8_c2_5 = t_r8_c2_0 + p_7_1;
  assign t_r8_c2_6 = t_r8_c2_1 + p_7_3;
  assign t_r8_c2_7 = t_r8_c2_2 + t_r8_c2_3;
  assign t_r8_c2_8 = t_r8_c2_4 + p_9_1;
  assign t_r8_c2_9 = t_r8_c2_5 + t_r8_c2_6;
  assign t_r8_c2_10 = t_r8_c2_7 + t_r8_c2_8;
  assign t_r8_c2_11 = t_r8_c2_9 + t_r8_c2_10;
  assign t_r8_c2_12 = t_r8_c2_11 + p_9_3;
  assign out_8_2 = t_r8_c2_12 >> 4;

  assign t_r8_c3_0 = p_7_3 << 1;
  assign t_r8_c3_1 = p_8_2 << 1;
  assign t_r8_c3_2 = p_8_3 << 2;
  assign t_r8_c3_3 = p_8_4 << 1;
  assign t_r8_c3_4 = p_9_3 << 1;
  assign t_r8_c3_5 = t_r8_c3_0 + p_7_2;
  assign t_r8_c3_6 = t_r8_c3_1 + p_7_4;
  assign t_r8_c3_7 = t_r8_c3_2 + t_r8_c3_3;
  assign t_r8_c3_8 = t_r8_c3_4 + p_9_2;
  assign t_r8_c3_9 = t_r8_c3_5 + t_r8_c3_6;
  assign t_r8_c3_10 = t_r8_c3_7 + t_r8_c3_8;
  assign t_r8_c3_11 = t_r8_c3_9 + t_r8_c3_10;
  assign t_r8_c3_12 = t_r8_c3_11 + p_9_4;
  assign out_8_3 = t_r8_c3_12 >> 4;

  assign t_r8_c4_0 = p_7_4 << 1;
  assign t_r8_c4_1 = p_8_3 << 1;
  assign t_r8_c4_2 = p_8_4 << 2;
  assign t_r8_c4_3 = p_8_5 << 1;
  assign t_r8_c4_4 = p_9_4 << 1;
  assign t_r8_c4_5 = t_r8_c4_0 + p_7_3;
  assign t_r8_c4_6 = t_r8_c4_1 + p_7_5;
  assign t_r8_c4_7 = t_r8_c4_2 + t_r8_c4_3;
  assign t_r8_c4_8 = t_r8_c4_4 + p_9_3;
  assign t_r8_c4_9 = t_r8_c4_5 + t_r8_c4_6;
  assign t_r8_c4_10 = t_r8_c4_7 + t_r8_c4_8;
  assign t_r8_c4_11 = t_r8_c4_9 + t_r8_c4_10;
  assign t_r8_c4_12 = t_r8_c4_11 + p_9_5;
  assign out_8_4 = t_r8_c4_12 >> 4;

  assign t_r8_c5_0 = p_7_5 << 1;
  assign t_r8_c5_1 = p_8_4 << 1;
  assign t_r8_c5_2 = p_8_5 << 2;
  assign t_r8_c5_3 = p_8_6 << 1;
  assign t_r8_c5_4 = p_9_5 << 1;
  assign t_r8_c5_5 = t_r8_c5_0 + p_7_4;
  assign t_r8_c5_6 = t_r8_c5_1 + p_7_6;
  assign t_r8_c5_7 = t_r8_c5_2 + t_r8_c5_3;
  assign t_r8_c5_8 = t_r8_c5_4 + p_9_4;
  assign t_r8_c5_9 = t_r8_c5_5 + t_r8_c5_6;
  assign t_r8_c5_10 = t_r8_c5_7 + t_r8_c5_8;
  assign t_r8_c5_11 = t_r8_c5_9 + t_r8_c5_10;
  assign t_r8_c5_12 = t_r8_c5_11 + p_9_6;
  assign out_8_5 = t_r8_c5_12 >> 4;

  assign t_r8_c6_0 = p_7_6 << 1;
  assign t_r8_c6_1 = p_8_5 << 1;
  assign t_r8_c6_2 = p_8_6 << 2;
  assign t_r8_c6_3 = p_8_7 << 1;
  assign t_r8_c6_4 = p_9_6 << 1;
  assign t_r8_c6_5 = t_r8_c6_0 + p_7_5;
  assign t_r8_c6_6 = t_r8_c6_1 + p_7_7;
  assign t_r8_c6_7 = t_r8_c6_2 + t_r8_c6_3;
  assign t_r8_c6_8 = t_r8_c6_4 + p_9_5;
  assign t_r8_c6_9 = t_r8_c6_5 + t_r8_c6_6;
  assign t_r8_c6_10 = t_r8_c6_7 + t_r8_c6_8;
  assign t_r8_c6_11 = t_r8_c6_9 + t_r8_c6_10;
  assign t_r8_c6_12 = t_r8_c6_11 + p_9_7;
  assign out_8_6 = t_r8_c6_12 >> 4;

  assign t_r8_c7_0 = p_7_7 << 1;
  assign t_r8_c7_1 = p_8_6 << 1;
  assign t_r8_c7_2 = p_8_7 << 2;
  assign t_r8_c7_3 = p_8_8 << 1;
  assign t_r8_c7_4 = p_9_7 << 1;
  assign t_r8_c7_5 = t_r8_c7_0 + p_7_6;
  assign t_r8_c7_6 = t_r8_c7_1 + p_7_8;
  assign t_r8_c7_7 = t_r8_c7_2 + t_r8_c7_3;
  assign t_r8_c7_8 = t_r8_c7_4 + p_9_6;
  assign t_r8_c7_9 = t_r8_c7_5 + t_r8_c7_6;
  assign t_r8_c7_10 = t_r8_c7_7 + t_r8_c7_8;
  assign t_r8_c7_11 = t_r8_c7_9 + t_r8_c7_10;
  assign t_r8_c7_12 = t_r8_c7_11 + p_9_8;
  assign out_8_7 = t_r8_c7_12 >> 4;

  assign t_r8_c8_0 = p_7_8 << 1;
  assign t_r8_c8_1 = p_8_7 << 1;
  assign t_r8_c8_2 = p_8_8 << 2;
  assign t_r8_c8_3 = p_8_9 << 1;
  assign t_r8_c8_4 = p_9_8 << 1;
  assign t_r8_c8_5 = t_r8_c8_0 + p_7_7;
  assign t_r8_c8_6 = t_r8_c8_1 + p_7_9;
  assign t_r8_c8_7 = t_r8_c8_2 + t_r8_c8_3;
  assign t_r8_c8_8 = t_r8_c8_4 + p_9_7;
  assign t_r8_c8_9 = t_r8_c8_5 + t_r8_c8_6;
  assign t_r8_c8_10 = t_r8_c8_7 + t_r8_c8_8;
  assign t_r8_c8_11 = t_r8_c8_9 + t_r8_c8_10;
  assign t_r8_c8_12 = t_r8_c8_11 + p_9_9;
  assign out_8_8 = t_r8_c8_12 >> 4;

  assign t_r8_c9_0 = p_7_9 << 1;
  assign t_r8_c9_1 = p_8_8 << 1;
  assign t_r8_c9_2 = p_8_9 << 2;
  assign t_r8_c9_3 = p_8_10 << 1;
  assign t_r8_c9_4 = p_9_9 << 1;
  assign t_r8_c9_5 = t_r8_c9_0 + p_7_8;
  assign t_r8_c9_6 = t_r8_c9_1 + p_7_10;
  assign t_r8_c9_7 = t_r8_c9_2 + t_r8_c9_3;
  assign t_r8_c9_8 = t_r8_c9_4 + p_9_8;
  assign t_r8_c9_9 = t_r8_c9_5 + t_r8_c9_6;
  assign t_r8_c9_10 = t_r8_c9_7 + t_r8_c9_8;
  assign t_r8_c9_11 = t_r8_c9_9 + t_r8_c9_10;
  assign t_r8_c9_12 = t_r8_c9_11 + p_9_10;
  assign out_8_9 = t_r8_c9_12 >> 4;

  assign t_r8_c10_0 = p_7_10 << 1;
  assign t_r8_c10_1 = p_8_9 << 1;
  assign t_r8_c10_2 = p_8_10 << 2;
  assign t_r8_c10_3 = p_8_11 << 1;
  assign t_r8_c10_4 = p_9_10 << 1;
  assign t_r8_c10_5 = t_r8_c10_0 + p_7_9;
  assign t_r8_c10_6 = t_r8_c10_1 + p_7_11;
  assign t_r8_c10_7 = t_r8_c10_2 + t_r8_c10_3;
  assign t_r8_c10_8 = t_r8_c10_4 + p_9_9;
  assign t_r8_c10_9 = t_r8_c10_5 + t_r8_c10_6;
  assign t_r8_c10_10 = t_r8_c10_7 + t_r8_c10_8;
  assign t_r8_c10_11 = t_r8_c10_9 + t_r8_c10_10;
  assign t_r8_c10_12 = t_r8_c10_11 + p_9_11;
  assign out_8_10 = t_r8_c10_12 >> 4;

  assign t_r8_c11_0 = p_7_11 << 1;
  assign t_r8_c11_1 = p_8_10 << 1;
  assign t_r8_c11_2 = p_8_11 << 2;
  assign t_r8_c11_3 = p_8_12 << 1;
  assign t_r8_c11_4 = p_9_11 << 1;
  assign t_r8_c11_5 = t_r8_c11_0 + p_7_10;
  assign t_r8_c11_6 = t_r8_c11_1 + p_7_12;
  assign t_r8_c11_7 = t_r8_c11_2 + t_r8_c11_3;
  assign t_r8_c11_8 = t_r8_c11_4 + p_9_10;
  assign t_r8_c11_9 = t_r8_c11_5 + t_r8_c11_6;
  assign t_r8_c11_10 = t_r8_c11_7 + t_r8_c11_8;
  assign t_r8_c11_11 = t_r8_c11_9 + t_r8_c11_10;
  assign t_r8_c11_12 = t_r8_c11_11 + p_9_12;
  assign out_8_11 = t_r8_c11_12 >> 4;

  assign t_r8_c12_0 = p_7_12 << 1;
  assign t_r8_c12_1 = p_8_11 << 1;
  assign t_r8_c12_2 = p_8_12 << 2;
  assign t_r8_c12_3 = p_8_13 << 1;
  assign t_r8_c12_4 = p_9_12 << 1;
  assign t_r8_c12_5 = t_r8_c12_0 + p_7_11;
  assign t_r8_c12_6 = t_r8_c12_1 + p_7_13;
  assign t_r8_c12_7 = t_r8_c12_2 + t_r8_c12_3;
  assign t_r8_c12_8 = t_r8_c12_4 + p_9_11;
  assign t_r8_c12_9 = t_r8_c12_5 + t_r8_c12_6;
  assign t_r8_c12_10 = t_r8_c12_7 + t_r8_c12_8;
  assign t_r8_c12_11 = t_r8_c12_9 + t_r8_c12_10;
  assign t_r8_c12_12 = t_r8_c12_11 + p_9_13;
  assign out_8_12 = t_r8_c12_12 >> 4;

  assign t_r8_c13_0 = p_7_13 << 1;
  assign t_r8_c13_1 = p_8_12 << 1;
  assign t_r8_c13_2 = p_8_13 << 2;
  assign t_r8_c13_3 = p_8_14 << 1;
  assign t_r8_c13_4 = p_9_13 << 1;
  assign t_r8_c13_5 = t_r8_c13_0 + p_7_12;
  assign t_r8_c13_6 = t_r8_c13_1 + p_7_14;
  assign t_r8_c13_7 = t_r8_c13_2 + t_r8_c13_3;
  assign t_r8_c13_8 = t_r8_c13_4 + p_9_12;
  assign t_r8_c13_9 = t_r8_c13_5 + t_r8_c13_6;
  assign t_r8_c13_10 = t_r8_c13_7 + t_r8_c13_8;
  assign t_r8_c13_11 = t_r8_c13_9 + t_r8_c13_10;
  assign t_r8_c13_12 = t_r8_c13_11 + p_9_14;
  assign out_8_13 = t_r8_c13_12 >> 4;

  assign t_r8_c14_0 = p_7_14 << 1;
  assign t_r8_c14_1 = p_8_13 << 1;
  assign t_r8_c14_2 = p_8_14 << 2;
  assign t_r8_c14_3 = p_8_15 << 1;
  assign t_r8_c14_4 = p_9_14 << 1;
  assign t_r8_c14_5 = t_r8_c14_0 + p_7_13;
  assign t_r8_c14_6 = t_r8_c14_1 + p_7_15;
  assign t_r8_c14_7 = t_r8_c14_2 + t_r8_c14_3;
  assign t_r8_c14_8 = t_r8_c14_4 + p_9_13;
  assign t_r8_c14_9 = t_r8_c14_5 + t_r8_c14_6;
  assign t_r8_c14_10 = t_r8_c14_7 + t_r8_c14_8;
  assign t_r8_c14_11 = t_r8_c14_9 + t_r8_c14_10;
  assign t_r8_c14_12 = t_r8_c14_11 + p_9_15;
  assign out_8_14 = t_r8_c14_12 >> 4;

  assign t_r8_c15_0 = p_7_15 << 1;
  assign t_r8_c15_1 = p_8_14 << 1;
  assign t_r8_c15_2 = p_8_15 << 2;
  assign t_r8_c15_3 = p_8_16 << 1;
  assign t_r8_c15_4 = p_9_15 << 1;
  assign t_r8_c15_5 = t_r8_c15_0 + p_7_14;
  assign t_r8_c15_6 = t_r8_c15_1 + p_7_16;
  assign t_r8_c15_7 = t_r8_c15_2 + t_r8_c15_3;
  assign t_r8_c15_8 = t_r8_c15_4 + p_9_14;
  assign t_r8_c15_9 = t_r8_c15_5 + t_r8_c15_6;
  assign t_r8_c15_10 = t_r8_c15_7 + t_r8_c15_8;
  assign t_r8_c15_11 = t_r8_c15_9 + t_r8_c15_10;
  assign t_r8_c15_12 = t_r8_c15_11 + p_9_16;
  assign out_8_15 = t_r8_c15_12 >> 4;

  assign t_r8_c16_0 = p_7_16 << 1;
  assign t_r8_c16_1 = p_8_15 << 1;
  assign t_r8_c16_2 = p_8_16 << 2;
  assign t_r8_c16_3 = p_8_17 << 1;
  assign t_r8_c16_4 = p_9_16 << 1;
  assign t_r8_c16_5 = t_r8_c16_0 + p_7_15;
  assign t_r8_c16_6 = t_r8_c16_1 + p_7_17;
  assign t_r8_c16_7 = t_r8_c16_2 + t_r8_c16_3;
  assign t_r8_c16_8 = t_r8_c16_4 + p_9_15;
  assign t_r8_c16_9 = t_r8_c16_5 + t_r8_c16_6;
  assign t_r8_c16_10 = t_r8_c16_7 + t_r8_c16_8;
  assign t_r8_c16_11 = t_r8_c16_9 + t_r8_c16_10;
  assign t_r8_c16_12 = t_r8_c16_11 + p_9_17;
  assign out_8_16 = t_r8_c16_12 >> 4;

  assign t_r8_c17_0 = p_7_17 << 1;
  assign t_r8_c17_1 = p_8_16 << 1;
  assign t_r8_c17_2 = p_8_17 << 2;
  assign t_r8_c17_3 = p_8_18 << 1;
  assign t_r8_c17_4 = p_9_17 << 1;
  assign t_r8_c17_5 = t_r8_c17_0 + p_7_16;
  assign t_r8_c17_6 = t_r8_c17_1 + p_7_18;
  assign t_r8_c17_7 = t_r8_c17_2 + t_r8_c17_3;
  assign t_r8_c17_8 = t_r8_c17_4 + p_9_16;
  assign t_r8_c17_9 = t_r8_c17_5 + t_r8_c17_6;
  assign t_r8_c17_10 = t_r8_c17_7 + t_r8_c17_8;
  assign t_r8_c17_11 = t_r8_c17_9 + t_r8_c17_10;
  assign t_r8_c17_12 = t_r8_c17_11 + p_9_18;
  assign out_8_17 = t_r8_c17_12 >> 4;

  assign t_r8_c18_0 = p_7_18 << 1;
  assign t_r8_c18_1 = p_8_17 << 1;
  assign t_r8_c18_2 = p_8_18 << 2;
  assign t_r8_c18_3 = p_8_19 << 1;
  assign t_r8_c18_4 = p_9_18 << 1;
  assign t_r8_c18_5 = t_r8_c18_0 + p_7_17;
  assign t_r8_c18_6 = t_r8_c18_1 + p_7_19;
  assign t_r8_c18_7 = t_r8_c18_2 + t_r8_c18_3;
  assign t_r8_c18_8 = t_r8_c18_4 + p_9_17;
  assign t_r8_c18_9 = t_r8_c18_5 + t_r8_c18_6;
  assign t_r8_c18_10 = t_r8_c18_7 + t_r8_c18_8;
  assign t_r8_c18_11 = t_r8_c18_9 + t_r8_c18_10;
  assign t_r8_c18_12 = t_r8_c18_11 + p_9_19;
  assign out_8_18 = t_r8_c18_12 >> 4;

  assign t_r8_c19_0 = p_7_19 << 1;
  assign t_r8_c19_1 = p_8_18 << 1;
  assign t_r8_c19_2 = p_8_19 << 2;
  assign t_r8_c19_3 = p_8_20 << 1;
  assign t_r8_c19_4 = p_9_19 << 1;
  assign t_r8_c19_5 = t_r8_c19_0 + p_7_18;
  assign t_r8_c19_6 = t_r8_c19_1 + p_7_20;
  assign t_r8_c19_7 = t_r8_c19_2 + t_r8_c19_3;
  assign t_r8_c19_8 = t_r8_c19_4 + p_9_18;
  assign t_r8_c19_9 = t_r8_c19_5 + t_r8_c19_6;
  assign t_r8_c19_10 = t_r8_c19_7 + t_r8_c19_8;
  assign t_r8_c19_11 = t_r8_c19_9 + t_r8_c19_10;
  assign t_r8_c19_12 = t_r8_c19_11 + p_9_20;
  assign out_8_19 = t_r8_c19_12 >> 4;

  assign t_r8_c20_0 = p_7_20 << 1;
  assign t_r8_c20_1 = p_8_19 << 1;
  assign t_r8_c20_2 = p_8_20 << 2;
  assign t_r8_c20_3 = p_8_21 << 1;
  assign t_r8_c20_4 = p_9_20 << 1;
  assign t_r8_c20_5 = t_r8_c20_0 + p_7_19;
  assign t_r8_c20_6 = t_r8_c20_1 + p_7_21;
  assign t_r8_c20_7 = t_r8_c20_2 + t_r8_c20_3;
  assign t_r8_c20_8 = t_r8_c20_4 + p_9_19;
  assign t_r8_c20_9 = t_r8_c20_5 + t_r8_c20_6;
  assign t_r8_c20_10 = t_r8_c20_7 + t_r8_c20_8;
  assign t_r8_c20_11 = t_r8_c20_9 + t_r8_c20_10;
  assign t_r8_c20_12 = t_r8_c20_11 + p_9_21;
  assign out_8_20 = t_r8_c20_12 >> 4;

  assign t_r8_c21_0 = p_7_21 << 1;
  assign t_r8_c21_1 = p_8_20 << 1;
  assign t_r8_c21_2 = p_8_21 << 2;
  assign t_r8_c21_3 = p_8_22 << 1;
  assign t_r8_c21_4 = p_9_21 << 1;
  assign t_r8_c21_5 = t_r8_c21_0 + p_7_20;
  assign t_r8_c21_6 = t_r8_c21_1 + p_7_22;
  assign t_r8_c21_7 = t_r8_c21_2 + t_r8_c21_3;
  assign t_r8_c21_8 = t_r8_c21_4 + p_9_20;
  assign t_r8_c21_9 = t_r8_c21_5 + t_r8_c21_6;
  assign t_r8_c21_10 = t_r8_c21_7 + t_r8_c21_8;
  assign t_r8_c21_11 = t_r8_c21_9 + t_r8_c21_10;
  assign t_r8_c21_12 = t_r8_c21_11 + p_9_22;
  assign out_8_21 = t_r8_c21_12 >> 4;

  assign t_r8_c22_0 = p_7_22 << 1;
  assign t_r8_c22_1 = p_8_21 << 1;
  assign t_r8_c22_2 = p_8_22 << 2;
  assign t_r8_c22_3 = p_8_23 << 1;
  assign t_r8_c22_4 = p_9_22 << 1;
  assign t_r8_c22_5 = t_r8_c22_0 + p_7_21;
  assign t_r8_c22_6 = t_r8_c22_1 + p_7_23;
  assign t_r8_c22_7 = t_r8_c22_2 + t_r8_c22_3;
  assign t_r8_c22_8 = t_r8_c22_4 + p_9_21;
  assign t_r8_c22_9 = t_r8_c22_5 + t_r8_c22_6;
  assign t_r8_c22_10 = t_r8_c22_7 + t_r8_c22_8;
  assign t_r8_c22_11 = t_r8_c22_9 + t_r8_c22_10;
  assign t_r8_c22_12 = t_r8_c22_11 + p_9_23;
  assign out_8_22 = t_r8_c22_12 >> 4;

  assign t_r8_c23_0 = p_7_23 << 1;
  assign t_r8_c23_1 = p_8_22 << 1;
  assign t_r8_c23_2 = p_8_23 << 2;
  assign t_r8_c23_3 = p_8_24 << 1;
  assign t_r8_c23_4 = p_9_23 << 1;
  assign t_r8_c23_5 = t_r8_c23_0 + p_7_22;
  assign t_r8_c23_6 = t_r8_c23_1 + p_7_24;
  assign t_r8_c23_7 = t_r8_c23_2 + t_r8_c23_3;
  assign t_r8_c23_8 = t_r8_c23_4 + p_9_22;
  assign t_r8_c23_9 = t_r8_c23_5 + t_r8_c23_6;
  assign t_r8_c23_10 = t_r8_c23_7 + t_r8_c23_8;
  assign t_r8_c23_11 = t_r8_c23_9 + t_r8_c23_10;
  assign t_r8_c23_12 = t_r8_c23_11 + p_9_24;
  assign out_8_23 = t_r8_c23_12 >> 4;

  assign t_r8_c24_0 = p_7_24 << 1;
  assign t_r8_c24_1 = p_8_23 << 1;
  assign t_r8_c24_2 = p_8_24 << 2;
  assign t_r8_c24_3 = p_8_25 << 1;
  assign t_r8_c24_4 = p_9_24 << 1;
  assign t_r8_c24_5 = t_r8_c24_0 + p_7_23;
  assign t_r8_c24_6 = t_r8_c24_1 + p_7_25;
  assign t_r8_c24_7 = t_r8_c24_2 + t_r8_c24_3;
  assign t_r8_c24_8 = t_r8_c24_4 + p_9_23;
  assign t_r8_c24_9 = t_r8_c24_5 + t_r8_c24_6;
  assign t_r8_c24_10 = t_r8_c24_7 + t_r8_c24_8;
  assign t_r8_c24_11 = t_r8_c24_9 + t_r8_c24_10;
  assign t_r8_c24_12 = t_r8_c24_11 + p_9_25;
  assign out_8_24 = t_r8_c24_12 >> 4;

  assign t_r8_c25_0 = p_7_25 << 1;
  assign t_r8_c25_1 = p_8_24 << 1;
  assign t_r8_c25_2 = p_8_25 << 2;
  assign t_r8_c25_3 = p_8_26 << 1;
  assign t_r8_c25_4 = p_9_25 << 1;
  assign t_r8_c25_5 = t_r8_c25_0 + p_7_24;
  assign t_r8_c25_6 = t_r8_c25_1 + p_7_26;
  assign t_r8_c25_7 = t_r8_c25_2 + t_r8_c25_3;
  assign t_r8_c25_8 = t_r8_c25_4 + p_9_24;
  assign t_r8_c25_9 = t_r8_c25_5 + t_r8_c25_6;
  assign t_r8_c25_10 = t_r8_c25_7 + t_r8_c25_8;
  assign t_r8_c25_11 = t_r8_c25_9 + t_r8_c25_10;
  assign t_r8_c25_12 = t_r8_c25_11 + p_9_26;
  assign out_8_25 = t_r8_c25_12 >> 4;

  assign t_r8_c26_0 = p_7_26 << 1;
  assign t_r8_c26_1 = p_8_25 << 1;
  assign t_r8_c26_2 = p_8_26 << 2;
  assign t_r8_c26_3 = p_8_27 << 1;
  assign t_r8_c26_4 = p_9_26 << 1;
  assign t_r8_c26_5 = t_r8_c26_0 + p_7_25;
  assign t_r8_c26_6 = t_r8_c26_1 + p_7_27;
  assign t_r8_c26_7 = t_r8_c26_2 + t_r8_c26_3;
  assign t_r8_c26_8 = t_r8_c26_4 + p_9_25;
  assign t_r8_c26_9 = t_r8_c26_5 + t_r8_c26_6;
  assign t_r8_c26_10 = t_r8_c26_7 + t_r8_c26_8;
  assign t_r8_c26_11 = t_r8_c26_9 + t_r8_c26_10;
  assign t_r8_c26_12 = t_r8_c26_11 + p_9_27;
  assign out_8_26 = t_r8_c26_12 >> 4;

  assign t_r8_c27_0 = p_7_27 << 1;
  assign t_r8_c27_1 = p_8_26 << 1;
  assign t_r8_c27_2 = p_8_27 << 2;
  assign t_r8_c27_3 = p_8_28 << 1;
  assign t_r8_c27_4 = p_9_27 << 1;
  assign t_r8_c27_5 = t_r8_c27_0 + p_7_26;
  assign t_r8_c27_6 = t_r8_c27_1 + p_7_28;
  assign t_r8_c27_7 = t_r8_c27_2 + t_r8_c27_3;
  assign t_r8_c27_8 = t_r8_c27_4 + p_9_26;
  assign t_r8_c27_9 = t_r8_c27_5 + t_r8_c27_6;
  assign t_r8_c27_10 = t_r8_c27_7 + t_r8_c27_8;
  assign t_r8_c27_11 = t_r8_c27_9 + t_r8_c27_10;
  assign t_r8_c27_12 = t_r8_c27_11 + p_9_28;
  assign out_8_27 = t_r8_c27_12 >> 4;

  assign t_r8_c28_0 = p_7_28 << 1;
  assign t_r8_c28_1 = p_8_27 << 1;
  assign t_r8_c28_2 = p_8_28 << 2;
  assign t_r8_c28_3 = p_8_29 << 1;
  assign t_r8_c28_4 = p_9_28 << 1;
  assign t_r8_c28_5 = t_r8_c28_0 + p_7_27;
  assign t_r8_c28_6 = t_r8_c28_1 + p_7_29;
  assign t_r8_c28_7 = t_r8_c28_2 + t_r8_c28_3;
  assign t_r8_c28_8 = t_r8_c28_4 + p_9_27;
  assign t_r8_c28_9 = t_r8_c28_5 + t_r8_c28_6;
  assign t_r8_c28_10 = t_r8_c28_7 + t_r8_c28_8;
  assign t_r8_c28_11 = t_r8_c28_9 + t_r8_c28_10;
  assign t_r8_c28_12 = t_r8_c28_11 + p_9_29;
  assign out_8_28 = t_r8_c28_12 >> 4;

  assign t_r8_c29_0 = p_7_29 << 1;
  assign t_r8_c29_1 = p_8_28 << 1;
  assign t_r8_c29_2 = p_8_29 << 2;
  assign t_r8_c29_3 = p_8_30 << 1;
  assign t_r8_c29_4 = p_9_29 << 1;
  assign t_r8_c29_5 = t_r8_c29_0 + p_7_28;
  assign t_r8_c29_6 = t_r8_c29_1 + p_7_30;
  assign t_r8_c29_7 = t_r8_c29_2 + t_r8_c29_3;
  assign t_r8_c29_8 = t_r8_c29_4 + p_9_28;
  assign t_r8_c29_9 = t_r8_c29_5 + t_r8_c29_6;
  assign t_r8_c29_10 = t_r8_c29_7 + t_r8_c29_8;
  assign t_r8_c29_11 = t_r8_c29_9 + t_r8_c29_10;
  assign t_r8_c29_12 = t_r8_c29_11 + p_9_30;
  assign out_8_29 = t_r8_c29_12 >> 4;

  assign t_r8_c30_0 = p_7_30 << 1;
  assign t_r8_c30_1 = p_8_29 << 1;
  assign t_r8_c30_2 = p_8_30 << 2;
  assign t_r8_c30_3 = p_8_31 << 1;
  assign t_r8_c30_4 = p_9_30 << 1;
  assign t_r8_c30_5 = t_r8_c30_0 + p_7_29;
  assign t_r8_c30_6 = t_r8_c30_1 + p_7_31;
  assign t_r8_c30_7 = t_r8_c30_2 + t_r8_c30_3;
  assign t_r8_c30_8 = t_r8_c30_4 + p_9_29;
  assign t_r8_c30_9 = t_r8_c30_5 + t_r8_c30_6;
  assign t_r8_c30_10 = t_r8_c30_7 + t_r8_c30_8;
  assign t_r8_c30_11 = t_r8_c30_9 + t_r8_c30_10;
  assign t_r8_c30_12 = t_r8_c30_11 + p_9_31;
  assign out_8_30 = t_r8_c30_12 >> 4;

  assign t_r8_c31_0 = p_7_31 << 1;
  assign t_r8_c31_1 = p_8_30 << 1;
  assign t_r8_c31_2 = p_8_31 << 2;
  assign t_r8_c31_3 = p_8_32 << 1;
  assign t_r8_c31_4 = p_9_31 << 1;
  assign t_r8_c31_5 = t_r8_c31_0 + p_7_30;
  assign t_r8_c31_6 = t_r8_c31_1 + p_7_32;
  assign t_r8_c31_7 = t_r8_c31_2 + t_r8_c31_3;
  assign t_r8_c31_8 = t_r8_c31_4 + p_9_30;
  assign t_r8_c31_9 = t_r8_c31_5 + t_r8_c31_6;
  assign t_r8_c31_10 = t_r8_c31_7 + t_r8_c31_8;
  assign t_r8_c31_11 = t_r8_c31_9 + t_r8_c31_10;
  assign t_r8_c31_12 = t_r8_c31_11 + p_9_32;
  assign out_8_31 = t_r8_c31_12 >> 4;

  assign t_r8_c32_0 = p_7_32 << 1;
  assign t_r8_c32_1 = p_8_31 << 1;
  assign t_r8_c32_2 = p_8_32 << 2;
  assign t_r8_c32_3 = p_8_33 << 1;
  assign t_r8_c32_4 = p_9_32 << 1;
  assign t_r8_c32_5 = t_r8_c32_0 + p_7_31;
  assign t_r8_c32_6 = t_r8_c32_1 + p_7_33;
  assign t_r8_c32_7 = t_r8_c32_2 + t_r8_c32_3;
  assign t_r8_c32_8 = t_r8_c32_4 + p_9_31;
  assign t_r8_c32_9 = t_r8_c32_5 + t_r8_c32_6;
  assign t_r8_c32_10 = t_r8_c32_7 + t_r8_c32_8;
  assign t_r8_c32_11 = t_r8_c32_9 + t_r8_c32_10;
  assign t_r8_c32_12 = t_r8_c32_11 + p_9_33;
  assign out_8_32 = t_r8_c32_12 >> 4;

  assign t_r8_c33_0 = p_7_33 << 1;
  assign t_r8_c33_1 = p_8_32 << 1;
  assign t_r8_c33_2 = p_8_33 << 2;
  assign t_r8_c33_3 = p_8_34 << 1;
  assign t_r8_c33_4 = p_9_33 << 1;
  assign t_r8_c33_5 = t_r8_c33_0 + p_7_32;
  assign t_r8_c33_6 = t_r8_c33_1 + p_7_34;
  assign t_r8_c33_7 = t_r8_c33_2 + t_r8_c33_3;
  assign t_r8_c33_8 = t_r8_c33_4 + p_9_32;
  assign t_r8_c33_9 = t_r8_c33_5 + t_r8_c33_6;
  assign t_r8_c33_10 = t_r8_c33_7 + t_r8_c33_8;
  assign t_r8_c33_11 = t_r8_c33_9 + t_r8_c33_10;
  assign t_r8_c33_12 = t_r8_c33_11 + p_9_34;
  assign out_8_33 = t_r8_c33_12 >> 4;

  assign t_r8_c34_0 = p_7_34 << 1;
  assign t_r8_c34_1 = p_8_33 << 1;
  assign t_r8_c34_2 = p_8_34 << 2;
  assign t_r8_c34_3 = p_8_35 << 1;
  assign t_r8_c34_4 = p_9_34 << 1;
  assign t_r8_c34_5 = t_r8_c34_0 + p_7_33;
  assign t_r8_c34_6 = t_r8_c34_1 + p_7_35;
  assign t_r8_c34_7 = t_r8_c34_2 + t_r8_c34_3;
  assign t_r8_c34_8 = t_r8_c34_4 + p_9_33;
  assign t_r8_c34_9 = t_r8_c34_5 + t_r8_c34_6;
  assign t_r8_c34_10 = t_r8_c34_7 + t_r8_c34_8;
  assign t_r8_c34_11 = t_r8_c34_9 + t_r8_c34_10;
  assign t_r8_c34_12 = t_r8_c34_11 + p_9_35;
  assign out_8_34 = t_r8_c34_12 >> 4;

  assign t_r8_c35_0 = p_7_35 << 1;
  assign t_r8_c35_1 = p_8_34 << 1;
  assign t_r8_c35_2 = p_8_35 << 2;
  assign t_r8_c35_3 = p_8_36 << 1;
  assign t_r8_c35_4 = p_9_35 << 1;
  assign t_r8_c35_5 = t_r8_c35_0 + p_7_34;
  assign t_r8_c35_6 = t_r8_c35_1 + p_7_36;
  assign t_r8_c35_7 = t_r8_c35_2 + t_r8_c35_3;
  assign t_r8_c35_8 = t_r8_c35_4 + p_9_34;
  assign t_r8_c35_9 = t_r8_c35_5 + t_r8_c35_6;
  assign t_r8_c35_10 = t_r8_c35_7 + t_r8_c35_8;
  assign t_r8_c35_11 = t_r8_c35_9 + t_r8_c35_10;
  assign t_r8_c35_12 = t_r8_c35_11 + p_9_36;
  assign out_8_35 = t_r8_c35_12 >> 4;

  assign t_r8_c36_0 = p_7_36 << 1;
  assign t_r8_c36_1 = p_8_35 << 1;
  assign t_r8_c36_2 = p_8_36 << 2;
  assign t_r8_c36_3 = p_8_37 << 1;
  assign t_r8_c36_4 = p_9_36 << 1;
  assign t_r8_c36_5 = t_r8_c36_0 + p_7_35;
  assign t_r8_c36_6 = t_r8_c36_1 + p_7_37;
  assign t_r8_c36_7 = t_r8_c36_2 + t_r8_c36_3;
  assign t_r8_c36_8 = t_r8_c36_4 + p_9_35;
  assign t_r8_c36_9 = t_r8_c36_5 + t_r8_c36_6;
  assign t_r8_c36_10 = t_r8_c36_7 + t_r8_c36_8;
  assign t_r8_c36_11 = t_r8_c36_9 + t_r8_c36_10;
  assign t_r8_c36_12 = t_r8_c36_11 + p_9_37;
  assign out_8_36 = t_r8_c36_12 >> 4;

  assign t_r8_c37_0 = p_7_37 << 1;
  assign t_r8_c37_1 = p_8_36 << 1;
  assign t_r8_c37_2 = p_8_37 << 2;
  assign t_r8_c37_3 = p_8_38 << 1;
  assign t_r8_c37_4 = p_9_37 << 1;
  assign t_r8_c37_5 = t_r8_c37_0 + p_7_36;
  assign t_r8_c37_6 = t_r8_c37_1 + p_7_38;
  assign t_r8_c37_7 = t_r8_c37_2 + t_r8_c37_3;
  assign t_r8_c37_8 = t_r8_c37_4 + p_9_36;
  assign t_r8_c37_9 = t_r8_c37_5 + t_r8_c37_6;
  assign t_r8_c37_10 = t_r8_c37_7 + t_r8_c37_8;
  assign t_r8_c37_11 = t_r8_c37_9 + t_r8_c37_10;
  assign t_r8_c37_12 = t_r8_c37_11 + p_9_38;
  assign out_8_37 = t_r8_c37_12 >> 4;

  assign t_r8_c38_0 = p_7_38 << 1;
  assign t_r8_c38_1 = p_8_37 << 1;
  assign t_r8_c38_2 = p_8_38 << 2;
  assign t_r8_c38_3 = p_8_39 << 1;
  assign t_r8_c38_4 = p_9_38 << 1;
  assign t_r8_c38_5 = t_r8_c38_0 + p_7_37;
  assign t_r8_c38_6 = t_r8_c38_1 + p_7_39;
  assign t_r8_c38_7 = t_r8_c38_2 + t_r8_c38_3;
  assign t_r8_c38_8 = t_r8_c38_4 + p_9_37;
  assign t_r8_c38_9 = t_r8_c38_5 + t_r8_c38_6;
  assign t_r8_c38_10 = t_r8_c38_7 + t_r8_c38_8;
  assign t_r8_c38_11 = t_r8_c38_9 + t_r8_c38_10;
  assign t_r8_c38_12 = t_r8_c38_11 + p_9_39;
  assign out_8_38 = t_r8_c38_12 >> 4;

  assign t_r8_c39_0 = p_7_39 << 1;
  assign t_r8_c39_1 = p_8_38 << 1;
  assign t_r8_c39_2 = p_8_39 << 2;
  assign t_r8_c39_3 = p_8_40 << 1;
  assign t_r8_c39_4 = p_9_39 << 1;
  assign t_r8_c39_5 = t_r8_c39_0 + p_7_38;
  assign t_r8_c39_6 = t_r8_c39_1 + p_7_40;
  assign t_r8_c39_7 = t_r8_c39_2 + t_r8_c39_3;
  assign t_r8_c39_8 = t_r8_c39_4 + p_9_38;
  assign t_r8_c39_9 = t_r8_c39_5 + t_r8_c39_6;
  assign t_r8_c39_10 = t_r8_c39_7 + t_r8_c39_8;
  assign t_r8_c39_11 = t_r8_c39_9 + t_r8_c39_10;
  assign t_r8_c39_12 = t_r8_c39_11 + p_9_40;
  assign out_8_39 = t_r8_c39_12 >> 4;

  assign t_r8_c40_0 = p_7_40 << 1;
  assign t_r8_c40_1 = p_8_39 << 1;
  assign t_r8_c40_2 = p_8_40 << 2;
  assign t_r8_c40_3 = p_8_41 << 1;
  assign t_r8_c40_4 = p_9_40 << 1;
  assign t_r8_c40_5 = t_r8_c40_0 + p_7_39;
  assign t_r8_c40_6 = t_r8_c40_1 + p_7_41;
  assign t_r8_c40_7 = t_r8_c40_2 + t_r8_c40_3;
  assign t_r8_c40_8 = t_r8_c40_4 + p_9_39;
  assign t_r8_c40_9 = t_r8_c40_5 + t_r8_c40_6;
  assign t_r8_c40_10 = t_r8_c40_7 + t_r8_c40_8;
  assign t_r8_c40_11 = t_r8_c40_9 + t_r8_c40_10;
  assign t_r8_c40_12 = t_r8_c40_11 + p_9_41;
  assign out_8_40 = t_r8_c40_12 >> 4;

  assign t_r8_c41_0 = p_7_41 << 1;
  assign t_r8_c41_1 = p_8_40 << 1;
  assign t_r8_c41_2 = p_8_41 << 2;
  assign t_r8_c41_3 = p_8_42 << 1;
  assign t_r8_c41_4 = p_9_41 << 1;
  assign t_r8_c41_5 = t_r8_c41_0 + p_7_40;
  assign t_r8_c41_6 = t_r8_c41_1 + p_7_42;
  assign t_r8_c41_7 = t_r8_c41_2 + t_r8_c41_3;
  assign t_r8_c41_8 = t_r8_c41_4 + p_9_40;
  assign t_r8_c41_9 = t_r8_c41_5 + t_r8_c41_6;
  assign t_r8_c41_10 = t_r8_c41_7 + t_r8_c41_8;
  assign t_r8_c41_11 = t_r8_c41_9 + t_r8_c41_10;
  assign t_r8_c41_12 = t_r8_c41_11 + p_9_42;
  assign out_8_41 = t_r8_c41_12 >> 4;

  assign t_r8_c42_0 = p_7_42 << 1;
  assign t_r8_c42_1 = p_8_41 << 1;
  assign t_r8_c42_2 = p_8_42 << 2;
  assign t_r8_c42_3 = p_8_43 << 1;
  assign t_r8_c42_4 = p_9_42 << 1;
  assign t_r8_c42_5 = t_r8_c42_0 + p_7_41;
  assign t_r8_c42_6 = t_r8_c42_1 + p_7_43;
  assign t_r8_c42_7 = t_r8_c42_2 + t_r8_c42_3;
  assign t_r8_c42_8 = t_r8_c42_4 + p_9_41;
  assign t_r8_c42_9 = t_r8_c42_5 + t_r8_c42_6;
  assign t_r8_c42_10 = t_r8_c42_7 + t_r8_c42_8;
  assign t_r8_c42_11 = t_r8_c42_9 + t_r8_c42_10;
  assign t_r8_c42_12 = t_r8_c42_11 + p_9_43;
  assign out_8_42 = t_r8_c42_12 >> 4;

  assign t_r8_c43_0 = p_7_43 << 1;
  assign t_r8_c43_1 = p_8_42 << 1;
  assign t_r8_c43_2 = p_8_43 << 2;
  assign t_r8_c43_3 = p_8_44 << 1;
  assign t_r8_c43_4 = p_9_43 << 1;
  assign t_r8_c43_5 = t_r8_c43_0 + p_7_42;
  assign t_r8_c43_6 = t_r8_c43_1 + p_7_44;
  assign t_r8_c43_7 = t_r8_c43_2 + t_r8_c43_3;
  assign t_r8_c43_8 = t_r8_c43_4 + p_9_42;
  assign t_r8_c43_9 = t_r8_c43_5 + t_r8_c43_6;
  assign t_r8_c43_10 = t_r8_c43_7 + t_r8_c43_8;
  assign t_r8_c43_11 = t_r8_c43_9 + t_r8_c43_10;
  assign t_r8_c43_12 = t_r8_c43_11 + p_9_44;
  assign out_8_43 = t_r8_c43_12 >> 4;

  assign t_r8_c44_0 = p_7_44 << 1;
  assign t_r8_c44_1 = p_8_43 << 1;
  assign t_r8_c44_2 = p_8_44 << 2;
  assign t_r8_c44_3 = p_8_45 << 1;
  assign t_r8_c44_4 = p_9_44 << 1;
  assign t_r8_c44_5 = t_r8_c44_0 + p_7_43;
  assign t_r8_c44_6 = t_r8_c44_1 + p_7_45;
  assign t_r8_c44_7 = t_r8_c44_2 + t_r8_c44_3;
  assign t_r8_c44_8 = t_r8_c44_4 + p_9_43;
  assign t_r8_c44_9 = t_r8_c44_5 + t_r8_c44_6;
  assign t_r8_c44_10 = t_r8_c44_7 + t_r8_c44_8;
  assign t_r8_c44_11 = t_r8_c44_9 + t_r8_c44_10;
  assign t_r8_c44_12 = t_r8_c44_11 + p_9_45;
  assign out_8_44 = t_r8_c44_12 >> 4;

  assign t_r8_c45_0 = p_7_45 << 1;
  assign t_r8_c45_1 = p_8_44 << 1;
  assign t_r8_c45_2 = p_8_45 << 2;
  assign t_r8_c45_3 = p_8_46 << 1;
  assign t_r8_c45_4 = p_9_45 << 1;
  assign t_r8_c45_5 = t_r8_c45_0 + p_7_44;
  assign t_r8_c45_6 = t_r8_c45_1 + p_7_46;
  assign t_r8_c45_7 = t_r8_c45_2 + t_r8_c45_3;
  assign t_r8_c45_8 = t_r8_c45_4 + p_9_44;
  assign t_r8_c45_9 = t_r8_c45_5 + t_r8_c45_6;
  assign t_r8_c45_10 = t_r8_c45_7 + t_r8_c45_8;
  assign t_r8_c45_11 = t_r8_c45_9 + t_r8_c45_10;
  assign t_r8_c45_12 = t_r8_c45_11 + p_9_46;
  assign out_8_45 = t_r8_c45_12 >> 4;

  assign t_r8_c46_0 = p_7_46 << 1;
  assign t_r8_c46_1 = p_8_45 << 1;
  assign t_r8_c46_2 = p_8_46 << 2;
  assign t_r8_c46_3 = p_8_47 << 1;
  assign t_r8_c46_4 = p_9_46 << 1;
  assign t_r8_c46_5 = t_r8_c46_0 + p_7_45;
  assign t_r8_c46_6 = t_r8_c46_1 + p_7_47;
  assign t_r8_c46_7 = t_r8_c46_2 + t_r8_c46_3;
  assign t_r8_c46_8 = t_r8_c46_4 + p_9_45;
  assign t_r8_c46_9 = t_r8_c46_5 + t_r8_c46_6;
  assign t_r8_c46_10 = t_r8_c46_7 + t_r8_c46_8;
  assign t_r8_c46_11 = t_r8_c46_9 + t_r8_c46_10;
  assign t_r8_c46_12 = t_r8_c46_11 + p_9_47;
  assign out_8_46 = t_r8_c46_12 >> 4;

  assign t_r8_c47_0 = p_7_47 << 1;
  assign t_r8_c47_1 = p_8_46 << 1;
  assign t_r8_c47_2 = p_8_47 << 2;
  assign t_r8_c47_3 = p_8_48 << 1;
  assign t_r8_c47_4 = p_9_47 << 1;
  assign t_r8_c47_5 = t_r8_c47_0 + p_7_46;
  assign t_r8_c47_6 = t_r8_c47_1 + p_7_48;
  assign t_r8_c47_7 = t_r8_c47_2 + t_r8_c47_3;
  assign t_r8_c47_8 = t_r8_c47_4 + p_9_46;
  assign t_r8_c47_9 = t_r8_c47_5 + t_r8_c47_6;
  assign t_r8_c47_10 = t_r8_c47_7 + t_r8_c47_8;
  assign t_r8_c47_11 = t_r8_c47_9 + t_r8_c47_10;
  assign t_r8_c47_12 = t_r8_c47_11 + p_9_48;
  assign out_8_47 = t_r8_c47_12 >> 4;

  assign t_r8_c48_0 = p_7_48 << 1;
  assign t_r8_c48_1 = p_8_47 << 1;
  assign t_r8_c48_2 = p_8_48 << 2;
  assign t_r8_c48_3 = p_8_49 << 1;
  assign t_r8_c48_4 = p_9_48 << 1;
  assign t_r8_c48_5 = t_r8_c48_0 + p_7_47;
  assign t_r8_c48_6 = t_r8_c48_1 + p_7_49;
  assign t_r8_c48_7 = t_r8_c48_2 + t_r8_c48_3;
  assign t_r8_c48_8 = t_r8_c48_4 + p_9_47;
  assign t_r8_c48_9 = t_r8_c48_5 + t_r8_c48_6;
  assign t_r8_c48_10 = t_r8_c48_7 + t_r8_c48_8;
  assign t_r8_c48_11 = t_r8_c48_9 + t_r8_c48_10;
  assign t_r8_c48_12 = t_r8_c48_11 + p_9_49;
  assign out_8_48 = t_r8_c48_12 >> 4;

  assign t_r8_c49_0 = p_7_49 << 1;
  assign t_r8_c49_1 = p_8_48 << 1;
  assign t_r8_c49_2 = p_8_49 << 2;
  assign t_r8_c49_3 = p_8_50 << 1;
  assign t_r8_c49_4 = p_9_49 << 1;
  assign t_r8_c49_5 = t_r8_c49_0 + p_7_48;
  assign t_r8_c49_6 = t_r8_c49_1 + p_7_50;
  assign t_r8_c49_7 = t_r8_c49_2 + t_r8_c49_3;
  assign t_r8_c49_8 = t_r8_c49_4 + p_9_48;
  assign t_r8_c49_9 = t_r8_c49_5 + t_r8_c49_6;
  assign t_r8_c49_10 = t_r8_c49_7 + t_r8_c49_8;
  assign t_r8_c49_11 = t_r8_c49_9 + t_r8_c49_10;
  assign t_r8_c49_12 = t_r8_c49_11 + p_9_50;
  assign out_8_49 = t_r8_c49_12 >> 4;

  assign t_r8_c50_0 = p_7_50 << 1;
  assign t_r8_c50_1 = p_8_49 << 1;
  assign t_r8_c50_2 = p_8_50 << 2;
  assign t_r8_c50_3 = p_8_51 << 1;
  assign t_r8_c50_4 = p_9_50 << 1;
  assign t_r8_c50_5 = t_r8_c50_0 + p_7_49;
  assign t_r8_c50_6 = t_r8_c50_1 + p_7_51;
  assign t_r8_c50_7 = t_r8_c50_2 + t_r8_c50_3;
  assign t_r8_c50_8 = t_r8_c50_4 + p_9_49;
  assign t_r8_c50_9 = t_r8_c50_5 + t_r8_c50_6;
  assign t_r8_c50_10 = t_r8_c50_7 + t_r8_c50_8;
  assign t_r8_c50_11 = t_r8_c50_9 + t_r8_c50_10;
  assign t_r8_c50_12 = t_r8_c50_11 + p_9_51;
  assign out_8_50 = t_r8_c50_12 >> 4;

  assign t_r8_c51_0 = p_7_51 << 1;
  assign t_r8_c51_1 = p_8_50 << 1;
  assign t_r8_c51_2 = p_8_51 << 2;
  assign t_r8_c51_3 = p_8_52 << 1;
  assign t_r8_c51_4 = p_9_51 << 1;
  assign t_r8_c51_5 = t_r8_c51_0 + p_7_50;
  assign t_r8_c51_6 = t_r8_c51_1 + p_7_52;
  assign t_r8_c51_7 = t_r8_c51_2 + t_r8_c51_3;
  assign t_r8_c51_8 = t_r8_c51_4 + p_9_50;
  assign t_r8_c51_9 = t_r8_c51_5 + t_r8_c51_6;
  assign t_r8_c51_10 = t_r8_c51_7 + t_r8_c51_8;
  assign t_r8_c51_11 = t_r8_c51_9 + t_r8_c51_10;
  assign t_r8_c51_12 = t_r8_c51_11 + p_9_52;
  assign out_8_51 = t_r8_c51_12 >> 4;

  assign t_r8_c52_0 = p_7_52 << 1;
  assign t_r8_c52_1 = p_8_51 << 1;
  assign t_r8_c52_2 = p_8_52 << 2;
  assign t_r8_c52_3 = p_8_53 << 1;
  assign t_r8_c52_4 = p_9_52 << 1;
  assign t_r8_c52_5 = t_r8_c52_0 + p_7_51;
  assign t_r8_c52_6 = t_r8_c52_1 + p_7_53;
  assign t_r8_c52_7 = t_r8_c52_2 + t_r8_c52_3;
  assign t_r8_c52_8 = t_r8_c52_4 + p_9_51;
  assign t_r8_c52_9 = t_r8_c52_5 + t_r8_c52_6;
  assign t_r8_c52_10 = t_r8_c52_7 + t_r8_c52_8;
  assign t_r8_c52_11 = t_r8_c52_9 + t_r8_c52_10;
  assign t_r8_c52_12 = t_r8_c52_11 + p_9_53;
  assign out_8_52 = t_r8_c52_12 >> 4;

  assign t_r8_c53_0 = p_7_53 << 1;
  assign t_r8_c53_1 = p_8_52 << 1;
  assign t_r8_c53_2 = p_8_53 << 2;
  assign t_r8_c53_3 = p_8_54 << 1;
  assign t_r8_c53_4 = p_9_53 << 1;
  assign t_r8_c53_5 = t_r8_c53_0 + p_7_52;
  assign t_r8_c53_6 = t_r8_c53_1 + p_7_54;
  assign t_r8_c53_7 = t_r8_c53_2 + t_r8_c53_3;
  assign t_r8_c53_8 = t_r8_c53_4 + p_9_52;
  assign t_r8_c53_9 = t_r8_c53_5 + t_r8_c53_6;
  assign t_r8_c53_10 = t_r8_c53_7 + t_r8_c53_8;
  assign t_r8_c53_11 = t_r8_c53_9 + t_r8_c53_10;
  assign t_r8_c53_12 = t_r8_c53_11 + p_9_54;
  assign out_8_53 = t_r8_c53_12 >> 4;

  assign t_r8_c54_0 = p_7_54 << 1;
  assign t_r8_c54_1 = p_8_53 << 1;
  assign t_r8_c54_2 = p_8_54 << 2;
  assign t_r8_c54_3 = p_8_55 << 1;
  assign t_r8_c54_4 = p_9_54 << 1;
  assign t_r8_c54_5 = t_r8_c54_0 + p_7_53;
  assign t_r8_c54_6 = t_r8_c54_1 + p_7_55;
  assign t_r8_c54_7 = t_r8_c54_2 + t_r8_c54_3;
  assign t_r8_c54_8 = t_r8_c54_4 + p_9_53;
  assign t_r8_c54_9 = t_r8_c54_5 + t_r8_c54_6;
  assign t_r8_c54_10 = t_r8_c54_7 + t_r8_c54_8;
  assign t_r8_c54_11 = t_r8_c54_9 + t_r8_c54_10;
  assign t_r8_c54_12 = t_r8_c54_11 + p_9_55;
  assign out_8_54 = t_r8_c54_12 >> 4;

  assign t_r8_c55_0 = p_7_55 << 1;
  assign t_r8_c55_1 = p_8_54 << 1;
  assign t_r8_c55_2 = p_8_55 << 2;
  assign t_r8_c55_3 = p_8_56 << 1;
  assign t_r8_c55_4 = p_9_55 << 1;
  assign t_r8_c55_5 = t_r8_c55_0 + p_7_54;
  assign t_r8_c55_6 = t_r8_c55_1 + p_7_56;
  assign t_r8_c55_7 = t_r8_c55_2 + t_r8_c55_3;
  assign t_r8_c55_8 = t_r8_c55_4 + p_9_54;
  assign t_r8_c55_9 = t_r8_c55_5 + t_r8_c55_6;
  assign t_r8_c55_10 = t_r8_c55_7 + t_r8_c55_8;
  assign t_r8_c55_11 = t_r8_c55_9 + t_r8_c55_10;
  assign t_r8_c55_12 = t_r8_c55_11 + p_9_56;
  assign out_8_55 = t_r8_c55_12 >> 4;

  assign t_r8_c56_0 = p_7_56 << 1;
  assign t_r8_c56_1 = p_8_55 << 1;
  assign t_r8_c56_2 = p_8_56 << 2;
  assign t_r8_c56_3 = p_8_57 << 1;
  assign t_r8_c56_4 = p_9_56 << 1;
  assign t_r8_c56_5 = t_r8_c56_0 + p_7_55;
  assign t_r8_c56_6 = t_r8_c56_1 + p_7_57;
  assign t_r8_c56_7 = t_r8_c56_2 + t_r8_c56_3;
  assign t_r8_c56_8 = t_r8_c56_4 + p_9_55;
  assign t_r8_c56_9 = t_r8_c56_5 + t_r8_c56_6;
  assign t_r8_c56_10 = t_r8_c56_7 + t_r8_c56_8;
  assign t_r8_c56_11 = t_r8_c56_9 + t_r8_c56_10;
  assign t_r8_c56_12 = t_r8_c56_11 + p_9_57;
  assign out_8_56 = t_r8_c56_12 >> 4;

  assign t_r8_c57_0 = p_7_57 << 1;
  assign t_r8_c57_1 = p_8_56 << 1;
  assign t_r8_c57_2 = p_8_57 << 2;
  assign t_r8_c57_3 = p_8_58 << 1;
  assign t_r8_c57_4 = p_9_57 << 1;
  assign t_r8_c57_5 = t_r8_c57_0 + p_7_56;
  assign t_r8_c57_6 = t_r8_c57_1 + p_7_58;
  assign t_r8_c57_7 = t_r8_c57_2 + t_r8_c57_3;
  assign t_r8_c57_8 = t_r8_c57_4 + p_9_56;
  assign t_r8_c57_9 = t_r8_c57_5 + t_r8_c57_6;
  assign t_r8_c57_10 = t_r8_c57_7 + t_r8_c57_8;
  assign t_r8_c57_11 = t_r8_c57_9 + t_r8_c57_10;
  assign t_r8_c57_12 = t_r8_c57_11 + p_9_58;
  assign out_8_57 = t_r8_c57_12 >> 4;

  assign t_r8_c58_0 = p_7_58 << 1;
  assign t_r8_c58_1 = p_8_57 << 1;
  assign t_r8_c58_2 = p_8_58 << 2;
  assign t_r8_c58_3 = p_8_59 << 1;
  assign t_r8_c58_4 = p_9_58 << 1;
  assign t_r8_c58_5 = t_r8_c58_0 + p_7_57;
  assign t_r8_c58_6 = t_r8_c58_1 + p_7_59;
  assign t_r8_c58_7 = t_r8_c58_2 + t_r8_c58_3;
  assign t_r8_c58_8 = t_r8_c58_4 + p_9_57;
  assign t_r8_c58_9 = t_r8_c58_5 + t_r8_c58_6;
  assign t_r8_c58_10 = t_r8_c58_7 + t_r8_c58_8;
  assign t_r8_c58_11 = t_r8_c58_9 + t_r8_c58_10;
  assign t_r8_c58_12 = t_r8_c58_11 + p_9_59;
  assign out_8_58 = t_r8_c58_12 >> 4;

  assign t_r8_c59_0 = p_7_59 << 1;
  assign t_r8_c59_1 = p_8_58 << 1;
  assign t_r8_c59_2 = p_8_59 << 2;
  assign t_r8_c59_3 = p_8_60 << 1;
  assign t_r8_c59_4 = p_9_59 << 1;
  assign t_r8_c59_5 = t_r8_c59_0 + p_7_58;
  assign t_r8_c59_6 = t_r8_c59_1 + p_7_60;
  assign t_r8_c59_7 = t_r8_c59_2 + t_r8_c59_3;
  assign t_r8_c59_8 = t_r8_c59_4 + p_9_58;
  assign t_r8_c59_9 = t_r8_c59_5 + t_r8_c59_6;
  assign t_r8_c59_10 = t_r8_c59_7 + t_r8_c59_8;
  assign t_r8_c59_11 = t_r8_c59_9 + t_r8_c59_10;
  assign t_r8_c59_12 = t_r8_c59_11 + p_9_60;
  assign out_8_59 = t_r8_c59_12 >> 4;

  assign t_r8_c60_0 = p_7_60 << 1;
  assign t_r8_c60_1 = p_8_59 << 1;
  assign t_r8_c60_2 = p_8_60 << 2;
  assign t_r8_c60_3 = p_8_61 << 1;
  assign t_r8_c60_4 = p_9_60 << 1;
  assign t_r8_c60_5 = t_r8_c60_0 + p_7_59;
  assign t_r8_c60_6 = t_r8_c60_1 + p_7_61;
  assign t_r8_c60_7 = t_r8_c60_2 + t_r8_c60_3;
  assign t_r8_c60_8 = t_r8_c60_4 + p_9_59;
  assign t_r8_c60_9 = t_r8_c60_5 + t_r8_c60_6;
  assign t_r8_c60_10 = t_r8_c60_7 + t_r8_c60_8;
  assign t_r8_c60_11 = t_r8_c60_9 + t_r8_c60_10;
  assign t_r8_c60_12 = t_r8_c60_11 + p_9_61;
  assign out_8_60 = t_r8_c60_12 >> 4;

  assign t_r8_c61_0 = p_7_61 << 1;
  assign t_r8_c61_1 = p_8_60 << 1;
  assign t_r8_c61_2 = p_8_61 << 2;
  assign t_r8_c61_3 = p_8_62 << 1;
  assign t_r8_c61_4 = p_9_61 << 1;
  assign t_r8_c61_5 = t_r8_c61_0 + p_7_60;
  assign t_r8_c61_6 = t_r8_c61_1 + p_7_62;
  assign t_r8_c61_7 = t_r8_c61_2 + t_r8_c61_3;
  assign t_r8_c61_8 = t_r8_c61_4 + p_9_60;
  assign t_r8_c61_9 = t_r8_c61_5 + t_r8_c61_6;
  assign t_r8_c61_10 = t_r8_c61_7 + t_r8_c61_8;
  assign t_r8_c61_11 = t_r8_c61_9 + t_r8_c61_10;
  assign t_r8_c61_12 = t_r8_c61_11 + p_9_62;
  assign out_8_61 = t_r8_c61_12 >> 4;

  assign t_r8_c62_0 = p_7_62 << 1;
  assign t_r8_c62_1 = p_8_61 << 1;
  assign t_r8_c62_2 = p_8_62 << 2;
  assign t_r8_c62_3 = p_8_63 << 1;
  assign t_r8_c62_4 = p_9_62 << 1;
  assign t_r8_c62_5 = t_r8_c62_0 + p_7_61;
  assign t_r8_c62_6 = t_r8_c62_1 + p_7_63;
  assign t_r8_c62_7 = t_r8_c62_2 + t_r8_c62_3;
  assign t_r8_c62_8 = t_r8_c62_4 + p_9_61;
  assign t_r8_c62_9 = t_r8_c62_5 + t_r8_c62_6;
  assign t_r8_c62_10 = t_r8_c62_7 + t_r8_c62_8;
  assign t_r8_c62_11 = t_r8_c62_9 + t_r8_c62_10;
  assign t_r8_c62_12 = t_r8_c62_11 + p_9_63;
  assign out_8_62 = t_r8_c62_12 >> 4;

  assign t_r8_c63_0 = p_7_63 << 1;
  assign t_r8_c63_1 = p_8_62 << 1;
  assign t_r8_c63_2 = p_8_63 << 2;
  assign t_r8_c63_3 = p_8_64 << 1;
  assign t_r8_c63_4 = p_9_63 << 1;
  assign t_r8_c63_5 = t_r8_c63_0 + p_7_62;
  assign t_r8_c63_6 = t_r8_c63_1 + p_7_64;
  assign t_r8_c63_7 = t_r8_c63_2 + t_r8_c63_3;
  assign t_r8_c63_8 = t_r8_c63_4 + p_9_62;
  assign t_r8_c63_9 = t_r8_c63_5 + t_r8_c63_6;
  assign t_r8_c63_10 = t_r8_c63_7 + t_r8_c63_8;
  assign t_r8_c63_11 = t_r8_c63_9 + t_r8_c63_10;
  assign t_r8_c63_12 = t_r8_c63_11 + p_9_64;
  assign out_8_63 = t_r8_c63_12 >> 4;

  assign t_r8_c64_0 = p_7_64 << 1;
  assign t_r8_c64_1 = p_8_63 << 1;
  assign t_r8_c64_2 = p_8_64 << 2;
  assign t_r8_c64_3 = p_8_65 << 1;
  assign t_r8_c64_4 = p_9_64 << 1;
  assign t_r8_c64_5 = t_r8_c64_0 + p_7_63;
  assign t_r8_c64_6 = t_r8_c64_1 + p_7_65;
  assign t_r8_c64_7 = t_r8_c64_2 + t_r8_c64_3;
  assign t_r8_c64_8 = t_r8_c64_4 + p_9_63;
  assign t_r8_c64_9 = t_r8_c64_5 + t_r8_c64_6;
  assign t_r8_c64_10 = t_r8_c64_7 + t_r8_c64_8;
  assign t_r8_c64_11 = t_r8_c64_9 + t_r8_c64_10;
  assign t_r8_c64_12 = t_r8_c64_11 + p_9_65;
  assign out_8_64 = t_r8_c64_12 >> 4;

  assign t_r9_c1_0 = p_8_1 << 1;
  assign t_r9_c1_1 = p_9_0 << 1;
  assign t_r9_c1_2 = p_9_1 << 2;
  assign t_r9_c1_3 = p_9_2 << 1;
  assign t_r9_c1_4 = p_10_1 << 1;
  assign t_r9_c1_5 = t_r9_c1_0 + p_8_0;
  assign t_r9_c1_6 = t_r9_c1_1 + p_8_2;
  assign t_r9_c1_7 = t_r9_c1_2 + t_r9_c1_3;
  assign t_r9_c1_8 = t_r9_c1_4 + p_10_0;
  assign t_r9_c1_9 = t_r9_c1_5 + t_r9_c1_6;
  assign t_r9_c1_10 = t_r9_c1_7 + t_r9_c1_8;
  assign t_r9_c1_11 = t_r9_c1_9 + t_r9_c1_10;
  assign t_r9_c1_12 = t_r9_c1_11 + p_10_2;
  assign out_9_1 = t_r9_c1_12 >> 4;

  assign t_r9_c2_0 = p_8_2 << 1;
  assign t_r9_c2_1 = p_9_1 << 1;
  assign t_r9_c2_2 = p_9_2 << 2;
  assign t_r9_c2_3 = p_9_3 << 1;
  assign t_r9_c2_4 = p_10_2 << 1;
  assign t_r9_c2_5 = t_r9_c2_0 + p_8_1;
  assign t_r9_c2_6 = t_r9_c2_1 + p_8_3;
  assign t_r9_c2_7 = t_r9_c2_2 + t_r9_c2_3;
  assign t_r9_c2_8 = t_r9_c2_4 + p_10_1;
  assign t_r9_c2_9 = t_r9_c2_5 + t_r9_c2_6;
  assign t_r9_c2_10 = t_r9_c2_7 + t_r9_c2_8;
  assign t_r9_c2_11 = t_r9_c2_9 + t_r9_c2_10;
  assign t_r9_c2_12 = t_r9_c2_11 + p_10_3;
  assign out_9_2 = t_r9_c2_12 >> 4;

  assign t_r9_c3_0 = p_8_3 << 1;
  assign t_r9_c3_1 = p_9_2 << 1;
  assign t_r9_c3_2 = p_9_3 << 2;
  assign t_r9_c3_3 = p_9_4 << 1;
  assign t_r9_c3_4 = p_10_3 << 1;
  assign t_r9_c3_5 = t_r9_c3_0 + p_8_2;
  assign t_r9_c3_6 = t_r9_c3_1 + p_8_4;
  assign t_r9_c3_7 = t_r9_c3_2 + t_r9_c3_3;
  assign t_r9_c3_8 = t_r9_c3_4 + p_10_2;
  assign t_r9_c3_9 = t_r9_c3_5 + t_r9_c3_6;
  assign t_r9_c3_10 = t_r9_c3_7 + t_r9_c3_8;
  assign t_r9_c3_11 = t_r9_c3_9 + t_r9_c3_10;
  assign t_r9_c3_12 = t_r9_c3_11 + p_10_4;
  assign out_9_3 = t_r9_c3_12 >> 4;

  assign t_r9_c4_0 = p_8_4 << 1;
  assign t_r9_c4_1 = p_9_3 << 1;
  assign t_r9_c4_2 = p_9_4 << 2;
  assign t_r9_c4_3 = p_9_5 << 1;
  assign t_r9_c4_4 = p_10_4 << 1;
  assign t_r9_c4_5 = t_r9_c4_0 + p_8_3;
  assign t_r9_c4_6 = t_r9_c4_1 + p_8_5;
  assign t_r9_c4_7 = t_r9_c4_2 + t_r9_c4_3;
  assign t_r9_c4_8 = t_r9_c4_4 + p_10_3;
  assign t_r9_c4_9 = t_r9_c4_5 + t_r9_c4_6;
  assign t_r9_c4_10 = t_r9_c4_7 + t_r9_c4_8;
  assign t_r9_c4_11 = t_r9_c4_9 + t_r9_c4_10;
  assign t_r9_c4_12 = t_r9_c4_11 + p_10_5;
  assign out_9_4 = t_r9_c4_12 >> 4;

  assign t_r9_c5_0 = p_8_5 << 1;
  assign t_r9_c5_1 = p_9_4 << 1;
  assign t_r9_c5_2 = p_9_5 << 2;
  assign t_r9_c5_3 = p_9_6 << 1;
  assign t_r9_c5_4 = p_10_5 << 1;
  assign t_r9_c5_5 = t_r9_c5_0 + p_8_4;
  assign t_r9_c5_6 = t_r9_c5_1 + p_8_6;
  assign t_r9_c5_7 = t_r9_c5_2 + t_r9_c5_3;
  assign t_r9_c5_8 = t_r9_c5_4 + p_10_4;
  assign t_r9_c5_9 = t_r9_c5_5 + t_r9_c5_6;
  assign t_r9_c5_10 = t_r9_c5_7 + t_r9_c5_8;
  assign t_r9_c5_11 = t_r9_c5_9 + t_r9_c5_10;
  assign t_r9_c5_12 = t_r9_c5_11 + p_10_6;
  assign out_9_5 = t_r9_c5_12 >> 4;

  assign t_r9_c6_0 = p_8_6 << 1;
  assign t_r9_c6_1 = p_9_5 << 1;
  assign t_r9_c6_2 = p_9_6 << 2;
  assign t_r9_c6_3 = p_9_7 << 1;
  assign t_r9_c6_4 = p_10_6 << 1;
  assign t_r9_c6_5 = t_r9_c6_0 + p_8_5;
  assign t_r9_c6_6 = t_r9_c6_1 + p_8_7;
  assign t_r9_c6_7 = t_r9_c6_2 + t_r9_c6_3;
  assign t_r9_c6_8 = t_r9_c6_4 + p_10_5;
  assign t_r9_c6_9 = t_r9_c6_5 + t_r9_c6_6;
  assign t_r9_c6_10 = t_r9_c6_7 + t_r9_c6_8;
  assign t_r9_c6_11 = t_r9_c6_9 + t_r9_c6_10;
  assign t_r9_c6_12 = t_r9_c6_11 + p_10_7;
  assign out_9_6 = t_r9_c6_12 >> 4;

  assign t_r9_c7_0 = p_8_7 << 1;
  assign t_r9_c7_1 = p_9_6 << 1;
  assign t_r9_c7_2 = p_9_7 << 2;
  assign t_r9_c7_3 = p_9_8 << 1;
  assign t_r9_c7_4 = p_10_7 << 1;
  assign t_r9_c7_5 = t_r9_c7_0 + p_8_6;
  assign t_r9_c7_6 = t_r9_c7_1 + p_8_8;
  assign t_r9_c7_7 = t_r9_c7_2 + t_r9_c7_3;
  assign t_r9_c7_8 = t_r9_c7_4 + p_10_6;
  assign t_r9_c7_9 = t_r9_c7_5 + t_r9_c7_6;
  assign t_r9_c7_10 = t_r9_c7_7 + t_r9_c7_8;
  assign t_r9_c7_11 = t_r9_c7_9 + t_r9_c7_10;
  assign t_r9_c7_12 = t_r9_c7_11 + p_10_8;
  assign out_9_7 = t_r9_c7_12 >> 4;

  assign t_r9_c8_0 = p_8_8 << 1;
  assign t_r9_c8_1 = p_9_7 << 1;
  assign t_r9_c8_2 = p_9_8 << 2;
  assign t_r9_c8_3 = p_9_9 << 1;
  assign t_r9_c8_4 = p_10_8 << 1;
  assign t_r9_c8_5 = t_r9_c8_0 + p_8_7;
  assign t_r9_c8_6 = t_r9_c8_1 + p_8_9;
  assign t_r9_c8_7 = t_r9_c8_2 + t_r9_c8_3;
  assign t_r9_c8_8 = t_r9_c8_4 + p_10_7;
  assign t_r9_c8_9 = t_r9_c8_5 + t_r9_c8_6;
  assign t_r9_c8_10 = t_r9_c8_7 + t_r9_c8_8;
  assign t_r9_c8_11 = t_r9_c8_9 + t_r9_c8_10;
  assign t_r9_c8_12 = t_r9_c8_11 + p_10_9;
  assign out_9_8 = t_r9_c8_12 >> 4;

  assign t_r9_c9_0 = p_8_9 << 1;
  assign t_r9_c9_1 = p_9_8 << 1;
  assign t_r9_c9_2 = p_9_9 << 2;
  assign t_r9_c9_3 = p_9_10 << 1;
  assign t_r9_c9_4 = p_10_9 << 1;
  assign t_r9_c9_5 = t_r9_c9_0 + p_8_8;
  assign t_r9_c9_6 = t_r9_c9_1 + p_8_10;
  assign t_r9_c9_7 = t_r9_c9_2 + t_r9_c9_3;
  assign t_r9_c9_8 = t_r9_c9_4 + p_10_8;
  assign t_r9_c9_9 = t_r9_c9_5 + t_r9_c9_6;
  assign t_r9_c9_10 = t_r9_c9_7 + t_r9_c9_8;
  assign t_r9_c9_11 = t_r9_c9_9 + t_r9_c9_10;
  assign t_r9_c9_12 = t_r9_c9_11 + p_10_10;
  assign out_9_9 = t_r9_c9_12 >> 4;

  assign t_r9_c10_0 = p_8_10 << 1;
  assign t_r9_c10_1 = p_9_9 << 1;
  assign t_r9_c10_2 = p_9_10 << 2;
  assign t_r9_c10_3 = p_9_11 << 1;
  assign t_r9_c10_4 = p_10_10 << 1;
  assign t_r9_c10_5 = t_r9_c10_0 + p_8_9;
  assign t_r9_c10_6 = t_r9_c10_1 + p_8_11;
  assign t_r9_c10_7 = t_r9_c10_2 + t_r9_c10_3;
  assign t_r9_c10_8 = t_r9_c10_4 + p_10_9;
  assign t_r9_c10_9 = t_r9_c10_5 + t_r9_c10_6;
  assign t_r9_c10_10 = t_r9_c10_7 + t_r9_c10_8;
  assign t_r9_c10_11 = t_r9_c10_9 + t_r9_c10_10;
  assign t_r9_c10_12 = t_r9_c10_11 + p_10_11;
  assign out_9_10 = t_r9_c10_12 >> 4;

  assign t_r9_c11_0 = p_8_11 << 1;
  assign t_r9_c11_1 = p_9_10 << 1;
  assign t_r9_c11_2 = p_9_11 << 2;
  assign t_r9_c11_3 = p_9_12 << 1;
  assign t_r9_c11_4 = p_10_11 << 1;
  assign t_r9_c11_5 = t_r9_c11_0 + p_8_10;
  assign t_r9_c11_6 = t_r9_c11_1 + p_8_12;
  assign t_r9_c11_7 = t_r9_c11_2 + t_r9_c11_3;
  assign t_r9_c11_8 = t_r9_c11_4 + p_10_10;
  assign t_r9_c11_9 = t_r9_c11_5 + t_r9_c11_6;
  assign t_r9_c11_10 = t_r9_c11_7 + t_r9_c11_8;
  assign t_r9_c11_11 = t_r9_c11_9 + t_r9_c11_10;
  assign t_r9_c11_12 = t_r9_c11_11 + p_10_12;
  assign out_9_11 = t_r9_c11_12 >> 4;

  assign t_r9_c12_0 = p_8_12 << 1;
  assign t_r9_c12_1 = p_9_11 << 1;
  assign t_r9_c12_2 = p_9_12 << 2;
  assign t_r9_c12_3 = p_9_13 << 1;
  assign t_r9_c12_4 = p_10_12 << 1;
  assign t_r9_c12_5 = t_r9_c12_0 + p_8_11;
  assign t_r9_c12_6 = t_r9_c12_1 + p_8_13;
  assign t_r9_c12_7 = t_r9_c12_2 + t_r9_c12_3;
  assign t_r9_c12_8 = t_r9_c12_4 + p_10_11;
  assign t_r9_c12_9 = t_r9_c12_5 + t_r9_c12_6;
  assign t_r9_c12_10 = t_r9_c12_7 + t_r9_c12_8;
  assign t_r9_c12_11 = t_r9_c12_9 + t_r9_c12_10;
  assign t_r9_c12_12 = t_r9_c12_11 + p_10_13;
  assign out_9_12 = t_r9_c12_12 >> 4;

  assign t_r9_c13_0 = p_8_13 << 1;
  assign t_r9_c13_1 = p_9_12 << 1;
  assign t_r9_c13_2 = p_9_13 << 2;
  assign t_r9_c13_3 = p_9_14 << 1;
  assign t_r9_c13_4 = p_10_13 << 1;
  assign t_r9_c13_5 = t_r9_c13_0 + p_8_12;
  assign t_r9_c13_6 = t_r9_c13_1 + p_8_14;
  assign t_r9_c13_7 = t_r9_c13_2 + t_r9_c13_3;
  assign t_r9_c13_8 = t_r9_c13_4 + p_10_12;
  assign t_r9_c13_9 = t_r9_c13_5 + t_r9_c13_6;
  assign t_r9_c13_10 = t_r9_c13_7 + t_r9_c13_8;
  assign t_r9_c13_11 = t_r9_c13_9 + t_r9_c13_10;
  assign t_r9_c13_12 = t_r9_c13_11 + p_10_14;
  assign out_9_13 = t_r9_c13_12 >> 4;

  assign t_r9_c14_0 = p_8_14 << 1;
  assign t_r9_c14_1 = p_9_13 << 1;
  assign t_r9_c14_2 = p_9_14 << 2;
  assign t_r9_c14_3 = p_9_15 << 1;
  assign t_r9_c14_4 = p_10_14 << 1;
  assign t_r9_c14_5 = t_r9_c14_0 + p_8_13;
  assign t_r9_c14_6 = t_r9_c14_1 + p_8_15;
  assign t_r9_c14_7 = t_r9_c14_2 + t_r9_c14_3;
  assign t_r9_c14_8 = t_r9_c14_4 + p_10_13;
  assign t_r9_c14_9 = t_r9_c14_5 + t_r9_c14_6;
  assign t_r9_c14_10 = t_r9_c14_7 + t_r9_c14_8;
  assign t_r9_c14_11 = t_r9_c14_9 + t_r9_c14_10;
  assign t_r9_c14_12 = t_r9_c14_11 + p_10_15;
  assign out_9_14 = t_r9_c14_12 >> 4;

  assign t_r9_c15_0 = p_8_15 << 1;
  assign t_r9_c15_1 = p_9_14 << 1;
  assign t_r9_c15_2 = p_9_15 << 2;
  assign t_r9_c15_3 = p_9_16 << 1;
  assign t_r9_c15_4 = p_10_15 << 1;
  assign t_r9_c15_5 = t_r9_c15_0 + p_8_14;
  assign t_r9_c15_6 = t_r9_c15_1 + p_8_16;
  assign t_r9_c15_7 = t_r9_c15_2 + t_r9_c15_3;
  assign t_r9_c15_8 = t_r9_c15_4 + p_10_14;
  assign t_r9_c15_9 = t_r9_c15_5 + t_r9_c15_6;
  assign t_r9_c15_10 = t_r9_c15_7 + t_r9_c15_8;
  assign t_r9_c15_11 = t_r9_c15_9 + t_r9_c15_10;
  assign t_r9_c15_12 = t_r9_c15_11 + p_10_16;
  assign out_9_15 = t_r9_c15_12 >> 4;

  assign t_r9_c16_0 = p_8_16 << 1;
  assign t_r9_c16_1 = p_9_15 << 1;
  assign t_r9_c16_2 = p_9_16 << 2;
  assign t_r9_c16_3 = p_9_17 << 1;
  assign t_r9_c16_4 = p_10_16 << 1;
  assign t_r9_c16_5 = t_r9_c16_0 + p_8_15;
  assign t_r9_c16_6 = t_r9_c16_1 + p_8_17;
  assign t_r9_c16_7 = t_r9_c16_2 + t_r9_c16_3;
  assign t_r9_c16_8 = t_r9_c16_4 + p_10_15;
  assign t_r9_c16_9 = t_r9_c16_5 + t_r9_c16_6;
  assign t_r9_c16_10 = t_r9_c16_7 + t_r9_c16_8;
  assign t_r9_c16_11 = t_r9_c16_9 + t_r9_c16_10;
  assign t_r9_c16_12 = t_r9_c16_11 + p_10_17;
  assign out_9_16 = t_r9_c16_12 >> 4;

  assign t_r9_c17_0 = p_8_17 << 1;
  assign t_r9_c17_1 = p_9_16 << 1;
  assign t_r9_c17_2 = p_9_17 << 2;
  assign t_r9_c17_3 = p_9_18 << 1;
  assign t_r9_c17_4 = p_10_17 << 1;
  assign t_r9_c17_5 = t_r9_c17_0 + p_8_16;
  assign t_r9_c17_6 = t_r9_c17_1 + p_8_18;
  assign t_r9_c17_7 = t_r9_c17_2 + t_r9_c17_3;
  assign t_r9_c17_8 = t_r9_c17_4 + p_10_16;
  assign t_r9_c17_9 = t_r9_c17_5 + t_r9_c17_6;
  assign t_r9_c17_10 = t_r9_c17_7 + t_r9_c17_8;
  assign t_r9_c17_11 = t_r9_c17_9 + t_r9_c17_10;
  assign t_r9_c17_12 = t_r9_c17_11 + p_10_18;
  assign out_9_17 = t_r9_c17_12 >> 4;

  assign t_r9_c18_0 = p_8_18 << 1;
  assign t_r9_c18_1 = p_9_17 << 1;
  assign t_r9_c18_2 = p_9_18 << 2;
  assign t_r9_c18_3 = p_9_19 << 1;
  assign t_r9_c18_4 = p_10_18 << 1;
  assign t_r9_c18_5 = t_r9_c18_0 + p_8_17;
  assign t_r9_c18_6 = t_r9_c18_1 + p_8_19;
  assign t_r9_c18_7 = t_r9_c18_2 + t_r9_c18_3;
  assign t_r9_c18_8 = t_r9_c18_4 + p_10_17;
  assign t_r9_c18_9 = t_r9_c18_5 + t_r9_c18_6;
  assign t_r9_c18_10 = t_r9_c18_7 + t_r9_c18_8;
  assign t_r9_c18_11 = t_r9_c18_9 + t_r9_c18_10;
  assign t_r9_c18_12 = t_r9_c18_11 + p_10_19;
  assign out_9_18 = t_r9_c18_12 >> 4;

  assign t_r9_c19_0 = p_8_19 << 1;
  assign t_r9_c19_1 = p_9_18 << 1;
  assign t_r9_c19_2 = p_9_19 << 2;
  assign t_r9_c19_3 = p_9_20 << 1;
  assign t_r9_c19_4 = p_10_19 << 1;
  assign t_r9_c19_5 = t_r9_c19_0 + p_8_18;
  assign t_r9_c19_6 = t_r9_c19_1 + p_8_20;
  assign t_r9_c19_7 = t_r9_c19_2 + t_r9_c19_3;
  assign t_r9_c19_8 = t_r9_c19_4 + p_10_18;
  assign t_r9_c19_9 = t_r9_c19_5 + t_r9_c19_6;
  assign t_r9_c19_10 = t_r9_c19_7 + t_r9_c19_8;
  assign t_r9_c19_11 = t_r9_c19_9 + t_r9_c19_10;
  assign t_r9_c19_12 = t_r9_c19_11 + p_10_20;
  assign out_9_19 = t_r9_c19_12 >> 4;

  assign t_r9_c20_0 = p_8_20 << 1;
  assign t_r9_c20_1 = p_9_19 << 1;
  assign t_r9_c20_2 = p_9_20 << 2;
  assign t_r9_c20_3 = p_9_21 << 1;
  assign t_r9_c20_4 = p_10_20 << 1;
  assign t_r9_c20_5 = t_r9_c20_0 + p_8_19;
  assign t_r9_c20_6 = t_r9_c20_1 + p_8_21;
  assign t_r9_c20_7 = t_r9_c20_2 + t_r9_c20_3;
  assign t_r9_c20_8 = t_r9_c20_4 + p_10_19;
  assign t_r9_c20_9 = t_r9_c20_5 + t_r9_c20_6;
  assign t_r9_c20_10 = t_r9_c20_7 + t_r9_c20_8;
  assign t_r9_c20_11 = t_r9_c20_9 + t_r9_c20_10;
  assign t_r9_c20_12 = t_r9_c20_11 + p_10_21;
  assign out_9_20 = t_r9_c20_12 >> 4;

  assign t_r9_c21_0 = p_8_21 << 1;
  assign t_r9_c21_1 = p_9_20 << 1;
  assign t_r9_c21_2 = p_9_21 << 2;
  assign t_r9_c21_3 = p_9_22 << 1;
  assign t_r9_c21_4 = p_10_21 << 1;
  assign t_r9_c21_5 = t_r9_c21_0 + p_8_20;
  assign t_r9_c21_6 = t_r9_c21_1 + p_8_22;
  assign t_r9_c21_7 = t_r9_c21_2 + t_r9_c21_3;
  assign t_r9_c21_8 = t_r9_c21_4 + p_10_20;
  assign t_r9_c21_9 = t_r9_c21_5 + t_r9_c21_6;
  assign t_r9_c21_10 = t_r9_c21_7 + t_r9_c21_8;
  assign t_r9_c21_11 = t_r9_c21_9 + t_r9_c21_10;
  assign t_r9_c21_12 = t_r9_c21_11 + p_10_22;
  assign out_9_21 = t_r9_c21_12 >> 4;

  assign t_r9_c22_0 = p_8_22 << 1;
  assign t_r9_c22_1 = p_9_21 << 1;
  assign t_r9_c22_2 = p_9_22 << 2;
  assign t_r9_c22_3 = p_9_23 << 1;
  assign t_r9_c22_4 = p_10_22 << 1;
  assign t_r9_c22_5 = t_r9_c22_0 + p_8_21;
  assign t_r9_c22_6 = t_r9_c22_1 + p_8_23;
  assign t_r9_c22_7 = t_r9_c22_2 + t_r9_c22_3;
  assign t_r9_c22_8 = t_r9_c22_4 + p_10_21;
  assign t_r9_c22_9 = t_r9_c22_5 + t_r9_c22_6;
  assign t_r9_c22_10 = t_r9_c22_7 + t_r9_c22_8;
  assign t_r9_c22_11 = t_r9_c22_9 + t_r9_c22_10;
  assign t_r9_c22_12 = t_r9_c22_11 + p_10_23;
  assign out_9_22 = t_r9_c22_12 >> 4;

  assign t_r9_c23_0 = p_8_23 << 1;
  assign t_r9_c23_1 = p_9_22 << 1;
  assign t_r9_c23_2 = p_9_23 << 2;
  assign t_r9_c23_3 = p_9_24 << 1;
  assign t_r9_c23_4 = p_10_23 << 1;
  assign t_r9_c23_5 = t_r9_c23_0 + p_8_22;
  assign t_r9_c23_6 = t_r9_c23_1 + p_8_24;
  assign t_r9_c23_7 = t_r9_c23_2 + t_r9_c23_3;
  assign t_r9_c23_8 = t_r9_c23_4 + p_10_22;
  assign t_r9_c23_9 = t_r9_c23_5 + t_r9_c23_6;
  assign t_r9_c23_10 = t_r9_c23_7 + t_r9_c23_8;
  assign t_r9_c23_11 = t_r9_c23_9 + t_r9_c23_10;
  assign t_r9_c23_12 = t_r9_c23_11 + p_10_24;
  assign out_9_23 = t_r9_c23_12 >> 4;

  assign t_r9_c24_0 = p_8_24 << 1;
  assign t_r9_c24_1 = p_9_23 << 1;
  assign t_r9_c24_2 = p_9_24 << 2;
  assign t_r9_c24_3 = p_9_25 << 1;
  assign t_r9_c24_4 = p_10_24 << 1;
  assign t_r9_c24_5 = t_r9_c24_0 + p_8_23;
  assign t_r9_c24_6 = t_r9_c24_1 + p_8_25;
  assign t_r9_c24_7 = t_r9_c24_2 + t_r9_c24_3;
  assign t_r9_c24_8 = t_r9_c24_4 + p_10_23;
  assign t_r9_c24_9 = t_r9_c24_5 + t_r9_c24_6;
  assign t_r9_c24_10 = t_r9_c24_7 + t_r9_c24_8;
  assign t_r9_c24_11 = t_r9_c24_9 + t_r9_c24_10;
  assign t_r9_c24_12 = t_r9_c24_11 + p_10_25;
  assign out_9_24 = t_r9_c24_12 >> 4;

  assign t_r9_c25_0 = p_8_25 << 1;
  assign t_r9_c25_1 = p_9_24 << 1;
  assign t_r9_c25_2 = p_9_25 << 2;
  assign t_r9_c25_3 = p_9_26 << 1;
  assign t_r9_c25_4 = p_10_25 << 1;
  assign t_r9_c25_5 = t_r9_c25_0 + p_8_24;
  assign t_r9_c25_6 = t_r9_c25_1 + p_8_26;
  assign t_r9_c25_7 = t_r9_c25_2 + t_r9_c25_3;
  assign t_r9_c25_8 = t_r9_c25_4 + p_10_24;
  assign t_r9_c25_9 = t_r9_c25_5 + t_r9_c25_6;
  assign t_r9_c25_10 = t_r9_c25_7 + t_r9_c25_8;
  assign t_r9_c25_11 = t_r9_c25_9 + t_r9_c25_10;
  assign t_r9_c25_12 = t_r9_c25_11 + p_10_26;
  assign out_9_25 = t_r9_c25_12 >> 4;

  assign t_r9_c26_0 = p_8_26 << 1;
  assign t_r9_c26_1 = p_9_25 << 1;
  assign t_r9_c26_2 = p_9_26 << 2;
  assign t_r9_c26_3 = p_9_27 << 1;
  assign t_r9_c26_4 = p_10_26 << 1;
  assign t_r9_c26_5 = t_r9_c26_0 + p_8_25;
  assign t_r9_c26_6 = t_r9_c26_1 + p_8_27;
  assign t_r9_c26_7 = t_r9_c26_2 + t_r9_c26_3;
  assign t_r9_c26_8 = t_r9_c26_4 + p_10_25;
  assign t_r9_c26_9 = t_r9_c26_5 + t_r9_c26_6;
  assign t_r9_c26_10 = t_r9_c26_7 + t_r9_c26_8;
  assign t_r9_c26_11 = t_r9_c26_9 + t_r9_c26_10;
  assign t_r9_c26_12 = t_r9_c26_11 + p_10_27;
  assign out_9_26 = t_r9_c26_12 >> 4;

  assign t_r9_c27_0 = p_8_27 << 1;
  assign t_r9_c27_1 = p_9_26 << 1;
  assign t_r9_c27_2 = p_9_27 << 2;
  assign t_r9_c27_3 = p_9_28 << 1;
  assign t_r9_c27_4 = p_10_27 << 1;
  assign t_r9_c27_5 = t_r9_c27_0 + p_8_26;
  assign t_r9_c27_6 = t_r9_c27_1 + p_8_28;
  assign t_r9_c27_7 = t_r9_c27_2 + t_r9_c27_3;
  assign t_r9_c27_8 = t_r9_c27_4 + p_10_26;
  assign t_r9_c27_9 = t_r9_c27_5 + t_r9_c27_6;
  assign t_r9_c27_10 = t_r9_c27_7 + t_r9_c27_8;
  assign t_r9_c27_11 = t_r9_c27_9 + t_r9_c27_10;
  assign t_r9_c27_12 = t_r9_c27_11 + p_10_28;
  assign out_9_27 = t_r9_c27_12 >> 4;

  assign t_r9_c28_0 = p_8_28 << 1;
  assign t_r9_c28_1 = p_9_27 << 1;
  assign t_r9_c28_2 = p_9_28 << 2;
  assign t_r9_c28_3 = p_9_29 << 1;
  assign t_r9_c28_4 = p_10_28 << 1;
  assign t_r9_c28_5 = t_r9_c28_0 + p_8_27;
  assign t_r9_c28_6 = t_r9_c28_1 + p_8_29;
  assign t_r9_c28_7 = t_r9_c28_2 + t_r9_c28_3;
  assign t_r9_c28_8 = t_r9_c28_4 + p_10_27;
  assign t_r9_c28_9 = t_r9_c28_5 + t_r9_c28_6;
  assign t_r9_c28_10 = t_r9_c28_7 + t_r9_c28_8;
  assign t_r9_c28_11 = t_r9_c28_9 + t_r9_c28_10;
  assign t_r9_c28_12 = t_r9_c28_11 + p_10_29;
  assign out_9_28 = t_r9_c28_12 >> 4;

  assign t_r9_c29_0 = p_8_29 << 1;
  assign t_r9_c29_1 = p_9_28 << 1;
  assign t_r9_c29_2 = p_9_29 << 2;
  assign t_r9_c29_3 = p_9_30 << 1;
  assign t_r9_c29_4 = p_10_29 << 1;
  assign t_r9_c29_5 = t_r9_c29_0 + p_8_28;
  assign t_r9_c29_6 = t_r9_c29_1 + p_8_30;
  assign t_r9_c29_7 = t_r9_c29_2 + t_r9_c29_3;
  assign t_r9_c29_8 = t_r9_c29_4 + p_10_28;
  assign t_r9_c29_9 = t_r9_c29_5 + t_r9_c29_6;
  assign t_r9_c29_10 = t_r9_c29_7 + t_r9_c29_8;
  assign t_r9_c29_11 = t_r9_c29_9 + t_r9_c29_10;
  assign t_r9_c29_12 = t_r9_c29_11 + p_10_30;
  assign out_9_29 = t_r9_c29_12 >> 4;

  assign t_r9_c30_0 = p_8_30 << 1;
  assign t_r9_c30_1 = p_9_29 << 1;
  assign t_r9_c30_2 = p_9_30 << 2;
  assign t_r9_c30_3 = p_9_31 << 1;
  assign t_r9_c30_4 = p_10_30 << 1;
  assign t_r9_c30_5 = t_r9_c30_0 + p_8_29;
  assign t_r9_c30_6 = t_r9_c30_1 + p_8_31;
  assign t_r9_c30_7 = t_r9_c30_2 + t_r9_c30_3;
  assign t_r9_c30_8 = t_r9_c30_4 + p_10_29;
  assign t_r9_c30_9 = t_r9_c30_5 + t_r9_c30_6;
  assign t_r9_c30_10 = t_r9_c30_7 + t_r9_c30_8;
  assign t_r9_c30_11 = t_r9_c30_9 + t_r9_c30_10;
  assign t_r9_c30_12 = t_r9_c30_11 + p_10_31;
  assign out_9_30 = t_r9_c30_12 >> 4;

  assign t_r9_c31_0 = p_8_31 << 1;
  assign t_r9_c31_1 = p_9_30 << 1;
  assign t_r9_c31_2 = p_9_31 << 2;
  assign t_r9_c31_3 = p_9_32 << 1;
  assign t_r9_c31_4 = p_10_31 << 1;
  assign t_r9_c31_5 = t_r9_c31_0 + p_8_30;
  assign t_r9_c31_6 = t_r9_c31_1 + p_8_32;
  assign t_r9_c31_7 = t_r9_c31_2 + t_r9_c31_3;
  assign t_r9_c31_8 = t_r9_c31_4 + p_10_30;
  assign t_r9_c31_9 = t_r9_c31_5 + t_r9_c31_6;
  assign t_r9_c31_10 = t_r9_c31_7 + t_r9_c31_8;
  assign t_r9_c31_11 = t_r9_c31_9 + t_r9_c31_10;
  assign t_r9_c31_12 = t_r9_c31_11 + p_10_32;
  assign out_9_31 = t_r9_c31_12 >> 4;

  assign t_r9_c32_0 = p_8_32 << 1;
  assign t_r9_c32_1 = p_9_31 << 1;
  assign t_r9_c32_2 = p_9_32 << 2;
  assign t_r9_c32_3 = p_9_33 << 1;
  assign t_r9_c32_4 = p_10_32 << 1;
  assign t_r9_c32_5 = t_r9_c32_0 + p_8_31;
  assign t_r9_c32_6 = t_r9_c32_1 + p_8_33;
  assign t_r9_c32_7 = t_r9_c32_2 + t_r9_c32_3;
  assign t_r9_c32_8 = t_r9_c32_4 + p_10_31;
  assign t_r9_c32_9 = t_r9_c32_5 + t_r9_c32_6;
  assign t_r9_c32_10 = t_r9_c32_7 + t_r9_c32_8;
  assign t_r9_c32_11 = t_r9_c32_9 + t_r9_c32_10;
  assign t_r9_c32_12 = t_r9_c32_11 + p_10_33;
  assign out_9_32 = t_r9_c32_12 >> 4;

  assign t_r9_c33_0 = p_8_33 << 1;
  assign t_r9_c33_1 = p_9_32 << 1;
  assign t_r9_c33_2 = p_9_33 << 2;
  assign t_r9_c33_3 = p_9_34 << 1;
  assign t_r9_c33_4 = p_10_33 << 1;
  assign t_r9_c33_5 = t_r9_c33_0 + p_8_32;
  assign t_r9_c33_6 = t_r9_c33_1 + p_8_34;
  assign t_r9_c33_7 = t_r9_c33_2 + t_r9_c33_3;
  assign t_r9_c33_8 = t_r9_c33_4 + p_10_32;
  assign t_r9_c33_9 = t_r9_c33_5 + t_r9_c33_6;
  assign t_r9_c33_10 = t_r9_c33_7 + t_r9_c33_8;
  assign t_r9_c33_11 = t_r9_c33_9 + t_r9_c33_10;
  assign t_r9_c33_12 = t_r9_c33_11 + p_10_34;
  assign out_9_33 = t_r9_c33_12 >> 4;

  assign t_r9_c34_0 = p_8_34 << 1;
  assign t_r9_c34_1 = p_9_33 << 1;
  assign t_r9_c34_2 = p_9_34 << 2;
  assign t_r9_c34_3 = p_9_35 << 1;
  assign t_r9_c34_4 = p_10_34 << 1;
  assign t_r9_c34_5 = t_r9_c34_0 + p_8_33;
  assign t_r9_c34_6 = t_r9_c34_1 + p_8_35;
  assign t_r9_c34_7 = t_r9_c34_2 + t_r9_c34_3;
  assign t_r9_c34_8 = t_r9_c34_4 + p_10_33;
  assign t_r9_c34_9 = t_r9_c34_5 + t_r9_c34_6;
  assign t_r9_c34_10 = t_r9_c34_7 + t_r9_c34_8;
  assign t_r9_c34_11 = t_r9_c34_9 + t_r9_c34_10;
  assign t_r9_c34_12 = t_r9_c34_11 + p_10_35;
  assign out_9_34 = t_r9_c34_12 >> 4;

  assign t_r9_c35_0 = p_8_35 << 1;
  assign t_r9_c35_1 = p_9_34 << 1;
  assign t_r9_c35_2 = p_9_35 << 2;
  assign t_r9_c35_3 = p_9_36 << 1;
  assign t_r9_c35_4 = p_10_35 << 1;
  assign t_r9_c35_5 = t_r9_c35_0 + p_8_34;
  assign t_r9_c35_6 = t_r9_c35_1 + p_8_36;
  assign t_r9_c35_7 = t_r9_c35_2 + t_r9_c35_3;
  assign t_r9_c35_8 = t_r9_c35_4 + p_10_34;
  assign t_r9_c35_9 = t_r9_c35_5 + t_r9_c35_6;
  assign t_r9_c35_10 = t_r9_c35_7 + t_r9_c35_8;
  assign t_r9_c35_11 = t_r9_c35_9 + t_r9_c35_10;
  assign t_r9_c35_12 = t_r9_c35_11 + p_10_36;
  assign out_9_35 = t_r9_c35_12 >> 4;

  assign t_r9_c36_0 = p_8_36 << 1;
  assign t_r9_c36_1 = p_9_35 << 1;
  assign t_r9_c36_2 = p_9_36 << 2;
  assign t_r9_c36_3 = p_9_37 << 1;
  assign t_r9_c36_4 = p_10_36 << 1;
  assign t_r9_c36_5 = t_r9_c36_0 + p_8_35;
  assign t_r9_c36_6 = t_r9_c36_1 + p_8_37;
  assign t_r9_c36_7 = t_r9_c36_2 + t_r9_c36_3;
  assign t_r9_c36_8 = t_r9_c36_4 + p_10_35;
  assign t_r9_c36_9 = t_r9_c36_5 + t_r9_c36_6;
  assign t_r9_c36_10 = t_r9_c36_7 + t_r9_c36_8;
  assign t_r9_c36_11 = t_r9_c36_9 + t_r9_c36_10;
  assign t_r9_c36_12 = t_r9_c36_11 + p_10_37;
  assign out_9_36 = t_r9_c36_12 >> 4;

  assign t_r9_c37_0 = p_8_37 << 1;
  assign t_r9_c37_1 = p_9_36 << 1;
  assign t_r9_c37_2 = p_9_37 << 2;
  assign t_r9_c37_3 = p_9_38 << 1;
  assign t_r9_c37_4 = p_10_37 << 1;
  assign t_r9_c37_5 = t_r9_c37_0 + p_8_36;
  assign t_r9_c37_6 = t_r9_c37_1 + p_8_38;
  assign t_r9_c37_7 = t_r9_c37_2 + t_r9_c37_3;
  assign t_r9_c37_8 = t_r9_c37_4 + p_10_36;
  assign t_r9_c37_9 = t_r9_c37_5 + t_r9_c37_6;
  assign t_r9_c37_10 = t_r9_c37_7 + t_r9_c37_8;
  assign t_r9_c37_11 = t_r9_c37_9 + t_r9_c37_10;
  assign t_r9_c37_12 = t_r9_c37_11 + p_10_38;
  assign out_9_37 = t_r9_c37_12 >> 4;

  assign t_r9_c38_0 = p_8_38 << 1;
  assign t_r9_c38_1 = p_9_37 << 1;
  assign t_r9_c38_2 = p_9_38 << 2;
  assign t_r9_c38_3 = p_9_39 << 1;
  assign t_r9_c38_4 = p_10_38 << 1;
  assign t_r9_c38_5 = t_r9_c38_0 + p_8_37;
  assign t_r9_c38_6 = t_r9_c38_1 + p_8_39;
  assign t_r9_c38_7 = t_r9_c38_2 + t_r9_c38_3;
  assign t_r9_c38_8 = t_r9_c38_4 + p_10_37;
  assign t_r9_c38_9 = t_r9_c38_5 + t_r9_c38_6;
  assign t_r9_c38_10 = t_r9_c38_7 + t_r9_c38_8;
  assign t_r9_c38_11 = t_r9_c38_9 + t_r9_c38_10;
  assign t_r9_c38_12 = t_r9_c38_11 + p_10_39;
  assign out_9_38 = t_r9_c38_12 >> 4;

  assign t_r9_c39_0 = p_8_39 << 1;
  assign t_r9_c39_1 = p_9_38 << 1;
  assign t_r9_c39_2 = p_9_39 << 2;
  assign t_r9_c39_3 = p_9_40 << 1;
  assign t_r9_c39_4 = p_10_39 << 1;
  assign t_r9_c39_5 = t_r9_c39_0 + p_8_38;
  assign t_r9_c39_6 = t_r9_c39_1 + p_8_40;
  assign t_r9_c39_7 = t_r9_c39_2 + t_r9_c39_3;
  assign t_r9_c39_8 = t_r9_c39_4 + p_10_38;
  assign t_r9_c39_9 = t_r9_c39_5 + t_r9_c39_6;
  assign t_r9_c39_10 = t_r9_c39_7 + t_r9_c39_8;
  assign t_r9_c39_11 = t_r9_c39_9 + t_r9_c39_10;
  assign t_r9_c39_12 = t_r9_c39_11 + p_10_40;
  assign out_9_39 = t_r9_c39_12 >> 4;

  assign t_r9_c40_0 = p_8_40 << 1;
  assign t_r9_c40_1 = p_9_39 << 1;
  assign t_r9_c40_2 = p_9_40 << 2;
  assign t_r9_c40_3 = p_9_41 << 1;
  assign t_r9_c40_4 = p_10_40 << 1;
  assign t_r9_c40_5 = t_r9_c40_0 + p_8_39;
  assign t_r9_c40_6 = t_r9_c40_1 + p_8_41;
  assign t_r9_c40_7 = t_r9_c40_2 + t_r9_c40_3;
  assign t_r9_c40_8 = t_r9_c40_4 + p_10_39;
  assign t_r9_c40_9 = t_r9_c40_5 + t_r9_c40_6;
  assign t_r9_c40_10 = t_r9_c40_7 + t_r9_c40_8;
  assign t_r9_c40_11 = t_r9_c40_9 + t_r9_c40_10;
  assign t_r9_c40_12 = t_r9_c40_11 + p_10_41;
  assign out_9_40 = t_r9_c40_12 >> 4;

  assign t_r9_c41_0 = p_8_41 << 1;
  assign t_r9_c41_1 = p_9_40 << 1;
  assign t_r9_c41_2 = p_9_41 << 2;
  assign t_r9_c41_3 = p_9_42 << 1;
  assign t_r9_c41_4 = p_10_41 << 1;
  assign t_r9_c41_5 = t_r9_c41_0 + p_8_40;
  assign t_r9_c41_6 = t_r9_c41_1 + p_8_42;
  assign t_r9_c41_7 = t_r9_c41_2 + t_r9_c41_3;
  assign t_r9_c41_8 = t_r9_c41_4 + p_10_40;
  assign t_r9_c41_9 = t_r9_c41_5 + t_r9_c41_6;
  assign t_r9_c41_10 = t_r9_c41_7 + t_r9_c41_8;
  assign t_r9_c41_11 = t_r9_c41_9 + t_r9_c41_10;
  assign t_r9_c41_12 = t_r9_c41_11 + p_10_42;
  assign out_9_41 = t_r9_c41_12 >> 4;

  assign t_r9_c42_0 = p_8_42 << 1;
  assign t_r9_c42_1 = p_9_41 << 1;
  assign t_r9_c42_2 = p_9_42 << 2;
  assign t_r9_c42_3 = p_9_43 << 1;
  assign t_r9_c42_4 = p_10_42 << 1;
  assign t_r9_c42_5 = t_r9_c42_0 + p_8_41;
  assign t_r9_c42_6 = t_r9_c42_1 + p_8_43;
  assign t_r9_c42_7 = t_r9_c42_2 + t_r9_c42_3;
  assign t_r9_c42_8 = t_r9_c42_4 + p_10_41;
  assign t_r9_c42_9 = t_r9_c42_5 + t_r9_c42_6;
  assign t_r9_c42_10 = t_r9_c42_7 + t_r9_c42_8;
  assign t_r9_c42_11 = t_r9_c42_9 + t_r9_c42_10;
  assign t_r9_c42_12 = t_r9_c42_11 + p_10_43;
  assign out_9_42 = t_r9_c42_12 >> 4;

  assign t_r9_c43_0 = p_8_43 << 1;
  assign t_r9_c43_1 = p_9_42 << 1;
  assign t_r9_c43_2 = p_9_43 << 2;
  assign t_r9_c43_3 = p_9_44 << 1;
  assign t_r9_c43_4 = p_10_43 << 1;
  assign t_r9_c43_5 = t_r9_c43_0 + p_8_42;
  assign t_r9_c43_6 = t_r9_c43_1 + p_8_44;
  assign t_r9_c43_7 = t_r9_c43_2 + t_r9_c43_3;
  assign t_r9_c43_8 = t_r9_c43_4 + p_10_42;
  assign t_r9_c43_9 = t_r9_c43_5 + t_r9_c43_6;
  assign t_r9_c43_10 = t_r9_c43_7 + t_r9_c43_8;
  assign t_r9_c43_11 = t_r9_c43_9 + t_r9_c43_10;
  assign t_r9_c43_12 = t_r9_c43_11 + p_10_44;
  assign out_9_43 = t_r9_c43_12 >> 4;

  assign t_r9_c44_0 = p_8_44 << 1;
  assign t_r9_c44_1 = p_9_43 << 1;
  assign t_r9_c44_2 = p_9_44 << 2;
  assign t_r9_c44_3 = p_9_45 << 1;
  assign t_r9_c44_4 = p_10_44 << 1;
  assign t_r9_c44_5 = t_r9_c44_0 + p_8_43;
  assign t_r9_c44_6 = t_r9_c44_1 + p_8_45;
  assign t_r9_c44_7 = t_r9_c44_2 + t_r9_c44_3;
  assign t_r9_c44_8 = t_r9_c44_4 + p_10_43;
  assign t_r9_c44_9 = t_r9_c44_5 + t_r9_c44_6;
  assign t_r9_c44_10 = t_r9_c44_7 + t_r9_c44_8;
  assign t_r9_c44_11 = t_r9_c44_9 + t_r9_c44_10;
  assign t_r9_c44_12 = t_r9_c44_11 + p_10_45;
  assign out_9_44 = t_r9_c44_12 >> 4;

  assign t_r9_c45_0 = p_8_45 << 1;
  assign t_r9_c45_1 = p_9_44 << 1;
  assign t_r9_c45_2 = p_9_45 << 2;
  assign t_r9_c45_3 = p_9_46 << 1;
  assign t_r9_c45_4 = p_10_45 << 1;
  assign t_r9_c45_5 = t_r9_c45_0 + p_8_44;
  assign t_r9_c45_6 = t_r9_c45_1 + p_8_46;
  assign t_r9_c45_7 = t_r9_c45_2 + t_r9_c45_3;
  assign t_r9_c45_8 = t_r9_c45_4 + p_10_44;
  assign t_r9_c45_9 = t_r9_c45_5 + t_r9_c45_6;
  assign t_r9_c45_10 = t_r9_c45_7 + t_r9_c45_8;
  assign t_r9_c45_11 = t_r9_c45_9 + t_r9_c45_10;
  assign t_r9_c45_12 = t_r9_c45_11 + p_10_46;
  assign out_9_45 = t_r9_c45_12 >> 4;

  assign t_r9_c46_0 = p_8_46 << 1;
  assign t_r9_c46_1 = p_9_45 << 1;
  assign t_r9_c46_2 = p_9_46 << 2;
  assign t_r9_c46_3 = p_9_47 << 1;
  assign t_r9_c46_4 = p_10_46 << 1;
  assign t_r9_c46_5 = t_r9_c46_0 + p_8_45;
  assign t_r9_c46_6 = t_r9_c46_1 + p_8_47;
  assign t_r9_c46_7 = t_r9_c46_2 + t_r9_c46_3;
  assign t_r9_c46_8 = t_r9_c46_4 + p_10_45;
  assign t_r9_c46_9 = t_r9_c46_5 + t_r9_c46_6;
  assign t_r9_c46_10 = t_r9_c46_7 + t_r9_c46_8;
  assign t_r9_c46_11 = t_r9_c46_9 + t_r9_c46_10;
  assign t_r9_c46_12 = t_r9_c46_11 + p_10_47;
  assign out_9_46 = t_r9_c46_12 >> 4;

  assign t_r9_c47_0 = p_8_47 << 1;
  assign t_r9_c47_1 = p_9_46 << 1;
  assign t_r9_c47_2 = p_9_47 << 2;
  assign t_r9_c47_3 = p_9_48 << 1;
  assign t_r9_c47_4 = p_10_47 << 1;
  assign t_r9_c47_5 = t_r9_c47_0 + p_8_46;
  assign t_r9_c47_6 = t_r9_c47_1 + p_8_48;
  assign t_r9_c47_7 = t_r9_c47_2 + t_r9_c47_3;
  assign t_r9_c47_8 = t_r9_c47_4 + p_10_46;
  assign t_r9_c47_9 = t_r9_c47_5 + t_r9_c47_6;
  assign t_r9_c47_10 = t_r9_c47_7 + t_r9_c47_8;
  assign t_r9_c47_11 = t_r9_c47_9 + t_r9_c47_10;
  assign t_r9_c47_12 = t_r9_c47_11 + p_10_48;
  assign out_9_47 = t_r9_c47_12 >> 4;

  assign t_r9_c48_0 = p_8_48 << 1;
  assign t_r9_c48_1 = p_9_47 << 1;
  assign t_r9_c48_2 = p_9_48 << 2;
  assign t_r9_c48_3 = p_9_49 << 1;
  assign t_r9_c48_4 = p_10_48 << 1;
  assign t_r9_c48_5 = t_r9_c48_0 + p_8_47;
  assign t_r9_c48_6 = t_r9_c48_1 + p_8_49;
  assign t_r9_c48_7 = t_r9_c48_2 + t_r9_c48_3;
  assign t_r9_c48_8 = t_r9_c48_4 + p_10_47;
  assign t_r9_c48_9 = t_r9_c48_5 + t_r9_c48_6;
  assign t_r9_c48_10 = t_r9_c48_7 + t_r9_c48_8;
  assign t_r9_c48_11 = t_r9_c48_9 + t_r9_c48_10;
  assign t_r9_c48_12 = t_r9_c48_11 + p_10_49;
  assign out_9_48 = t_r9_c48_12 >> 4;

  assign t_r9_c49_0 = p_8_49 << 1;
  assign t_r9_c49_1 = p_9_48 << 1;
  assign t_r9_c49_2 = p_9_49 << 2;
  assign t_r9_c49_3 = p_9_50 << 1;
  assign t_r9_c49_4 = p_10_49 << 1;
  assign t_r9_c49_5 = t_r9_c49_0 + p_8_48;
  assign t_r9_c49_6 = t_r9_c49_1 + p_8_50;
  assign t_r9_c49_7 = t_r9_c49_2 + t_r9_c49_3;
  assign t_r9_c49_8 = t_r9_c49_4 + p_10_48;
  assign t_r9_c49_9 = t_r9_c49_5 + t_r9_c49_6;
  assign t_r9_c49_10 = t_r9_c49_7 + t_r9_c49_8;
  assign t_r9_c49_11 = t_r9_c49_9 + t_r9_c49_10;
  assign t_r9_c49_12 = t_r9_c49_11 + p_10_50;
  assign out_9_49 = t_r9_c49_12 >> 4;

  assign t_r9_c50_0 = p_8_50 << 1;
  assign t_r9_c50_1 = p_9_49 << 1;
  assign t_r9_c50_2 = p_9_50 << 2;
  assign t_r9_c50_3 = p_9_51 << 1;
  assign t_r9_c50_4 = p_10_50 << 1;
  assign t_r9_c50_5 = t_r9_c50_0 + p_8_49;
  assign t_r9_c50_6 = t_r9_c50_1 + p_8_51;
  assign t_r9_c50_7 = t_r9_c50_2 + t_r9_c50_3;
  assign t_r9_c50_8 = t_r9_c50_4 + p_10_49;
  assign t_r9_c50_9 = t_r9_c50_5 + t_r9_c50_6;
  assign t_r9_c50_10 = t_r9_c50_7 + t_r9_c50_8;
  assign t_r9_c50_11 = t_r9_c50_9 + t_r9_c50_10;
  assign t_r9_c50_12 = t_r9_c50_11 + p_10_51;
  assign out_9_50 = t_r9_c50_12 >> 4;

  assign t_r9_c51_0 = p_8_51 << 1;
  assign t_r9_c51_1 = p_9_50 << 1;
  assign t_r9_c51_2 = p_9_51 << 2;
  assign t_r9_c51_3 = p_9_52 << 1;
  assign t_r9_c51_4 = p_10_51 << 1;
  assign t_r9_c51_5 = t_r9_c51_0 + p_8_50;
  assign t_r9_c51_6 = t_r9_c51_1 + p_8_52;
  assign t_r9_c51_7 = t_r9_c51_2 + t_r9_c51_3;
  assign t_r9_c51_8 = t_r9_c51_4 + p_10_50;
  assign t_r9_c51_9 = t_r9_c51_5 + t_r9_c51_6;
  assign t_r9_c51_10 = t_r9_c51_7 + t_r9_c51_8;
  assign t_r9_c51_11 = t_r9_c51_9 + t_r9_c51_10;
  assign t_r9_c51_12 = t_r9_c51_11 + p_10_52;
  assign out_9_51 = t_r9_c51_12 >> 4;

  assign t_r9_c52_0 = p_8_52 << 1;
  assign t_r9_c52_1 = p_9_51 << 1;
  assign t_r9_c52_2 = p_9_52 << 2;
  assign t_r9_c52_3 = p_9_53 << 1;
  assign t_r9_c52_4 = p_10_52 << 1;
  assign t_r9_c52_5 = t_r9_c52_0 + p_8_51;
  assign t_r9_c52_6 = t_r9_c52_1 + p_8_53;
  assign t_r9_c52_7 = t_r9_c52_2 + t_r9_c52_3;
  assign t_r9_c52_8 = t_r9_c52_4 + p_10_51;
  assign t_r9_c52_9 = t_r9_c52_5 + t_r9_c52_6;
  assign t_r9_c52_10 = t_r9_c52_7 + t_r9_c52_8;
  assign t_r9_c52_11 = t_r9_c52_9 + t_r9_c52_10;
  assign t_r9_c52_12 = t_r9_c52_11 + p_10_53;
  assign out_9_52 = t_r9_c52_12 >> 4;

  assign t_r9_c53_0 = p_8_53 << 1;
  assign t_r9_c53_1 = p_9_52 << 1;
  assign t_r9_c53_2 = p_9_53 << 2;
  assign t_r9_c53_3 = p_9_54 << 1;
  assign t_r9_c53_4 = p_10_53 << 1;
  assign t_r9_c53_5 = t_r9_c53_0 + p_8_52;
  assign t_r9_c53_6 = t_r9_c53_1 + p_8_54;
  assign t_r9_c53_7 = t_r9_c53_2 + t_r9_c53_3;
  assign t_r9_c53_8 = t_r9_c53_4 + p_10_52;
  assign t_r9_c53_9 = t_r9_c53_5 + t_r9_c53_6;
  assign t_r9_c53_10 = t_r9_c53_7 + t_r9_c53_8;
  assign t_r9_c53_11 = t_r9_c53_9 + t_r9_c53_10;
  assign t_r9_c53_12 = t_r9_c53_11 + p_10_54;
  assign out_9_53 = t_r9_c53_12 >> 4;

  assign t_r9_c54_0 = p_8_54 << 1;
  assign t_r9_c54_1 = p_9_53 << 1;
  assign t_r9_c54_2 = p_9_54 << 2;
  assign t_r9_c54_3 = p_9_55 << 1;
  assign t_r9_c54_4 = p_10_54 << 1;
  assign t_r9_c54_5 = t_r9_c54_0 + p_8_53;
  assign t_r9_c54_6 = t_r9_c54_1 + p_8_55;
  assign t_r9_c54_7 = t_r9_c54_2 + t_r9_c54_3;
  assign t_r9_c54_8 = t_r9_c54_4 + p_10_53;
  assign t_r9_c54_9 = t_r9_c54_5 + t_r9_c54_6;
  assign t_r9_c54_10 = t_r9_c54_7 + t_r9_c54_8;
  assign t_r9_c54_11 = t_r9_c54_9 + t_r9_c54_10;
  assign t_r9_c54_12 = t_r9_c54_11 + p_10_55;
  assign out_9_54 = t_r9_c54_12 >> 4;

  assign t_r9_c55_0 = p_8_55 << 1;
  assign t_r9_c55_1 = p_9_54 << 1;
  assign t_r9_c55_2 = p_9_55 << 2;
  assign t_r9_c55_3 = p_9_56 << 1;
  assign t_r9_c55_4 = p_10_55 << 1;
  assign t_r9_c55_5 = t_r9_c55_0 + p_8_54;
  assign t_r9_c55_6 = t_r9_c55_1 + p_8_56;
  assign t_r9_c55_7 = t_r9_c55_2 + t_r9_c55_3;
  assign t_r9_c55_8 = t_r9_c55_4 + p_10_54;
  assign t_r9_c55_9 = t_r9_c55_5 + t_r9_c55_6;
  assign t_r9_c55_10 = t_r9_c55_7 + t_r9_c55_8;
  assign t_r9_c55_11 = t_r9_c55_9 + t_r9_c55_10;
  assign t_r9_c55_12 = t_r9_c55_11 + p_10_56;
  assign out_9_55 = t_r9_c55_12 >> 4;

  assign t_r9_c56_0 = p_8_56 << 1;
  assign t_r9_c56_1 = p_9_55 << 1;
  assign t_r9_c56_2 = p_9_56 << 2;
  assign t_r9_c56_3 = p_9_57 << 1;
  assign t_r9_c56_4 = p_10_56 << 1;
  assign t_r9_c56_5 = t_r9_c56_0 + p_8_55;
  assign t_r9_c56_6 = t_r9_c56_1 + p_8_57;
  assign t_r9_c56_7 = t_r9_c56_2 + t_r9_c56_3;
  assign t_r9_c56_8 = t_r9_c56_4 + p_10_55;
  assign t_r9_c56_9 = t_r9_c56_5 + t_r9_c56_6;
  assign t_r9_c56_10 = t_r9_c56_7 + t_r9_c56_8;
  assign t_r9_c56_11 = t_r9_c56_9 + t_r9_c56_10;
  assign t_r9_c56_12 = t_r9_c56_11 + p_10_57;
  assign out_9_56 = t_r9_c56_12 >> 4;

  assign t_r9_c57_0 = p_8_57 << 1;
  assign t_r9_c57_1 = p_9_56 << 1;
  assign t_r9_c57_2 = p_9_57 << 2;
  assign t_r9_c57_3 = p_9_58 << 1;
  assign t_r9_c57_4 = p_10_57 << 1;
  assign t_r9_c57_5 = t_r9_c57_0 + p_8_56;
  assign t_r9_c57_6 = t_r9_c57_1 + p_8_58;
  assign t_r9_c57_7 = t_r9_c57_2 + t_r9_c57_3;
  assign t_r9_c57_8 = t_r9_c57_4 + p_10_56;
  assign t_r9_c57_9 = t_r9_c57_5 + t_r9_c57_6;
  assign t_r9_c57_10 = t_r9_c57_7 + t_r9_c57_8;
  assign t_r9_c57_11 = t_r9_c57_9 + t_r9_c57_10;
  assign t_r9_c57_12 = t_r9_c57_11 + p_10_58;
  assign out_9_57 = t_r9_c57_12 >> 4;

  assign t_r9_c58_0 = p_8_58 << 1;
  assign t_r9_c58_1 = p_9_57 << 1;
  assign t_r9_c58_2 = p_9_58 << 2;
  assign t_r9_c58_3 = p_9_59 << 1;
  assign t_r9_c58_4 = p_10_58 << 1;
  assign t_r9_c58_5 = t_r9_c58_0 + p_8_57;
  assign t_r9_c58_6 = t_r9_c58_1 + p_8_59;
  assign t_r9_c58_7 = t_r9_c58_2 + t_r9_c58_3;
  assign t_r9_c58_8 = t_r9_c58_4 + p_10_57;
  assign t_r9_c58_9 = t_r9_c58_5 + t_r9_c58_6;
  assign t_r9_c58_10 = t_r9_c58_7 + t_r9_c58_8;
  assign t_r9_c58_11 = t_r9_c58_9 + t_r9_c58_10;
  assign t_r9_c58_12 = t_r9_c58_11 + p_10_59;
  assign out_9_58 = t_r9_c58_12 >> 4;

  assign t_r9_c59_0 = p_8_59 << 1;
  assign t_r9_c59_1 = p_9_58 << 1;
  assign t_r9_c59_2 = p_9_59 << 2;
  assign t_r9_c59_3 = p_9_60 << 1;
  assign t_r9_c59_4 = p_10_59 << 1;
  assign t_r9_c59_5 = t_r9_c59_0 + p_8_58;
  assign t_r9_c59_6 = t_r9_c59_1 + p_8_60;
  assign t_r9_c59_7 = t_r9_c59_2 + t_r9_c59_3;
  assign t_r9_c59_8 = t_r9_c59_4 + p_10_58;
  assign t_r9_c59_9 = t_r9_c59_5 + t_r9_c59_6;
  assign t_r9_c59_10 = t_r9_c59_7 + t_r9_c59_8;
  assign t_r9_c59_11 = t_r9_c59_9 + t_r9_c59_10;
  assign t_r9_c59_12 = t_r9_c59_11 + p_10_60;
  assign out_9_59 = t_r9_c59_12 >> 4;

  assign t_r9_c60_0 = p_8_60 << 1;
  assign t_r9_c60_1 = p_9_59 << 1;
  assign t_r9_c60_2 = p_9_60 << 2;
  assign t_r9_c60_3 = p_9_61 << 1;
  assign t_r9_c60_4 = p_10_60 << 1;
  assign t_r9_c60_5 = t_r9_c60_0 + p_8_59;
  assign t_r9_c60_6 = t_r9_c60_1 + p_8_61;
  assign t_r9_c60_7 = t_r9_c60_2 + t_r9_c60_3;
  assign t_r9_c60_8 = t_r9_c60_4 + p_10_59;
  assign t_r9_c60_9 = t_r9_c60_5 + t_r9_c60_6;
  assign t_r9_c60_10 = t_r9_c60_7 + t_r9_c60_8;
  assign t_r9_c60_11 = t_r9_c60_9 + t_r9_c60_10;
  assign t_r9_c60_12 = t_r9_c60_11 + p_10_61;
  assign out_9_60 = t_r9_c60_12 >> 4;

  assign t_r9_c61_0 = p_8_61 << 1;
  assign t_r9_c61_1 = p_9_60 << 1;
  assign t_r9_c61_2 = p_9_61 << 2;
  assign t_r9_c61_3 = p_9_62 << 1;
  assign t_r9_c61_4 = p_10_61 << 1;
  assign t_r9_c61_5 = t_r9_c61_0 + p_8_60;
  assign t_r9_c61_6 = t_r9_c61_1 + p_8_62;
  assign t_r9_c61_7 = t_r9_c61_2 + t_r9_c61_3;
  assign t_r9_c61_8 = t_r9_c61_4 + p_10_60;
  assign t_r9_c61_9 = t_r9_c61_5 + t_r9_c61_6;
  assign t_r9_c61_10 = t_r9_c61_7 + t_r9_c61_8;
  assign t_r9_c61_11 = t_r9_c61_9 + t_r9_c61_10;
  assign t_r9_c61_12 = t_r9_c61_11 + p_10_62;
  assign out_9_61 = t_r9_c61_12 >> 4;

  assign t_r9_c62_0 = p_8_62 << 1;
  assign t_r9_c62_1 = p_9_61 << 1;
  assign t_r9_c62_2 = p_9_62 << 2;
  assign t_r9_c62_3 = p_9_63 << 1;
  assign t_r9_c62_4 = p_10_62 << 1;
  assign t_r9_c62_5 = t_r9_c62_0 + p_8_61;
  assign t_r9_c62_6 = t_r9_c62_1 + p_8_63;
  assign t_r9_c62_7 = t_r9_c62_2 + t_r9_c62_3;
  assign t_r9_c62_8 = t_r9_c62_4 + p_10_61;
  assign t_r9_c62_9 = t_r9_c62_5 + t_r9_c62_6;
  assign t_r9_c62_10 = t_r9_c62_7 + t_r9_c62_8;
  assign t_r9_c62_11 = t_r9_c62_9 + t_r9_c62_10;
  assign t_r9_c62_12 = t_r9_c62_11 + p_10_63;
  assign out_9_62 = t_r9_c62_12 >> 4;

  assign t_r9_c63_0 = p_8_63 << 1;
  assign t_r9_c63_1 = p_9_62 << 1;
  assign t_r9_c63_2 = p_9_63 << 2;
  assign t_r9_c63_3 = p_9_64 << 1;
  assign t_r9_c63_4 = p_10_63 << 1;
  assign t_r9_c63_5 = t_r9_c63_0 + p_8_62;
  assign t_r9_c63_6 = t_r9_c63_1 + p_8_64;
  assign t_r9_c63_7 = t_r9_c63_2 + t_r9_c63_3;
  assign t_r9_c63_8 = t_r9_c63_4 + p_10_62;
  assign t_r9_c63_9 = t_r9_c63_5 + t_r9_c63_6;
  assign t_r9_c63_10 = t_r9_c63_7 + t_r9_c63_8;
  assign t_r9_c63_11 = t_r9_c63_9 + t_r9_c63_10;
  assign t_r9_c63_12 = t_r9_c63_11 + p_10_64;
  assign out_9_63 = t_r9_c63_12 >> 4;

  assign t_r9_c64_0 = p_8_64 << 1;
  assign t_r9_c64_1 = p_9_63 << 1;
  assign t_r9_c64_2 = p_9_64 << 2;
  assign t_r9_c64_3 = p_9_65 << 1;
  assign t_r9_c64_4 = p_10_64 << 1;
  assign t_r9_c64_5 = t_r9_c64_0 + p_8_63;
  assign t_r9_c64_6 = t_r9_c64_1 + p_8_65;
  assign t_r9_c64_7 = t_r9_c64_2 + t_r9_c64_3;
  assign t_r9_c64_8 = t_r9_c64_4 + p_10_63;
  assign t_r9_c64_9 = t_r9_c64_5 + t_r9_c64_6;
  assign t_r9_c64_10 = t_r9_c64_7 + t_r9_c64_8;
  assign t_r9_c64_11 = t_r9_c64_9 + t_r9_c64_10;
  assign t_r9_c64_12 = t_r9_c64_11 + p_10_65;
  assign out_9_64 = t_r9_c64_12 >> 4;

  assign t_r10_c1_0 = p_9_1 << 1;
  assign t_r10_c1_1 = p_10_0 << 1;
  assign t_r10_c1_2 = p_10_1 << 2;
  assign t_r10_c1_3 = p_10_2 << 1;
  assign t_r10_c1_4 = p_11_1 << 1;
  assign t_r10_c1_5 = t_r10_c1_0 + p_9_0;
  assign t_r10_c1_6 = t_r10_c1_1 + p_9_2;
  assign t_r10_c1_7 = t_r10_c1_2 + t_r10_c1_3;
  assign t_r10_c1_8 = t_r10_c1_4 + p_11_0;
  assign t_r10_c1_9 = t_r10_c1_5 + t_r10_c1_6;
  assign t_r10_c1_10 = t_r10_c1_7 + t_r10_c1_8;
  assign t_r10_c1_11 = t_r10_c1_9 + t_r10_c1_10;
  assign t_r10_c1_12 = t_r10_c1_11 + p_11_2;
  assign out_10_1 = t_r10_c1_12 >> 4;

  assign t_r10_c2_0 = p_9_2 << 1;
  assign t_r10_c2_1 = p_10_1 << 1;
  assign t_r10_c2_2 = p_10_2 << 2;
  assign t_r10_c2_3 = p_10_3 << 1;
  assign t_r10_c2_4 = p_11_2 << 1;
  assign t_r10_c2_5 = t_r10_c2_0 + p_9_1;
  assign t_r10_c2_6 = t_r10_c2_1 + p_9_3;
  assign t_r10_c2_7 = t_r10_c2_2 + t_r10_c2_3;
  assign t_r10_c2_8 = t_r10_c2_4 + p_11_1;
  assign t_r10_c2_9 = t_r10_c2_5 + t_r10_c2_6;
  assign t_r10_c2_10 = t_r10_c2_7 + t_r10_c2_8;
  assign t_r10_c2_11 = t_r10_c2_9 + t_r10_c2_10;
  assign t_r10_c2_12 = t_r10_c2_11 + p_11_3;
  assign out_10_2 = t_r10_c2_12 >> 4;

  assign t_r10_c3_0 = p_9_3 << 1;
  assign t_r10_c3_1 = p_10_2 << 1;
  assign t_r10_c3_2 = p_10_3 << 2;
  assign t_r10_c3_3 = p_10_4 << 1;
  assign t_r10_c3_4 = p_11_3 << 1;
  assign t_r10_c3_5 = t_r10_c3_0 + p_9_2;
  assign t_r10_c3_6 = t_r10_c3_1 + p_9_4;
  assign t_r10_c3_7 = t_r10_c3_2 + t_r10_c3_3;
  assign t_r10_c3_8 = t_r10_c3_4 + p_11_2;
  assign t_r10_c3_9 = t_r10_c3_5 + t_r10_c3_6;
  assign t_r10_c3_10 = t_r10_c3_7 + t_r10_c3_8;
  assign t_r10_c3_11 = t_r10_c3_9 + t_r10_c3_10;
  assign t_r10_c3_12 = t_r10_c3_11 + p_11_4;
  assign out_10_3 = t_r10_c3_12 >> 4;

  assign t_r10_c4_0 = p_9_4 << 1;
  assign t_r10_c4_1 = p_10_3 << 1;
  assign t_r10_c4_2 = p_10_4 << 2;
  assign t_r10_c4_3 = p_10_5 << 1;
  assign t_r10_c4_4 = p_11_4 << 1;
  assign t_r10_c4_5 = t_r10_c4_0 + p_9_3;
  assign t_r10_c4_6 = t_r10_c4_1 + p_9_5;
  assign t_r10_c4_7 = t_r10_c4_2 + t_r10_c4_3;
  assign t_r10_c4_8 = t_r10_c4_4 + p_11_3;
  assign t_r10_c4_9 = t_r10_c4_5 + t_r10_c4_6;
  assign t_r10_c4_10 = t_r10_c4_7 + t_r10_c4_8;
  assign t_r10_c4_11 = t_r10_c4_9 + t_r10_c4_10;
  assign t_r10_c4_12 = t_r10_c4_11 + p_11_5;
  assign out_10_4 = t_r10_c4_12 >> 4;

  assign t_r10_c5_0 = p_9_5 << 1;
  assign t_r10_c5_1 = p_10_4 << 1;
  assign t_r10_c5_2 = p_10_5 << 2;
  assign t_r10_c5_3 = p_10_6 << 1;
  assign t_r10_c5_4 = p_11_5 << 1;
  assign t_r10_c5_5 = t_r10_c5_0 + p_9_4;
  assign t_r10_c5_6 = t_r10_c5_1 + p_9_6;
  assign t_r10_c5_7 = t_r10_c5_2 + t_r10_c5_3;
  assign t_r10_c5_8 = t_r10_c5_4 + p_11_4;
  assign t_r10_c5_9 = t_r10_c5_5 + t_r10_c5_6;
  assign t_r10_c5_10 = t_r10_c5_7 + t_r10_c5_8;
  assign t_r10_c5_11 = t_r10_c5_9 + t_r10_c5_10;
  assign t_r10_c5_12 = t_r10_c5_11 + p_11_6;
  assign out_10_5 = t_r10_c5_12 >> 4;

  assign t_r10_c6_0 = p_9_6 << 1;
  assign t_r10_c6_1 = p_10_5 << 1;
  assign t_r10_c6_2 = p_10_6 << 2;
  assign t_r10_c6_3 = p_10_7 << 1;
  assign t_r10_c6_4 = p_11_6 << 1;
  assign t_r10_c6_5 = t_r10_c6_0 + p_9_5;
  assign t_r10_c6_6 = t_r10_c6_1 + p_9_7;
  assign t_r10_c6_7 = t_r10_c6_2 + t_r10_c6_3;
  assign t_r10_c6_8 = t_r10_c6_4 + p_11_5;
  assign t_r10_c6_9 = t_r10_c6_5 + t_r10_c6_6;
  assign t_r10_c6_10 = t_r10_c6_7 + t_r10_c6_8;
  assign t_r10_c6_11 = t_r10_c6_9 + t_r10_c6_10;
  assign t_r10_c6_12 = t_r10_c6_11 + p_11_7;
  assign out_10_6 = t_r10_c6_12 >> 4;

  assign t_r10_c7_0 = p_9_7 << 1;
  assign t_r10_c7_1 = p_10_6 << 1;
  assign t_r10_c7_2 = p_10_7 << 2;
  assign t_r10_c7_3 = p_10_8 << 1;
  assign t_r10_c7_4 = p_11_7 << 1;
  assign t_r10_c7_5 = t_r10_c7_0 + p_9_6;
  assign t_r10_c7_6 = t_r10_c7_1 + p_9_8;
  assign t_r10_c7_7 = t_r10_c7_2 + t_r10_c7_3;
  assign t_r10_c7_8 = t_r10_c7_4 + p_11_6;
  assign t_r10_c7_9 = t_r10_c7_5 + t_r10_c7_6;
  assign t_r10_c7_10 = t_r10_c7_7 + t_r10_c7_8;
  assign t_r10_c7_11 = t_r10_c7_9 + t_r10_c7_10;
  assign t_r10_c7_12 = t_r10_c7_11 + p_11_8;
  assign out_10_7 = t_r10_c7_12 >> 4;

  assign t_r10_c8_0 = p_9_8 << 1;
  assign t_r10_c8_1 = p_10_7 << 1;
  assign t_r10_c8_2 = p_10_8 << 2;
  assign t_r10_c8_3 = p_10_9 << 1;
  assign t_r10_c8_4 = p_11_8 << 1;
  assign t_r10_c8_5 = t_r10_c8_0 + p_9_7;
  assign t_r10_c8_6 = t_r10_c8_1 + p_9_9;
  assign t_r10_c8_7 = t_r10_c8_2 + t_r10_c8_3;
  assign t_r10_c8_8 = t_r10_c8_4 + p_11_7;
  assign t_r10_c8_9 = t_r10_c8_5 + t_r10_c8_6;
  assign t_r10_c8_10 = t_r10_c8_7 + t_r10_c8_8;
  assign t_r10_c8_11 = t_r10_c8_9 + t_r10_c8_10;
  assign t_r10_c8_12 = t_r10_c8_11 + p_11_9;
  assign out_10_8 = t_r10_c8_12 >> 4;

  assign t_r10_c9_0 = p_9_9 << 1;
  assign t_r10_c9_1 = p_10_8 << 1;
  assign t_r10_c9_2 = p_10_9 << 2;
  assign t_r10_c9_3 = p_10_10 << 1;
  assign t_r10_c9_4 = p_11_9 << 1;
  assign t_r10_c9_5 = t_r10_c9_0 + p_9_8;
  assign t_r10_c9_6 = t_r10_c9_1 + p_9_10;
  assign t_r10_c9_7 = t_r10_c9_2 + t_r10_c9_3;
  assign t_r10_c9_8 = t_r10_c9_4 + p_11_8;
  assign t_r10_c9_9 = t_r10_c9_5 + t_r10_c9_6;
  assign t_r10_c9_10 = t_r10_c9_7 + t_r10_c9_8;
  assign t_r10_c9_11 = t_r10_c9_9 + t_r10_c9_10;
  assign t_r10_c9_12 = t_r10_c9_11 + p_11_10;
  assign out_10_9 = t_r10_c9_12 >> 4;

  assign t_r10_c10_0 = p_9_10 << 1;
  assign t_r10_c10_1 = p_10_9 << 1;
  assign t_r10_c10_2 = p_10_10 << 2;
  assign t_r10_c10_3 = p_10_11 << 1;
  assign t_r10_c10_4 = p_11_10 << 1;
  assign t_r10_c10_5 = t_r10_c10_0 + p_9_9;
  assign t_r10_c10_6 = t_r10_c10_1 + p_9_11;
  assign t_r10_c10_7 = t_r10_c10_2 + t_r10_c10_3;
  assign t_r10_c10_8 = t_r10_c10_4 + p_11_9;
  assign t_r10_c10_9 = t_r10_c10_5 + t_r10_c10_6;
  assign t_r10_c10_10 = t_r10_c10_7 + t_r10_c10_8;
  assign t_r10_c10_11 = t_r10_c10_9 + t_r10_c10_10;
  assign t_r10_c10_12 = t_r10_c10_11 + p_11_11;
  assign out_10_10 = t_r10_c10_12 >> 4;

  assign t_r10_c11_0 = p_9_11 << 1;
  assign t_r10_c11_1 = p_10_10 << 1;
  assign t_r10_c11_2 = p_10_11 << 2;
  assign t_r10_c11_3 = p_10_12 << 1;
  assign t_r10_c11_4 = p_11_11 << 1;
  assign t_r10_c11_5 = t_r10_c11_0 + p_9_10;
  assign t_r10_c11_6 = t_r10_c11_1 + p_9_12;
  assign t_r10_c11_7 = t_r10_c11_2 + t_r10_c11_3;
  assign t_r10_c11_8 = t_r10_c11_4 + p_11_10;
  assign t_r10_c11_9 = t_r10_c11_5 + t_r10_c11_6;
  assign t_r10_c11_10 = t_r10_c11_7 + t_r10_c11_8;
  assign t_r10_c11_11 = t_r10_c11_9 + t_r10_c11_10;
  assign t_r10_c11_12 = t_r10_c11_11 + p_11_12;
  assign out_10_11 = t_r10_c11_12 >> 4;

  assign t_r10_c12_0 = p_9_12 << 1;
  assign t_r10_c12_1 = p_10_11 << 1;
  assign t_r10_c12_2 = p_10_12 << 2;
  assign t_r10_c12_3 = p_10_13 << 1;
  assign t_r10_c12_4 = p_11_12 << 1;
  assign t_r10_c12_5 = t_r10_c12_0 + p_9_11;
  assign t_r10_c12_6 = t_r10_c12_1 + p_9_13;
  assign t_r10_c12_7 = t_r10_c12_2 + t_r10_c12_3;
  assign t_r10_c12_8 = t_r10_c12_4 + p_11_11;
  assign t_r10_c12_9 = t_r10_c12_5 + t_r10_c12_6;
  assign t_r10_c12_10 = t_r10_c12_7 + t_r10_c12_8;
  assign t_r10_c12_11 = t_r10_c12_9 + t_r10_c12_10;
  assign t_r10_c12_12 = t_r10_c12_11 + p_11_13;
  assign out_10_12 = t_r10_c12_12 >> 4;

  assign t_r10_c13_0 = p_9_13 << 1;
  assign t_r10_c13_1 = p_10_12 << 1;
  assign t_r10_c13_2 = p_10_13 << 2;
  assign t_r10_c13_3 = p_10_14 << 1;
  assign t_r10_c13_4 = p_11_13 << 1;
  assign t_r10_c13_5 = t_r10_c13_0 + p_9_12;
  assign t_r10_c13_6 = t_r10_c13_1 + p_9_14;
  assign t_r10_c13_7 = t_r10_c13_2 + t_r10_c13_3;
  assign t_r10_c13_8 = t_r10_c13_4 + p_11_12;
  assign t_r10_c13_9 = t_r10_c13_5 + t_r10_c13_6;
  assign t_r10_c13_10 = t_r10_c13_7 + t_r10_c13_8;
  assign t_r10_c13_11 = t_r10_c13_9 + t_r10_c13_10;
  assign t_r10_c13_12 = t_r10_c13_11 + p_11_14;
  assign out_10_13 = t_r10_c13_12 >> 4;

  assign t_r10_c14_0 = p_9_14 << 1;
  assign t_r10_c14_1 = p_10_13 << 1;
  assign t_r10_c14_2 = p_10_14 << 2;
  assign t_r10_c14_3 = p_10_15 << 1;
  assign t_r10_c14_4 = p_11_14 << 1;
  assign t_r10_c14_5 = t_r10_c14_0 + p_9_13;
  assign t_r10_c14_6 = t_r10_c14_1 + p_9_15;
  assign t_r10_c14_7 = t_r10_c14_2 + t_r10_c14_3;
  assign t_r10_c14_8 = t_r10_c14_4 + p_11_13;
  assign t_r10_c14_9 = t_r10_c14_5 + t_r10_c14_6;
  assign t_r10_c14_10 = t_r10_c14_7 + t_r10_c14_8;
  assign t_r10_c14_11 = t_r10_c14_9 + t_r10_c14_10;
  assign t_r10_c14_12 = t_r10_c14_11 + p_11_15;
  assign out_10_14 = t_r10_c14_12 >> 4;

  assign t_r10_c15_0 = p_9_15 << 1;
  assign t_r10_c15_1 = p_10_14 << 1;
  assign t_r10_c15_2 = p_10_15 << 2;
  assign t_r10_c15_3 = p_10_16 << 1;
  assign t_r10_c15_4 = p_11_15 << 1;
  assign t_r10_c15_5 = t_r10_c15_0 + p_9_14;
  assign t_r10_c15_6 = t_r10_c15_1 + p_9_16;
  assign t_r10_c15_7 = t_r10_c15_2 + t_r10_c15_3;
  assign t_r10_c15_8 = t_r10_c15_4 + p_11_14;
  assign t_r10_c15_9 = t_r10_c15_5 + t_r10_c15_6;
  assign t_r10_c15_10 = t_r10_c15_7 + t_r10_c15_8;
  assign t_r10_c15_11 = t_r10_c15_9 + t_r10_c15_10;
  assign t_r10_c15_12 = t_r10_c15_11 + p_11_16;
  assign out_10_15 = t_r10_c15_12 >> 4;

  assign t_r10_c16_0 = p_9_16 << 1;
  assign t_r10_c16_1 = p_10_15 << 1;
  assign t_r10_c16_2 = p_10_16 << 2;
  assign t_r10_c16_3 = p_10_17 << 1;
  assign t_r10_c16_4 = p_11_16 << 1;
  assign t_r10_c16_5 = t_r10_c16_0 + p_9_15;
  assign t_r10_c16_6 = t_r10_c16_1 + p_9_17;
  assign t_r10_c16_7 = t_r10_c16_2 + t_r10_c16_3;
  assign t_r10_c16_8 = t_r10_c16_4 + p_11_15;
  assign t_r10_c16_9 = t_r10_c16_5 + t_r10_c16_6;
  assign t_r10_c16_10 = t_r10_c16_7 + t_r10_c16_8;
  assign t_r10_c16_11 = t_r10_c16_9 + t_r10_c16_10;
  assign t_r10_c16_12 = t_r10_c16_11 + p_11_17;
  assign out_10_16 = t_r10_c16_12 >> 4;

  assign t_r10_c17_0 = p_9_17 << 1;
  assign t_r10_c17_1 = p_10_16 << 1;
  assign t_r10_c17_2 = p_10_17 << 2;
  assign t_r10_c17_3 = p_10_18 << 1;
  assign t_r10_c17_4 = p_11_17 << 1;
  assign t_r10_c17_5 = t_r10_c17_0 + p_9_16;
  assign t_r10_c17_6 = t_r10_c17_1 + p_9_18;
  assign t_r10_c17_7 = t_r10_c17_2 + t_r10_c17_3;
  assign t_r10_c17_8 = t_r10_c17_4 + p_11_16;
  assign t_r10_c17_9 = t_r10_c17_5 + t_r10_c17_6;
  assign t_r10_c17_10 = t_r10_c17_7 + t_r10_c17_8;
  assign t_r10_c17_11 = t_r10_c17_9 + t_r10_c17_10;
  assign t_r10_c17_12 = t_r10_c17_11 + p_11_18;
  assign out_10_17 = t_r10_c17_12 >> 4;

  assign t_r10_c18_0 = p_9_18 << 1;
  assign t_r10_c18_1 = p_10_17 << 1;
  assign t_r10_c18_2 = p_10_18 << 2;
  assign t_r10_c18_3 = p_10_19 << 1;
  assign t_r10_c18_4 = p_11_18 << 1;
  assign t_r10_c18_5 = t_r10_c18_0 + p_9_17;
  assign t_r10_c18_6 = t_r10_c18_1 + p_9_19;
  assign t_r10_c18_7 = t_r10_c18_2 + t_r10_c18_3;
  assign t_r10_c18_8 = t_r10_c18_4 + p_11_17;
  assign t_r10_c18_9 = t_r10_c18_5 + t_r10_c18_6;
  assign t_r10_c18_10 = t_r10_c18_7 + t_r10_c18_8;
  assign t_r10_c18_11 = t_r10_c18_9 + t_r10_c18_10;
  assign t_r10_c18_12 = t_r10_c18_11 + p_11_19;
  assign out_10_18 = t_r10_c18_12 >> 4;

  assign t_r10_c19_0 = p_9_19 << 1;
  assign t_r10_c19_1 = p_10_18 << 1;
  assign t_r10_c19_2 = p_10_19 << 2;
  assign t_r10_c19_3 = p_10_20 << 1;
  assign t_r10_c19_4 = p_11_19 << 1;
  assign t_r10_c19_5 = t_r10_c19_0 + p_9_18;
  assign t_r10_c19_6 = t_r10_c19_1 + p_9_20;
  assign t_r10_c19_7 = t_r10_c19_2 + t_r10_c19_3;
  assign t_r10_c19_8 = t_r10_c19_4 + p_11_18;
  assign t_r10_c19_9 = t_r10_c19_5 + t_r10_c19_6;
  assign t_r10_c19_10 = t_r10_c19_7 + t_r10_c19_8;
  assign t_r10_c19_11 = t_r10_c19_9 + t_r10_c19_10;
  assign t_r10_c19_12 = t_r10_c19_11 + p_11_20;
  assign out_10_19 = t_r10_c19_12 >> 4;

  assign t_r10_c20_0 = p_9_20 << 1;
  assign t_r10_c20_1 = p_10_19 << 1;
  assign t_r10_c20_2 = p_10_20 << 2;
  assign t_r10_c20_3 = p_10_21 << 1;
  assign t_r10_c20_4 = p_11_20 << 1;
  assign t_r10_c20_5 = t_r10_c20_0 + p_9_19;
  assign t_r10_c20_6 = t_r10_c20_1 + p_9_21;
  assign t_r10_c20_7 = t_r10_c20_2 + t_r10_c20_3;
  assign t_r10_c20_8 = t_r10_c20_4 + p_11_19;
  assign t_r10_c20_9 = t_r10_c20_5 + t_r10_c20_6;
  assign t_r10_c20_10 = t_r10_c20_7 + t_r10_c20_8;
  assign t_r10_c20_11 = t_r10_c20_9 + t_r10_c20_10;
  assign t_r10_c20_12 = t_r10_c20_11 + p_11_21;
  assign out_10_20 = t_r10_c20_12 >> 4;

  assign t_r10_c21_0 = p_9_21 << 1;
  assign t_r10_c21_1 = p_10_20 << 1;
  assign t_r10_c21_2 = p_10_21 << 2;
  assign t_r10_c21_3 = p_10_22 << 1;
  assign t_r10_c21_4 = p_11_21 << 1;
  assign t_r10_c21_5 = t_r10_c21_0 + p_9_20;
  assign t_r10_c21_6 = t_r10_c21_1 + p_9_22;
  assign t_r10_c21_7 = t_r10_c21_2 + t_r10_c21_3;
  assign t_r10_c21_8 = t_r10_c21_4 + p_11_20;
  assign t_r10_c21_9 = t_r10_c21_5 + t_r10_c21_6;
  assign t_r10_c21_10 = t_r10_c21_7 + t_r10_c21_8;
  assign t_r10_c21_11 = t_r10_c21_9 + t_r10_c21_10;
  assign t_r10_c21_12 = t_r10_c21_11 + p_11_22;
  assign out_10_21 = t_r10_c21_12 >> 4;

  assign t_r10_c22_0 = p_9_22 << 1;
  assign t_r10_c22_1 = p_10_21 << 1;
  assign t_r10_c22_2 = p_10_22 << 2;
  assign t_r10_c22_3 = p_10_23 << 1;
  assign t_r10_c22_4 = p_11_22 << 1;
  assign t_r10_c22_5 = t_r10_c22_0 + p_9_21;
  assign t_r10_c22_6 = t_r10_c22_1 + p_9_23;
  assign t_r10_c22_7 = t_r10_c22_2 + t_r10_c22_3;
  assign t_r10_c22_8 = t_r10_c22_4 + p_11_21;
  assign t_r10_c22_9 = t_r10_c22_5 + t_r10_c22_6;
  assign t_r10_c22_10 = t_r10_c22_7 + t_r10_c22_8;
  assign t_r10_c22_11 = t_r10_c22_9 + t_r10_c22_10;
  assign t_r10_c22_12 = t_r10_c22_11 + p_11_23;
  assign out_10_22 = t_r10_c22_12 >> 4;

  assign t_r10_c23_0 = p_9_23 << 1;
  assign t_r10_c23_1 = p_10_22 << 1;
  assign t_r10_c23_2 = p_10_23 << 2;
  assign t_r10_c23_3 = p_10_24 << 1;
  assign t_r10_c23_4 = p_11_23 << 1;
  assign t_r10_c23_5 = t_r10_c23_0 + p_9_22;
  assign t_r10_c23_6 = t_r10_c23_1 + p_9_24;
  assign t_r10_c23_7 = t_r10_c23_2 + t_r10_c23_3;
  assign t_r10_c23_8 = t_r10_c23_4 + p_11_22;
  assign t_r10_c23_9 = t_r10_c23_5 + t_r10_c23_6;
  assign t_r10_c23_10 = t_r10_c23_7 + t_r10_c23_8;
  assign t_r10_c23_11 = t_r10_c23_9 + t_r10_c23_10;
  assign t_r10_c23_12 = t_r10_c23_11 + p_11_24;
  assign out_10_23 = t_r10_c23_12 >> 4;

  assign t_r10_c24_0 = p_9_24 << 1;
  assign t_r10_c24_1 = p_10_23 << 1;
  assign t_r10_c24_2 = p_10_24 << 2;
  assign t_r10_c24_3 = p_10_25 << 1;
  assign t_r10_c24_4 = p_11_24 << 1;
  assign t_r10_c24_5 = t_r10_c24_0 + p_9_23;
  assign t_r10_c24_6 = t_r10_c24_1 + p_9_25;
  assign t_r10_c24_7 = t_r10_c24_2 + t_r10_c24_3;
  assign t_r10_c24_8 = t_r10_c24_4 + p_11_23;
  assign t_r10_c24_9 = t_r10_c24_5 + t_r10_c24_6;
  assign t_r10_c24_10 = t_r10_c24_7 + t_r10_c24_8;
  assign t_r10_c24_11 = t_r10_c24_9 + t_r10_c24_10;
  assign t_r10_c24_12 = t_r10_c24_11 + p_11_25;
  assign out_10_24 = t_r10_c24_12 >> 4;

  assign t_r10_c25_0 = p_9_25 << 1;
  assign t_r10_c25_1 = p_10_24 << 1;
  assign t_r10_c25_2 = p_10_25 << 2;
  assign t_r10_c25_3 = p_10_26 << 1;
  assign t_r10_c25_4 = p_11_25 << 1;
  assign t_r10_c25_5 = t_r10_c25_0 + p_9_24;
  assign t_r10_c25_6 = t_r10_c25_1 + p_9_26;
  assign t_r10_c25_7 = t_r10_c25_2 + t_r10_c25_3;
  assign t_r10_c25_8 = t_r10_c25_4 + p_11_24;
  assign t_r10_c25_9 = t_r10_c25_5 + t_r10_c25_6;
  assign t_r10_c25_10 = t_r10_c25_7 + t_r10_c25_8;
  assign t_r10_c25_11 = t_r10_c25_9 + t_r10_c25_10;
  assign t_r10_c25_12 = t_r10_c25_11 + p_11_26;
  assign out_10_25 = t_r10_c25_12 >> 4;

  assign t_r10_c26_0 = p_9_26 << 1;
  assign t_r10_c26_1 = p_10_25 << 1;
  assign t_r10_c26_2 = p_10_26 << 2;
  assign t_r10_c26_3 = p_10_27 << 1;
  assign t_r10_c26_4 = p_11_26 << 1;
  assign t_r10_c26_5 = t_r10_c26_0 + p_9_25;
  assign t_r10_c26_6 = t_r10_c26_1 + p_9_27;
  assign t_r10_c26_7 = t_r10_c26_2 + t_r10_c26_3;
  assign t_r10_c26_8 = t_r10_c26_4 + p_11_25;
  assign t_r10_c26_9 = t_r10_c26_5 + t_r10_c26_6;
  assign t_r10_c26_10 = t_r10_c26_7 + t_r10_c26_8;
  assign t_r10_c26_11 = t_r10_c26_9 + t_r10_c26_10;
  assign t_r10_c26_12 = t_r10_c26_11 + p_11_27;
  assign out_10_26 = t_r10_c26_12 >> 4;

  assign t_r10_c27_0 = p_9_27 << 1;
  assign t_r10_c27_1 = p_10_26 << 1;
  assign t_r10_c27_2 = p_10_27 << 2;
  assign t_r10_c27_3 = p_10_28 << 1;
  assign t_r10_c27_4 = p_11_27 << 1;
  assign t_r10_c27_5 = t_r10_c27_0 + p_9_26;
  assign t_r10_c27_6 = t_r10_c27_1 + p_9_28;
  assign t_r10_c27_7 = t_r10_c27_2 + t_r10_c27_3;
  assign t_r10_c27_8 = t_r10_c27_4 + p_11_26;
  assign t_r10_c27_9 = t_r10_c27_5 + t_r10_c27_6;
  assign t_r10_c27_10 = t_r10_c27_7 + t_r10_c27_8;
  assign t_r10_c27_11 = t_r10_c27_9 + t_r10_c27_10;
  assign t_r10_c27_12 = t_r10_c27_11 + p_11_28;
  assign out_10_27 = t_r10_c27_12 >> 4;

  assign t_r10_c28_0 = p_9_28 << 1;
  assign t_r10_c28_1 = p_10_27 << 1;
  assign t_r10_c28_2 = p_10_28 << 2;
  assign t_r10_c28_3 = p_10_29 << 1;
  assign t_r10_c28_4 = p_11_28 << 1;
  assign t_r10_c28_5 = t_r10_c28_0 + p_9_27;
  assign t_r10_c28_6 = t_r10_c28_1 + p_9_29;
  assign t_r10_c28_7 = t_r10_c28_2 + t_r10_c28_3;
  assign t_r10_c28_8 = t_r10_c28_4 + p_11_27;
  assign t_r10_c28_9 = t_r10_c28_5 + t_r10_c28_6;
  assign t_r10_c28_10 = t_r10_c28_7 + t_r10_c28_8;
  assign t_r10_c28_11 = t_r10_c28_9 + t_r10_c28_10;
  assign t_r10_c28_12 = t_r10_c28_11 + p_11_29;
  assign out_10_28 = t_r10_c28_12 >> 4;

  assign t_r10_c29_0 = p_9_29 << 1;
  assign t_r10_c29_1 = p_10_28 << 1;
  assign t_r10_c29_2 = p_10_29 << 2;
  assign t_r10_c29_3 = p_10_30 << 1;
  assign t_r10_c29_4 = p_11_29 << 1;
  assign t_r10_c29_5 = t_r10_c29_0 + p_9_28;
  assign t_r10_c29_6 = t_r10_c29_1 + p_9_30;
  assign t_r10_c29_7 = t_r10_c29_2 + t_r10_c29_3;
  assign t_r10_c29_8 = t_r10_c29_4 + p_11_28;
  assign t_r10_c29_9 = t_r10_c29_5 + t_r10_c29_6;
  assign t_r10_c29_10 = t_r10_c29_7 + t_r10_c29_8;
  assign t_r10_c29_11 = t_r10_c29_9 + t_r10_c29_10;
  assign t_r10_c29_12 = t_r10_c29_11 + p_11_30;
  assign out_10_29 = t_r10_c29_12 >> 4;

  assign t_r10_c30_0 = p_9_30 << 1;
  assign t_r10_c30_1 = p_10_29 << 1;
  assign t_r10_c30_2 = p_10_30 << 2;
  assign t_r10_c30_3 = p_10_31 << 1;
  assign t_r10_c30_4 = p_11_30 << 1;
  assign t_r10_c30_5 = t_r10_c30_0 + p_9_29;
  assign t_r10_c30_6 = t_r10_c30_1 + p_9_31;
  assign t_r10_c30_7 = t_r10_c30_2 + t_r10_c30_3;
  assign t_r10_c30_8 = t_r10_c30_4 + p_11_29;
  assign t_r10_c30_9 = t_r10_c30_5 + t_r10_c30_6;
  assign t_r10_c30_10 = t_r10_c30_7 + t_r10_c30_8;
  assign t_r10_c30_11 = t_r10_c30_9 + t_r10_c30_10;
  assign t_r10_c30_12 = t_r10_c30_11 + p_11_31;
  assign out_10_30 = t_r10_c30_12 >> 4;

  assign t_r10_c31_0 = p_9_31 << 1;
  assign t_r10_c31_1 = p_10_30 << 1;
  assign t_r10_c31_2 = p_10_31 << 2;
  assign t_r10_c31_3 = p_10_32 << 1;
  assign t_r10_c31_4 = p_11_31 << 1;
  assign t_r10_c31_5 = t_r10_c31_0 + p_9_30;
  assign t_r10_c31_6 = t_r10_c31_1 + p_9_32;
  assign t_r10_c31_7 = t_r10_c31_2 + t_r10_c31_3;
  assign t_r10_c31_8 = t_r10_c31_4 + p_11_30;
  assign t_r10_c31_9 = t_r10_c31_5 + t_r10_c31_6;
  assign t_r10_c31_10 = t_r10_c31_7 + t_r10_c31_8;
  assign t_r10_c31_11 = t_r10_c31_9 + t_r10_c31_10;
  assign t_r10_c31_12 = t_r10_c31_11 + p_11_32;
  assign out_10_31 = t_r10_c31_12 >> 4;

  assign t_r10_c32_0 = p_9_32 << 1;
  assign t_r10_c32_1 = p_10_31 << 1;
  assign t_r10_c32_2 = p_10_32 << 2;
  assign t_r10_c32_3 = p_10_33 << 1;
  assign t_r10_c32_4 = p_11_32 << 1;
  assign t_r10_c32_5 = t_r10_c32_0 + p_9_31;
  assign t_r10_c32_6 = t_r10_c32_1 + p_9_33;
  assign t_r10_c32_7 = t_r10_c32_2 + t_r10_c32_3;
  assign t_r10_c32_8 = t_r10_c32_4 + p_11_31;
  assign t_r10_c32_9 = t_r10_c32_5 + t_r10_c32_6;
  assign t_r10_c32_10 = t_r10_c32_7 + t_r10_c32_8;
  assign t_r10_c32_11 = t_r10_c32_9 + t_r10_c32_10;
  assign t_r10_c32_12 = t_r10_c32_11 + p_11_33;
  assign out_10_32 = t_r10_c32_12 >> 4;

  assign t_r10_c33_0 = p_9_33 << 1;
  assign t_r10_c33_1 = p_10_32 << 1;
  assign t_r10_c33_2 = p_10_33 << 2;
  assign t_r10_c33_3 = p_10_34 << 1;
  assign t_r10_c33_4 = p_11_33 << 1;
  assign t_r10_c33_5 = t_r10_c33_0 + p_9_32;
  assign t_r10_c33_6 = t_r10_c33_1 + p_9_34;
  assign t_r10_c33_7 = t_r10_c33_2 + t_r10_c33_3;
  assign t_r10_c33_8 = t_r10_c33_4 + p_11_32;
  assign t_r10_c33_9 = t_r10_c33_5 + t_r10_c33_6;
  assign t_r10_c33_10 = t_r10_c33_7 + t_r10_c33_8;
  assign t_r10_c33_11 = t_r10_c33_9 + t_r10_c33_10;
  assign t_r10_c33_12 = t_r10_c33_11 + p_11_34;
  assign out_10_33 = t_r10_c33_12 >> 4;

  assign t_r10_c34_0 = p_9_34 << 1;
  assign t_r10_c34_1 = p_10_33 << 1;
  assign t_r10_c34_2 = p_10_34 << 2;
  assign t_r10_c34_3 = p_10_35 << 1;
  assign t_r10_c34_4 = p_11_34 << 1;
  assign t_r10_c34_5 = t_r10_c34_0 + p_9_33;
  assign t_r10_c34_6 = t_r10_c34_1 + p_9_35;
  assign t_r10_c34_7 = t_r10_c34_2 + t_r10_c34_3;
  assign t_r10_c34_8 = t_r10_c34_4 + p_11_33;
  assign t_r10_c34_9 = t_r10_c34_5 + t_r10_c34_6;
  assign t_r10_c34_10 = t_r10_c34_7 + t_r10_c34_8;
  assign t_r10_c34_11 = t_r10_c34_9 + t_r10_c34_10;
  assign t_r10_c34_12 = t_r10_c34_11 + p_11_35;
  assign out_10_34 = t_r10_c34_12 >> 4;

  assign t_r10_c35_0 = p_9_35 << 1;
  assign t_r10_c35_1 = p_10_34 << 1;
  assign t_r10_c35_2 = p_10_35 << 2;
  assign t_r10_c35_3 = p_10_36 << 1;
  assign t_r10_c35_4 = p_11_35 << 1;
  assign t_r10_c35_5 = t_r10_c35_0 + p_9_34;
  assign t_r10_c35_6 = t_r10_c35_1 + p_9_36;
  assign t_r10_c35_7 = t_r10_c35_2 + t_r10_c35_3;
  assign t_r10_c35_8 = t_r10_c35_4 + p_11_34;
  assign t_r10_c35_9 = t_r10_c35_5 + t_r10_c35_6;
  assign t_r10_c35_10 = t_r10_c35_7 + t_r10_c35_8;
  assign t_r10_c35_11 = t_r10_c35_9 + t_r10_c35_10;
  assign t_r10_c35_12 = t_r10_c35_11 + p_11_36;
  assign out_10_35 = t_r10_c35_12 >> 4;

  assign t_r10_c36_0 = p_9_36 << 1;
  assign t_r10_c36_1 = p_10_35 << 1;
  assign t_r10_c36_2 = p_10_36 << 2;
  assign t_r10_c36_3 = p_10_37 << 1;
  assign t_r10_c36_4 = p_11_36 << 1;
  assign t_r10_c36_5 = t_r10_c36_0 + p_9_35;
  assign t_r10_c36_6 = t_r10_c36_1 + p_9_37;
  assign t_r10_c36_7 = t_r10_c36_2 + t_r10_c36_3;
  assign t_r10_c36_8 = t_r10_c36_4 + p_11_35;
  assign t_r10_c36_9 = t_r10_c36_5 + t_r10_c36_6;
  assign t_r10_c36_10 = t_r10_c36_7 + t_r10_c36_8;
  assign t_r10_c36_11 = t_r10_c36_9 + t_r10_c36_10;
  assign t_r10_c36_12 = t_r10_c36_11 + p_11_37;
  assign out_10_36 = t_r10_c36_12 >> 4;

  assign t_r10_c37_0 = p_9_37 << 1;
  assign t_r10_c37_1 = p_10_36 << 1;
  assign t_r10_c37_2 = p_10_37 << 2;
  assign t_r10_c37_3 = p_10_38 << 1;
  assign t_r10_c37_4 = p_11_37 << 1;
  assign t_r10_c37_5 = t_r10_c37_0 + p_9_36;
  assign t_r10_c37_6 = t_r10_c37_1 + p_9_38;
  assign t_r10_c37_7 = t_r10_c37_2 + t_r10_c37_3;
  assign t_r10_c37_8 = t_r10_c37_4 + p_11_36;
  assign t_r10_c37_9 = t_r10_c37_5 + t_r10_c37_6;
  assign t_r10_c37_10 = t_r10_c37_7 + t_r10_c37_8;
  assign t_r10_c37_11 = t_r10_c37_9 + t_r10_c37_10;
  assign t_r10_c37_12 = t_r10_c37_11 + p_11_38;
  assign out_10_37 = t_r10_c37_12 >> 4;

  assign t_r10_c38_0 = p_9_38 << 1;
  assign t_r10_c38_1 = p_10_37 << 1;
  assign t_r10_c38_2 = p_10_38 << 2;
  assign t_r10_c38_3 = p_10_39 << 1;
  assign t_r10_c38_4 = p_11_38 << 1;
  assign t_r10_c38_5 = t_r10_c38_0 + p_9_37;
  assign t_r10_c38_6 = t_r10_c38_1 + p_9_39;
  assign t_r10_c38_7 = t_r10_c38_2 + t_r10_c38_3;
  assign t_r10_c38_8 = t_r10_c38_4 + p_11_37;
  assign t_r10_c38_9 = t_r10_c38_5 + t_r10_c38_6;
  assign t_r10_c38_10 = t_r10_c38_7 + t_r10_c38_8;
  assign t_r10_c38_11 = t_r10_c38_9 + t_r10_c38_10;
  assign t_r10_c38_12 = t_r10_c38_11 + p_11_39;
  assign out_10_38 = t_r10_c38_12 >> 4;

  assign t_r10_c39_0 = p_9_39 << 1;
  assign t_r10_c39_1 = p_10_38 << 1;
  assign t_r10_c39_2 = p_10_39 << 2;
  assign t_r10_c39_3 = p_10_40 << 1;
  assign t_r10_c39_4 = p_11_39 << 1;
  assign t_r10_c39_5 = t_r10_c39_0 + p_9_38;
  assign t_r10_c39_6 = t_r10_c39_1 + p_9_40;
  assign t_r10_c39_7 = t_r10_c39_2 + t_r10_c39_3;
  assign t_r10_c39_8 = t_r10_c39_4 + p_11_38;
  assign t_r10_c39_9 = t_r10_c39_5 + t_r10_c39_6;
  assign t_r10_c39_10 = t_r10_c39_7 + t_r10_c39_8;
  assign t_r10_c39_11 = t_r10_c39_9 + t_r10_c39_10;
  assign t_r10_c39_12 = t_r10_c39_11 + p_11_40;
  assign out_10_39 = t_r10_c39_12 >> 4;

  assign t_r10_c40_0 = p_9_40 << 1;
  assign t_r10_c40_1 = p_10_39 << 1;
  assign t_r10_c40_2 = p_10_40 << 2;
  assign t_r10_c40_3 = p_10_41 << 1;
  assign t_r10_c40_4 = p_11_40 << 1;
  assign t_r10_c40_5 = t_r10_c40_0 + p_9_39;
  assign t_r10_c40_6 = t_r10_c40_1 + p_9_41;
  assign t_r10_c40_7 = t_r10_c40_2 + t_r10_c40_3;
  assign t_r10_c40_8 = t_r10_c40_4 + p_11_39;
  assign t_r10_c40_9 = t_r10_c40_5 + t_r10_c40_6;
  assign t_r10_c40_10 = t_r10_c40_7 + t_r10_c40_8;
  assign t_r10_c40_11 = t_r10_c40_9 + t_r10_c40_10;
  assign t_r10_c40_12 = t_r10_c40_11 + p_11_41;
  assign out_10_40 = t_r10_c40_12 >> 4;

  assign t_r10_c41_0 = p_9_41 << 1;
  assign t_r10_c41_1 = p_10_40 << 1;
  assign t_r10_c41_2 = p_10_41 << 2;
  assign t_r10_c41_3 = p_10_42 << 1;
  assign t_r10_c41_4 = p_11_41 << 1;
  assign t_r10_c41_5 = t_r10_c41_0 + p_9_40;
  assign t_r10_c41_6 = t_r10_c41_1 + p_9_42;
  assign t_r10_c41_7 = t_r10_c41_2 + t_r10_c41_3;
  assign t_r10_c41_8 = t_r10_c41_4 + p_11_40;
  assign t_r10_c41_9 = t_r10_c41_5 + t_r10_c41_6;
  assign t_r10_c41_10 = t_r10_c41_7 + t_r10_c41_8;
  assign t_r10_c41_11 = t_r10_c41_9 + t_r10_c41_10;
  assign t_r10_c41_12 = t_r10_c41_11 + p_11_42;
  assign out_10_41 = t_r10_c41_12 >> 4;

  assign t_r10_c42_0 = p_9_42 << 1;
  assign t_r10_c42_1 = p_10_41 << 1;
  assign t_r10_c42_2 = p_10_42 << 2;
  assign t_r10_c42_3 = p_10_43 << 1;
  assign t_r10_c42_4 = p_11_42 << 1;
  assign t_r10_c42_5 = t_r10_c42_0 + p_9_41;
  assign t_r10_c42_6 = t_r10_c42_1 + p_9_43;
  assign t_r10_c42_7 = t_r10_c42_2 + t_r10_c42_3;
  assign t_r10_c42_8 = t_r10_c42_4 + p_11_41;
  assign t_r10_c42_9 = t_r10_c42_5 + t_r10_c42_6;
  assign t_r10_c42_10 = t_r10_c42_7 + t_r10_c42_8;
  assign t_r10_c42_11 = t_r10_c42_9 + t_r10_c42_10;
  assign t_r10_c42_12 = t_r10_c42_11 + p_11_43;
  assign out_10_42 = t_r10_c42_12 >> 4;

  assign t_r10_c43_0 = p_9_43 << 1;
  assign t_r10_c43_1 = p_10_42 << 1;
  assign t_r10_c43_2 = p_10_43 << 2;
  assign t_r10_c43_3 = p_10_44 << 1;
  assign t_r10_c43_4 = p_11_43 << 1;
  assign t_r10_c43_5 = t_r10_c43_0 + p_9_42;
  assign t_r10_c43_6 = t_r10_c43_1 + p_9_44;
  assign t_r10_c43_7 = t_r10_c43_2 + t_r10_c43_3;
  assign t_r10_c43_8 = t_r10_c43_4 + p_11_42;
  assign t_r10_c43_9 = t_r10_c43_5 + t_r10_c43_6;
  assign t_r10_c43_10 = t_r10_c43_7 + t_r10_c43_8;
  assign t_r10_c43_11 = t_r10_c43_9 + t_r10_c43_10;
  assign t_r10_c43_12 = t_r10_c43_11 + p_11_44;
  assign out_10_43 = t_r10_c43_12 >> 4;

  assign t_r10_c44_0 = p_9_44 << 1;
  assign t_r10_c44_1 = p_10_43 << 1;
  assign t_r10_c44_2 = p_10_44 << 2;
  assign t_r10_c44_3 = p_10_45 << 1;
  assign t_r10_c44_4 = p_11_44 << 1;
  assign t_r10_c44_5 = t_r10_c44_0 + p_9_43;
  assign t_r10_c44_6 = t_r10_c44_1 + p_9_45;
  assign t_r10_c44_7 = t_r10_c44_2 + t_r10_c44_3;
  assign t_r10_c44_8 = t_r10_c44_4 + p_11_43;
  assign t_r10_c44_9 = t_r10_c44_5 + t_r10_c44_6;
  assign t_r10_c44_10 = t_r10_c44_7 + t_r10_c44_8;
  assign t_r10_c44_11 = t_r10_c44_9 + t_r10_c44_10;
  assign t_r10_c44_12 = t_r10_c44_11 + p_11_45;
  assign out_10_44 = t_r10_c44_12 >> 4;

  assign t_r10_c45_0 = p_9_45 << 1;
  assign t_r10_c45_1 = p_10_44 << 1;
  assign t_r10_c45_2 = p_10_45 << 2;
  assign t_r10_c45_3 = p_10_46 << 1;
  assign t_r10_c45_4 = p_11_45 << 1;
  assign t_r10_c45_5 = t_r10_c45_0 + p_9_44;
  assign t_r10_c45_6 = t_r10_c45_1 + p_9_46;
  assign t_r10_c45_7 = t_r10_c45_2 + t_r10_c45_3;
  assign t_r10_c45_8 = t_r10_c45_4 + p_11_44;
  assign t_r10_c45_9 = t_r10_c45_5 + t_r10_c45_6;
  assign t_r10_c45_10 = t_r10_c45_7 + t_r10_c45_8;
  assign t_r10_c45_11 = t_r10_c45_9 + t_r10_c45_10;
  assign t_r10_c45_12 = t_r10_c45_11 + p_11_46;
  assign out_10_45 = t_r10_c45_12 >> 4;

  assign t_r10_c46_0 = p_9_46 << 1;
  assign t_r10_c46_1 = p_10_45 << 1;
  assign t_r10_c46_2 = p_10_46 << 2;
  assign t_r10_c46_3 = p_10_47 << 1;
  assign t_r10_c46_4 = p_11_46 << 1;
  assign t_r10_c46_5 = t_r10_c46_0 + p_9_45;
  assign t_r10_c46_6 = t_r10_c46_1 + p_9_47;
  assign t_r10_c46_7 = t_r10_c46_2 + t_r10_c46_3;
  assign t_r10_c46_8 = t_r10_c46_4 + p_11_45;
  assign t_r10_c46_9 = t_r10_c46_5 + t_r10_c46_6;
  assign t_r10_c46_10 = t_r10_c46_7 + t_r10_c46_8;
  assign t_r10_c46_11 = t_r10_c46_9 + t_r10_c46_10;
  assign t_r10_c46_12 = t_r10_c46_11 + p_11_47;
  assign out_10_46 = t_r10_c46_12 >> 4;

  assign t_r10_c47_0 = p_9_47 << 1;
  assign t_r10_c47_1 = p_10_46 << 1;
  assign t_r10_c47_2 = p_10_47 << 2;
  assign t_r10_c47_3 = p_10_48 << 1;
  assign t_r10_c47_4 = p_11_47 << 1;
  assign t_r10_c47_5 = t_r10_c47_0 + p_9_46;
  assign t_r10_c47_6 = t_r10_c47_1 + p_9_48;
  assign t_r10_c47_7 = t_r10_c47_2 + t_r10_c47_3;
  assign t_r10_c47_8 = t_r10_c47_4 + p_11_46;
  assign t_r10_c47_9 = t_r10_c47_5 + t_r10_c47_6;
  assign t_r10_c47_10 = t_r10_c47_7 + t_r10_c47_8;
  assign t_r10_c47_11 = t_r10_c47_9 + t_r10_c47_10;
  assign t_r10_c47_12 = t_r10_c47_11 + p_11_48;
  assign out_10_47 = t_r10_c47_12 >> 4;

  assign t_r10_c48_0 = p_9_48 << 1;
  assign t_r10_c48_1 = p_10_47 << 1;
  assign t_r10_c48_2 = p_10_48 << 2;
  assign t_r10_c48_3 = p_10_49 << 1;
  assign t_r10_c48_4 = p_11_48 << 1;
  assign t_r10_c48_5 = t_r10_c48_0 + p_9_47;
  assign t_r10_c48_6 = t_r10_c48_1 + p_9_49;
  assign t_r10_c48_7 = t_r10_c48_2 + t_r10_c48_3;
  assign t_r10_c48_8 = t_r10_c48_4 + p_11_47;
  assign t_r10_c48_9 = t_r10_c48_5 + t_r10_c48_6;
  assign t_r10_c48_10 = t_r10_c48_7 + t_r10_c48_8;
  assign t_r10_c48_11 = t_r10_c48_9 + t_r10_c48_10;
  assign t_r10_c48_12 = t_r10_c48_11 + p_11_49;
  assign out_10_48 = t_r10_c48_12 >> 4;

  assign t_r10_c49_0 = p_9_49 << 1;
  assign t_r10_c49_1 = p_10_48 << 1;
  assign t_r10_c49_2 = p_10_49 << 2;
  assign t_r10_c49_3 = p_10_50 << 1;
  assign t_r10_c49_4 = p_11_49 << 1;
  assign t_r10_c49_5 = t_r10_c49_0 + p_9_48;
  assign t_r10_c49_6 = t_r10_c49_1 + p_9_50;
  assign t_r10_c49_7 = t_r10_c49_2 + t_r10_c49_3;
  assign t_r10_c49_8 = t_r10_c49_4 + p_11_48;
  assign t_r10_c49_9 = t_r10_c49_5 + t_r10_c49_6;
  assign t_r10_c49_10 = t_r10_c49_7 + t_r10_c49_8;
  assign t_r10_c49_11 = t_r10_c49_9 + t_r10_c49_10;
  assign t_r10_c49_12 = t_r10_c49_11 + p_11_50;
  assign out_10_49 = t_r10_c49_12 >> 4;

  assign t_r10_c50_0 = p_9_50 << 1;
  assign t_r10_c50_1 = p_10_49 << 1;
  assign t_r10_c50_2 = p_10_50 << 2;
  assign t_r10_c50_3 = p_10_51 << 1;
  assign t_r10_c50_4 = p_11_50 << 1;
  assign t_r10_c50_5 = t_r10_c50_0 + p_9_49;
  assign t_r10_c50_6 = t_r10_c50_1 + p_9_51;
  assign t_r10_c50_7 = t_r10_c50_2 + t_r10_c50_3;
  assign t_r10_c50_8 = t_r10_c50_4 + p_11_49;
  assign t_r10_c50_9 = t_r10_c50_5 + t_r10_c50_6;
  assign t_r10_c50_10 = t_r10_c50_7 + t_r10_c50_8;
  assign t_r10_c50_11 = t_r10_c50_9 + t_r10_c50_10;
  assign t_r10_c50_12 = t_r10_c50_11 + p_11_51;
  assign out_10_50 = t_r10_c50_12 >> 4;

  assign t_r10_c51_0 = p_9_51 << 1;
  assign t_r10_c51_1 = p_10_50 << 1;
  assign t_r10_c51_2 = p_10_51 << 2;
  assign t_r10_c51_3 = p_10_52 << 1;
  assign t_r10_c51_4 = p_11_51 << 1;
  assign t_r10_c51_5 = t_r10_c51_0 + p_9_50;
  assign t_r10_c51_6 = t_r10_c51_1 + p_9_52;
  assign t_r10_c51_7 = t_r10_c51_2 + t_r10_c51_3;
  assign t_r10_c51_8 = t_r10_c51_4 + p_11_50;
  assign t_r10_c51_9 = t_r10_c51_5 + t_r10_c51_6;
  assign t_r10_c51_10 = t_r10_c51_7 + t_r10_c51_8;
  assign t_r10_c51_11 = t_r10_c51_9 + t_r10_c51_10;
  assign t_r10_c51_12 = t_r10_c51_11 + p_11_52;
  assign out_10_51 = t_r10_c51_12 >> 4;

  assign t_r10_c52_0 = p_9_52 << 1;
  assign t_r10_c52_1 = p_10_51 << 1;
  assign t_r10_c52_2 = p_10_52 << 2;
  assign t_r10_c52_3 = p_10_53 << 1;
  assign t_r10_c52_4 = p_11_52 << 1;
  assign t_r10_c52_5 = t_r10_c52_0 + p_9_51;
  assign t_r10_c52_6 = t_r10_c52_1 + p_9_53;
  assign t_r10_c52_7 = t_r10_c52_2 + t_r10_c52_3;
  assign t_r10_c52_8 = t_r10_c52_4 + p_11_51;
  assign t_r10_c52_9 = t_r10_c52_5 + t_r10_c52_6;
  assign t_r10_c52_10 = t_r10_c52_7 + t_r10_c52_8;
  assign t_r10_c52_11 = t_r10_c52_9 + t_r10_c52_10;
  assign t_r10_c52_12 = t_r10_c52_11 + p_11_53;
  assign out_10_52 = t_r10_c52_12 >> 4;

  assign t_r10_c53_0 = p_9_53 << 1;
  assign t_r10_c53_1 = p_10_52 << 1;
  assign t_r10_c53_2 = p_10_53 << 2;
  assign t_r10_c53_3 = p_10_54 << 1;
  assign t_r10_c53_4 = p_11_53 << 1;
  assign t_r10_c53_5 = t_r10_c53_0 + p_9_52;
  assign t_r10_c53_6 = t_r10_c53_1 + p_9_54;
  assign t_r10_c53_7 = t_r10_c53_2 + t_r10_c53_3;
  assign t_r10_c53_8 = t_r10_c53_4 + p_11_52;
  assign t_r10_c53_9 = t_r10_c53_5 + t_r10_c53_6;
  assign t_r10_c53_10 = t_r10_c53_7 + t_r10_c53_8;
  assign t_r10_c53_11 = t_r10_c53_9 + t_r10_c53_10;
  assign t_r10_c53_12 = t_r10_c53_11 + p_11_54;
  assign out_10_53 = t_r10_c53_12 >> 4;

  assign t_r10_c54_0 = p_9_54 << 1;
  assign t_r10_c54_1 = p_10_53 << 1;
  assign t_r10_c54_2 = p_10_54 << 2;
  assign t_r10_c54_3 = p_10_55 << 1;
  assign t_r10_c54_4 = p_11_54 << 1;
  assign t_r10_c54_5 = t_r10_c54_0 + p_9_53;
  assign t_r10_c54_6 = t_r10_c54_1 + p_9_55;
  assign t_r10_c54_7 = t_r10_c54_2 + t_r10_c54_3;
  assign t_r10_c54_8 = t_r10_c54_4 + p_11_53;
  assign t_r10_c54_9 = t_r10_c54_5 + t_r10_c54_6;
  assign t_r10_c54_10 = t_r10_c54_7 + t_r10_c54_8;
  assign t_r10_c54_11 = t_r10_c54_9 + t_r10_c54_10;
  assign t_r10_c54_12 = t_r10_c54_11 + p_11_55;
  assign out_10_54 = t_r10_c54_12 >> 4;

  assign t_r10_c55_0 = p_9_55 << 1;
  assign t_r10_c55_1 = p_10_54 << 1;
  assign t_r10_c55_2 = p_10_55 << 2;
  assign t_r10_c55_3 = p_10_56 << 1;
  assign t_r10_c55_4 = p_11_55 << 1;
  assign t_r10_c55_5 = t_r10_c55_0 + p_9_54;
  assign t_r10_c55_6 = t_r10_c55_1 + p_9_56;
  assign t_r10_c55_7 = t_r10_c55_2 + t_r10_c55_3;
  assign t_r10_c55_8 = t_r10_c55_4 + p_11_54;
  assign t_r10_c55_9 = t_r10_c55_5 + t_r10_c55_6;
  assign t_r10_c55_10 = t_r10_c55_7 + t_r10_c55_8;
  assign t_r10_c55_11 = t_r10_c55_9 + t_r10_c55_10;
  assign t_r10_c55_12 = t_r10_c55_11 + p_11_56;
  assign out_10_55 = t_r10_c55_12 >> 4;

  assign t_r10_c56_0 = p_9_56 << 1;
  assign t_r10_c56_1 = p_10_55 << 1;
  assign t_r10_c56_2 = p_10_56 << 2;
  assign t_r10_c56_3 = p_10_57 << 1;
  assign t_r10_c56_4 = p_11_56 << 1;
  assign t_r10_c56_5 = t_r10_c56_0 + p_9_55;
  assign t_r10_c56_6 = t_r10_c56_1 + p_9_57;
  assign t_r10_c56_7 = t_r10_c56_2 + t_r10_c56_3;
  assign t_r10_c56_8 = t_r10_c56_4 + p_11_55;
  assign t_r10_c56_9 = t_r10_c56_5 + t_r10_c56_6;
  assign t_r10_c56_10 = t_r10_c56_7 + t_r10_c56_8;
  assign t_r10_c56_11 = t_r10_c56_9 + t_r10_c56_10;
  assign t_r10_c56_12 = t_r10_c56_11 + p_11_57;
  assign out_10_56 = t_r10_c56_12 >> 4;

  assign t_r10_c57_0 = p_9_57 << 1;
  assign t_r10_c57_1 = p_10_56 << 1;
  assign t_r10_c57_2 = p_10_57 << 2;
  assign t_r10_c57_3 = p_10_58 << 1;
  assign t_r10_c57_4 = p_11_57 << 1;
  assign t_r10_c57_5 = t_r10_c57_0 + p_9_56;
  assign t_r10_c57_6 = t_r10_c57_1 + p_9_58;
  assign t_r10_c57_7 = t_r10_c57_2 + t_r10_c57_3;
  assign t_r10_c57_8 = t_r10_c57_4 + p_11_56;
  assign t_r10_c57_9 = t_r10_c57_5 + t_r10_c57_6;
  assign t_r10_c57_10 = t_r10_c57_7 + t_r10_c57_8;
  assign t_r10_c57_11 = t_r10_c57_9 + t_r10_c57_10;
  assign t_r10_c57_12 = t_r10_c57_11 + p_11_58;
  assign out_10_57 = t_r10_c57_12 >> 4;

  assign t_r10_c58_0 = p_9_58 << 1;
  assign t_r10_c58_1 = p_10_57 << 1;
  assign t_r10_c58_2 = p_10_58 << 2;
  assign t_r10_c58_3 = p_10_59 << 1;
  assign t_r10_c58_4 = p_11_58 << 1;
  assign t_r10_c58_5 = t_r10_c58_0 + p_9_57;
  assign t_r10_c58_6 = t_r10_c58_1 + p_9_59;
  assign t_r10_c58_7 = t_r10_c58_2 + t_r10_c58_3;
  assign t_r10_c58_8 = t_r10_c58_4 + p_11_57;
  assign t_r10_c58_9 = t_r10_c58_5 + t_r10_c58_6;
  assign t_r10_c58_10 = t_r10_c58_7 + t_r10_c58_8;
  assign t_r10_c58_11 = t_r10_c58_9 + t_r10_c58_10;
  assign t_r10_c58_12 = t_r10_c58_11 + p_11_59;
  assign out_10_58 = t_r10_c58_12 >> 4;

  assign t_r10_c59_0 = p_9_59 << 1;
  assign t_r10_c59_1 = p_10_58 << 1;
  assign t_r10_c59_2 = p_10_59 << 2;
  assign t_r10_c59_3 = p_10_60 << 1;
  assign t_r10_c59_4 = p_11_59 << 1;
  assign t_r10_c59_5 = t_r10_c59_0 + p_9_58;
  assign t_r10_c59_6 = t_r10_c59_1 + p_9_60;
  assign t_r10_c59_7 = t_r10_c59_2 + t_r10_c59_3;
  assign t_r10_c59_8 = t_r10_c59_4 + p_11_58;
  assign t_r10_c59_9 = t_r10_c59_5 + t_r10_c59_6;
  assign t_r10_c59_10 = t_r10_c59_7 + t_r10_c59_8;
  assign t_r10_c59_11 = t_r10_c59_9 + t_r10_c59_10;
  assign t_r10_c59_12 = t_r10_c59_11 + p_11_60;
  assign out_10_59 = t_r10_c59_12 >> 4;

  assign t_r10_c60_0 = p_9_60 << 1;
  assign t_r10_c60_1 = p_10_59 << 1;
  assign t_r10_c60_2 = p_10_60 << 2;
  assign t_r10_c60_3 = p_10_61 << 1;
  assign t_r10_c60_4 = p_11_60 << 1;
  assign t_r10_c60_5 = t_r10_c60_0 + p_9_59;
  assign t_r10_c60_6 = t_r10_c60_1 + p_9_61;
  assign t_r10_c60_7 = t_r10_c60_2 + t_r10_c60_3;
  assign t_r10_c60_8 = t_r10_c60_4 + p_11_59;
  assign t_r10_c60_9 = t_r10_c60_5 + t_r10_c60_6;
  assign t_r10_c60_10 = t_r10_c60_7 + t_r10_c60_8;
  assign t_r10_c60_11 = t_r10_c60_9 + t_r10_c60_10;
  assign t_r10_c60_12 = t_r10_c60_11 + p_11_61;
  assign out_10_60 = t_r10_c60_12 >> 4;

  assign t_r10_c61_0 = p_9_61 << 1;
  assign t_r10_c61_1 = p_10_60 << 1;
  assign t_r10_c61_2 = p_10_61 << 2;
  assign t_r10_c61_3 = p_10_62 << 1;
  assign t_r10_c61_4 = p_11_61 << 1;
  assign t_r10_c61_5 = t_r10_c61_0 + p_9_60;
  assign t_r10_c61_6 = t_r10_c61_1 + p_9_62;
  assign t_r10_c61_7 = t_r10_c61_2 + t_r10_c61_3;
  assign t_r10_c61_8 = t_r10_c61_4 + p_11_60;
  assign t_r10_c61_9 = t_r10_c61_5 + t_r10_c61_6;
  assign t_r10_c61_10 = t_r10_c61_7 + t_r10_c61_8;
  assign t_r10_c61_11 = t_r10_c61_9 + t_r10_c61_10;
  assign t_r10_c61_12 = t_r10_c61_11 + p_11_62;
  assign out_10_61 = t_r10_c61_12 >> 4;

  assign t_r10_c62_0 = p_9_62 << 1;
  assign t_r10_c62_1 = p_10_61 << 1;
  assign t_r10_c62_2 = p_10_62 << 2;
  assign t_r10_c62_3 = p_10_63 << 1;
  assign t_r10_c62_4 = p_11_62 << 1;
  assign t_r10_c62_5 = t_r10_c62_0 + p_9_61;
  assign t_r10_c62_6 = t_r10_c62_1 + p_9_63;
  assign t_r10_c62_7 = t_r10_c62_2 + t_r10_c62_3;
  assign t_r10_c62_8 = t_r10_c62_4 + p_11_61;
  assign t_r10_c62_9 = t_r10_c62_5 + t_r10_c62_6;
  assign t_r10_c62_10 = t_r10_c62_7 + t_r10_c62_8;
  assign t_r10_c62_11 = t_r10_c62_9 + t_r10_c62_10;
  assign t_r10_c62_12 = t_r10_c62_11 + p_11_63;
  assign out_10_62 = t_r10_c62_12 >> 4;

  assign t_r10_c63_0 = p_9_63 << 1;
  assign t_r10_c63_1 = p_10_62 << 1;
  assign t_r10_c63_2 = p_10_63 << 2;
  assign t_r10_c63_3 = p_10_64 << 1;
  assign t_r10_c63_4 = p_11_63 << 1;
  assign t_r10_c63_5 = t_r10_c63_0 + p_9_62;
  assign t_r10_c63_6 = t_r10_c63_1 + p_9_64;
  assign t_r10_c63_7 = t_r10_c63_2 + t_r10_c63_3;
  assign t_r10_c63_8 = t_r10_c63_4 + p_11_62;
  assign t_r10_c63_9 = t_r10_c63_5 + t_r10_c63_6;
  assign t_r10_c63_10 = t_r10_c63_7 + t_r10_c63_8;
  assign t_r10_c63_11 = t_r10_c63_9 + t_r10_c63_10;
  assign t_r10_c63_12 = t_r10_c63_11 + p_11_64;
  assign out_10_63 = t_r10_c63_12 >> 4;

  assign t_r10_c64_0 = p_9_64 << 1;
  assign t_r10_c64_1 = p_10_63 << 1;
  assign t_r10_c64_2 = p_10_64 << 2;
  assign t_r10_c64_3 = p_10_65 << 1;
  assign t_r10_c64_4 = p_11_64 << 1;
  assign t_r10_c64_5 = t_r10_c64_0 + p_9_63;
  assign t_r10_c64_6 = t_r10_c64_1 + p_9_65;
  assign t_r10_c64_7 = t_r10_c64_2 + t_r10_c64_3;
  assign t_r10_c64_8 = t_r10_c64_4 + p_11_63;
  assign t_r10_c64_9 = t_r10_c64_5 + t_r10_c64_6;
  assign t_r10_c64_10 = t_r10_c64_7 + t_r10_c64_8;
  assign t_r10_c64_11 = t_r10_c64_9 + t_r10_c64_10;
  assign t_r10_c64_12 = t_r10_c64_11 + p_11_65;
  assign out_10_64 = t_r10_c64_12 >> 4;

  assign t_r11_c1_0 = p_10_1 << 1;
  assign t_r11_c1_1 = p_11_0 << 1;
  assign t_r11_c1_2 = p_11_1 << 2;
  assign t_r11_c1_3 = p_11_2 << 1;
  assign t_r11_c1_4 = p_12_1 << 1;
  assign t_r11_c1_5 = t_r11_c1_0 + p_10_0;
  assign t_r11_c1_6 = t_r11_c1_1 + p_10_2;
  assign t_r11_c1_7 = t_r11_c1_2 + t_r11_c1_3;
  assign t_r11_c1_8 = t_r11_c1_4 + p_12_0;
  assign t_r11_c1_9 = t_r11_c1_5 + t_r11_c1_6;
  assign t_r11_c1_10 = t_r11_c1_7 + t_r11_c1_8;
  assign t_r11_c1_11 = t_r11_c1_9 + t_r11_c1_10;
  assign t_r11_c1_12 = t_r11_c1_11 + p_12_2;
  assign out_11_1 = t_r11_c1_12 >> 4;

  assign t_r11_c2_0 = p_10_2 << 1;
  assign t_r11_c2_1 = p_11_1 << 1;
  assign t_r11_c2_2 = p_11_2 << 2;
  assign t_r11_c2_3 = p_11_3 << 1;
  assign t_r11_c2_4 = p_12_2 << 1;
  assign t_r11_c2_5 = t_r11_c2_0 + p_10_1;
  assign t_r11_c2_6 = t_r11_c2_1 + p_10_3;
  assign t_r11_c2_7 = t_r11_c2_2 + t_r11_c2_3;
  assign t_r11_c2_8 = t_r11_c2_4 + p_12_1;
  assign t_r11_c2_9 = t_r11_c2_5 + t_r11_c2_6;
  assign t_r11_c2_10 = t_r11_c2_7 + t_r11_c2_8;
  assign t_r11_c2_11 = t_r11_c2_9 + t_r11_c2_10;
  assign t_r11_c2_12 = t_r11_c2_11 + p_12_3;
  assign out_11_2 = t_r11_c2_12 >> 4;

  assign t_r11_c3_0 = p_10_3 << 1;
  assign t_r11_c3_1 = p_11_2 << 1;
  assign t_r11_c3_2 = p_11_3 << 2;
  assign t_r11_c3_3 = p_11_4 << 1;
  assign t_r11_c3_4 = p_12_3 << 1;
  assign t_r11_c3_5 = t_r11_c3_0 + p_10_2;
  assign t_r11_c3_6 = t_r11_c3_1 + p_10_4;
  assign t_r11_c3_7 = t_r11_c3_2 + t_r11_c3_3;
  assign t_r11_c3_8 = t_r11_c3_4 + p_12_2;
  assign t_r11_c3_9 = t_r11_c3_5 + t_r11_c3_6;
  assign t_r11_c3_10 = t_r11_c3_7 + t_r11_c3_8;
  assign t_r11_c3_11 = t_r11_c3_9 + t_r11_c3_10;
  assign t_r11_c3_12 = t_r11_c3_11 + p_12_4;
  assign out_11_3 = t_r11_c3_12 >> 4;

  assign t_r11_c4_0 = p_10_4 << 1;
  assign t_r11_c4_1 = p_11_3 << 1;
  assign t_r11_c4_2 = p_11_4 << 2;
  assign t_r11_c4_3 = p_11_5 << 1;
  assign t_r11_c4_4 = p_12_4 << 1;
  assign t_r11_c4_5 = t_r11_c4_0 + p_10_3;
  assign t_r11_c4_6 = t_r11_c4_1 + p_10_5;
  assign t_r11_c4_7 = t_r11_c4_2 + t_r11_c4_3;
  assign t_r11_c4_8 = t_r11_c4_4 + p_12_3;
  assign t_r11_c4_9 = t_r11_c4_5 + t_r11_c4_6;
  assign t_r11_c4_10 = t_r11_c4_7 + t_r11_c4_8;
  assign t_r11_c4_11 = t_r11_c4_9 + t_r11_c4_10;
  assign t_r11_c4_12 = t_r11_c4_11 + p_12_5;
  assign out_11_4 = t_r11_c4_12 >> 4;

  assign t_r11_c5_0 = p_10_5 << 1;
  assign t_r11_c5_1 = p_11_4 << 1;
  assign t_r11_c5_2 = p_11_5 << 2;
  assign t_r11_c5_3 = p_11_6 << 1;
  assign t_r11_c5_4 = p_12_5 << 1;
  assign t_r11_c5_5 = t_r11_c5_0 + p_10_4;
  assign t_r11_c5_6 = t_r11_c5_1 + p_10_6;
  assign t_r11_c5_7 = t_r11_c5_2 + t_r11_c5_3;
  assign t_r11_c5_8 = t_r11_c5_4 + p_12_4;
  assign t_r11_c5_9 = t_r11_c5_5 + t_r11_c5_6;
  assign t_r11_c5_10 = t_r11_c5_7 + t_r11_c5_8;
  assign t_r11_c5_11 = t_r11_c5_9 + t_r11_c5_10;
  assign t_r11_c5_12 = t_r11_c5_11 + p_12_6;
  assign out_11_5 = t_r11_c5_12 >> 4;

  assign t_r11_c6_0 = p_10_6 << 1;
  assign t_r11_c6_1 = p_11_5 << 1;
  assign t_r11_c6_2 = p_11_6 << 2;
  assign t_r11_c6_3 = p_11_7 << 1;
  assign t_r11_c6_4 = p_12_6 << 1;
  assign t_r11_c6_5 = t_r11_c6_0 + p_10_5;
  assign t_r11_c6_6 = t_r11_c6_1 + p_10_7;
  assign t_r11_c6_7 = t_r11_c6_2 + t_r11_c6_3;
  assign t_r11_c6_8 = t_r11_c6_4 + p_12_5;
  assign t_r11_c6_9 = t_r11_c6_5 + t_r11_c6_6;
  assign t_r11_c6_10 = t_r11_c6_7 + t_r11_c6_8;
  assign t_r11_c6_11 = t_r11_c6_9 + t_r11_c6_10;
  assign t_r11_c6_12 = t_r11_c6_11 + p_12_7;
  assign out_11_6 = t_r11_c6_12 >> 4;

  assign t_r11_c7_0 = p_10_7 << 1;
  assign t_r11_c7_1 = p_11_6 << 1;
  assign t_r11_c7_2 = p_11_7 << 2;
  assign t_r11_c7_3 = p_11_8 << 1;
  assign t_r11_c7_4 = p_12_7 << 1;
  assign t_r11_c7_5 = t_r11_c7_0 + p_10_6;
  assign t_r11_c7_6 = t_r11_c7_1 + p_10_8;
  assign t_r11_c7_7 = t_r11_c7_2 + t_r11_c7_3;
  assign t_r11_c7_8 = t_r11_c7_4 + p_12_6;
  assign t_r11_c7_9 = t_r11_c7_5 + t_r11_c7_6;
  assign t_r11_c7_10 = t_r11_c7_7 + t_r11_c7_8;
  assign t_r11_c7_11 = t_r11_c7_9 + t_r11_c7_10;
  assign t_r11_c7_12 = t_r11_c7_11 + p_12_8;
  assign out_11_7 = t_r11_c7_12 >> 4;

  assign t_r11_c8_0 = p_10_8 << 1;
  assign t_r11_c8_1 = p_11_7 << 1;
  assign t_r11_c8_2 = p_11_8 << 2;
  assign t_r11_c8_3 = p_11_9 << 1;
  assign t_r11_c8_4 = p_12_8 << 1;
  assign t_r11_c8_5 = t_r11_c8_0 + p_10_7;
  assign t_r11_c8_6 = t_r11_c8_1 + p_10_9;
  assign t_r11_c8_7 = t_r11_c8_2 + t_r11_c8_3;
  assign t_r11_c8_8 = t_r11_c8_4 + p_12_7;
  assign t_r11_c8_9 = t_r11_c8_5 + t_r11_c8_6;
  assign t_r11_c8_10 = t_r11_c8_7 + t_r11_c8_8;
  assign t_r11_c8_11 = t_r11_c8_9 + t_r11_c8_10;
  assign t_r11_c8_12 = t_r11_c8_11 + p_12_9;
  assign out_11_8 = t_r11_c8_12 >> 4;

  assign t_r11_c9_0 = p_10_9 << 1;
  assign t_r11_c9_1 = p_11_8 << 1;
  assign t_r11_c9_2 = p_11_9 << 2;
  assign t_r11_c9_3 = p_11_10 << 1;
  assign t_r11_c9_4 = p_12_9 << 1;
  assign t_r11_c9_5 = t_r11_c9_0 + p_10_8;
  assign t_r11_c9_6 = t_r11_c9_1 + p_10_10;
  assign t_r11_c9_7 = t_r11_c9_2 + t_r11_c9_3;
  assign t_r11_c9_8 = t_r11_c9_4 + p_12_8;
  assign t_r11_c9_9 = t_r11_c9_5 + t_r11_c9_6;
  assign t_r11_c9_10 = t_r11_c9_7 + t_r11_c9_8;
  assign t_r11_c9_11 = t_r11_c9_9 + t_r11_c9_10;
  assign t_r11_c9_12 = t_r11_c9_11 + p_12_10;
  assign out_11_9 = t_r11_c9_12 >> 4;

  assign t_r11_c10_0 = p_10_10 << 1;
  assign t_r11_c10_1 = p_11_9 << 1;
  assign t_r11_c10_2 = p_11_10 << 2;
  assign t_r11_c10_3 = p_11_11 << 1;
  assign t_r11_c10_4 = p_12_10 << 1;
  assign t_r11_c10_5 = t_r11_c10_0 + p_10_9;
  assign t_r11_c10_6 = t_r11_c10_1 + p_10_11;
  assign t_r11_c10_7 = t_r11_c10_2 + t_r11_c10_3;
  assign t_r11_c10_8 = t_r11_c10_4 + p_12_9;
  assign t_r11_c10_9 = t_r11_c10_5 + t_r11_c10_6;
  assign t_r11_c10_10 = t_r11_c10_7 + t_r11_c10_8;
  assign t_r11_c10_11 = t_r11_c10_9 + t_r11_c10_10;
  assign t_r11_c10_12 = t_r11_c10_11 + p_12_11;
  assign out_11_10 = t_r11_c10_12 >> 4;

  assign t_r11_c11_0 = p_10_11 << 1;
  assign t_r11_c11_1 = p_11_10 << 1;
  assign t_r11_c11_2 = p_11_11 << 2;
  assign t_r11_c11_3 = p_11_12 << 1;
  assign t_r11_c11_4 = p_12_11 << 1;
  assign t_r11_c11_5 = t_r11_c11_0 + p_10_10;
  assign t_r11_c11_6 = t_r11_c11_1 + p_10_12;
  assign t_r11_c11_7 = t_r11_c11_2 + t_r11_c11_3;
  assign t_r11_c11_8 = t_r11_c11_4 + p_12_10;
  assign t_r11_c11_9 = t_r11_c11_5 + t_r11_c11_6;
  assign t_r11_c11_10 = t_r11_c11_7 + t_r11_c11_8;
  assign t_r11_c11_11 = t_r11_c11_9 + t_r11_c11_10;
  assign t_r11_c11_12 = t_r11_c11_11 + p_12_12;
  assign out_11_11 = t_r11_c11_12 >> 4;

  assign t_r11_c12_0 = p_10_12 << 1;
  assign t_r11_c12_1 = p_11_11 << 1;
  assign t_r11_c12_2 = p_11_12 << 2;
  assign t_r11_c12_3 = p_11_13 << 1;
  assign t_r11_c12_4 = p_12_12 << 1;
  assign t_r11_c12_5 = t_r11_c12_0 + p_10_11;
  assign t_r11_c12_6 = t_r11_c12_1 + p_10_13;
  assign t_r11_c12_7 = t_r11_c12_2 + t_r11_c12_3;
  assign t_r11_c12_8 = t_r11_c12_4 + p_12_11;
  assign t_r11_c12_9 = t_r11_c12_5 + t_r11_c12_6;
  assign t_r11_c12_10 = t_r11_c12_7 + t_r11_c12_8;
  assign t_r11_c12_11 = t_r11_c12_9 + t_r11_c12_10;
  assign t_r11_c12_12 = t_r11_c12_11 + p_12_13;
  assign out_11_12 = t_r11_c12_12 >> 4;

  assign t_r11_c13_0 = p_10_13 << 1;
  assign t_r11_c13_1 = p_11_12 << 1;
  assign t_r11_c13_2 = p_11_13 << 2;
  assign t_r11_c13_3 = p_11_14 << 1;
  assign t_r11_c13_4 = p_12_13 << 1;
  assign t_r11_c13_5 = t_r11_c13_0 + p_10_12;
  assign t_r11_c13_6 = t_r11_c13_1 + p_10_14;
  assign t_r11_c13_7 = t_r11_c13_2 + t_r11_c13_3;
  assign t_r11_c13_8 = t_r11_c13_4 + p_12_12;
  assign t_r11_c13_9 = t_r11_c13_5 + t_r11_c13_6;
  assign t_r11_c13_10 = t_r11_c13_7 + t_r11_c13_8;
  assign t_r11_c13_11 = t_r11_c13_9 + t_r11_c13_10;
  assign t_r11_c13_12 = t_r11_c13_11 + p_12_14;
  assign out_11_13 = t_r11_c13_12 >> 4;

  assign t_r11_c14_0 = p_10_14 << 1;
  assign t_r11_c14_1 = p_11_13 << 1;
  assign t_r11_c14_2 = p_11_14 << 2;
  assign t_r11_c14_3 = p_11_15 << 1;
  assign t_r11_c14_4 = p_12_14 << 1;
  assign t_r11_c14_5 = t_r11_c14_0 + p_10_13;
  assign t_r11_c14_6 = t_r11_c14_1 + p_10_15;
  assign t_r11_c14_7 = t_r11_c14_2 + t_r11_c14_3;
  assign t_r11_c14_8 = t_r11_c14_4 + p_12_13;
  assign t_r11_c14_9 = t_r11_c14_5 + t_r11_c14_6;
  assign t_r11_c14_10 = t_r11_c14_7 + t_r11_c14_8;
  assign t_r11_c14_11 = t_r11_c14_9 + t_r11_c14_10;
  assign t_r11_c14_12 = t_r11_c14_11 + p_12_15;
  assign out_11_14 = t_r11_c14_12 >> 4;

  assign t_r11_c15_0 = p_10_15 << 1;
  assign t_r11_c15_1 = p_11_14 << 1;
  assign t_r11_c15_2 = p_11_15 << 2;
  assign t_r11_c15_3 = p_11_16 << 1;
  assign t_r11_c15_4 = p_12_15 << 1;
  assign t_r11_c15_5 = t_r11_c15_0 + p_10_14;
  assign t_r11_c15_6 = t_r11_c15_1 + p_10_16;
  assign t_r11_c15_7 = t_r11_c15_2 + t_r11_c15_3;
  assign t_r11_c15_8 = t_r11_c15_4 + p_12_14;
  assign t_r11_c15_9 = t_r11_c15_5 + t_r11_c15_6;
  assign t_r11_c15_10 = t_r11_c15_7 + t_r11_c15_8;
  assign t_r11_c15_11 = t_r11_c15_9 + t_r11_c15_10;
  assign t_r11_c15_12 = t_r11_c15_11 + p_12_16;
  assign out_11_15 = t_r11_c15_12 >> 4;

  assign t_r11_c16_0 = p_10_16 << 1;
  assign t_r11_c16_1 = p_11_15 << 1;
  assign t_r11_c16_2 = p_11_16 << 2;
  assign t_r11_c16_3 = p_11_17 << 1;
  assign t_r11_c16_4 = p_12_16 << 1;
  assign t_r11_c16_5 = t_r11_c16_0 + p_10_15;
  assign t_r11_c16_6 = t_r11_c16_1 + p_10_17;
  assign t_r11_c16_7 = t_r11_c16_2 + t_r11_c16_3;
  assign t_r11_c16_8 = t_r11_c16_4 + p_12_15;
  assign t_r11_c16_9 = t_r11_c16_5 + t_r11_c16_6;
  assign t_r11_c16_10 = t_r11_c16_7 + t_r11_c16_8;
  assign t_r11_c16_11 = t_r11_c16_9 + t_r11_c16_10;
  assign t_r11_c16_12 = t_r11_c16_11 + p_12_17;
  assign out_11_16 = t_r11_c16_12 >> 4;

  assign t_r11_c17_0 = p_10_17 << 1;
  assign t_r11_c17_1 = p_11_16 << 1;
  assign t_r11_c17_2 = p_11_17 << 2;
  assign t_r11_c17_3 = p_11_18 << 1;
  assign t_r11_c17_4 = p_12_17 << 1;
  assign t_r11_c17_5 = t_r11_c17_0 + p_10_16;
  assign t_r11_c17_6 = t_r11_c17_1 + p_10_18;
  assign t_r11_c17_7 = t_r11_c17_2 + t_r11_c17_3;
  assign t_r11_c17_8 = t_r11_c17_4 + p_12_16;
  assign t_r11_c17_9 = t_r11_c17_5 + t_r11_c17_6;
  assign t_r11_c17_10 = t_r11_c17_7 + t_r11_c17_8;
  assign t_r11_c17_11 = t_r11_c17_9 + t_r11_c17_10;
  assign t_r11_c17_12 = t_r11_c17_11 + p_12_18;
  assign out_11_17 = t_r11_c17_12 >> 4;

  assign t_r11_c18_0 = p_10_18 << 1;
  assign t_r11_c18_1 = p_11_17 << 1;
  assign t_r11_c18_2 = p_11_18 << 2;
  assign t_r11_c18_3 = p_11_19 << 1;
  assign t_r11_c18_4 = p_12_18 << 1;
  assign t_r11_c18_5 = t_r11_c18_0 + p_10_17;
  assign t_r11_c18_6 = t_r11_c18_1 + p_10_19;
  assign t_r11_c18_7 = t_r11_c18_2 + t_r11_c18_3;
  assign t_r11_c18_8 = t_r11_c18_4 + p_12_17;
  assign t_r11_c18_9 = t_r11_c18_5 + t_r11_c18_6;
  assign t_r11_c18_10 = t_r11_c18_7 + t_r11_c18_8;
  assign t_r11_c18_11 = t_r11_c18_9 + t_r11_c18_10;
  assign t_r11_c18_12 = t_r11_c18_11 + p_12_19;
  assign out_11_18 = t_r11_c18_12 >> 4;

  assign t_r11_c19_0 = p_10_19 << 1;
  assign t_r11_c19_1 = p_11_18 << 1;
  assign t_r11_c19_2 = p_11_19 << 2;
  assign t_r11_c19_3 = p_11_20 << 1;
  assign t_r11_c19_4 = p_12_19 << 1;
  assign t_r11_c19_5 = t_r11_c19_0 + p_10_18;
  assign t_r11_c19_6 = t_r11_c19_1 + p_10_20;
  assign t_r11_c19_7 = t_r11_c19_2 + t_r11_c19_3;
  assign t_r11_c19_8 = t_r11_c19_4 + p_12_18;
  assign t_r11_c19_9 = t_r11_c19_5 + t_r11_c19_6;
  assign t_r11_c19_10 = t_r11_c19_7 + t_r11_c19_8;
  assign t_r11_c19_11 = t_r11_c19_9 + t_r11_c19_10;
  assign t_r11_c19_12 = t_r11_c19_11 + p_12_20;
  assign out_11_19 = t_r11_c19_12 >> 4;

  assign t_r11_c20_0 = p_10_20 << 1;
  assign t_r11_c20_1 = p_11_19 << 1;
  assign t_r11_c20_2 = p_11_20 << 2;
  assign t_r11_c20_3 = p_11_21 << 1;
  assign t_r11_c20_4 = p_12_20 << 1;
  assign t_r11_c20_5 = t_r11_c20_0 + p_10_19;
  assign t_r11_c20_6 = t_r11_c20_1 + p_10_21;
  assign t_r11_c20_7 = t_r11_c20_2 + t_r11_c20_3;
  assign t_r11_c20_8 = t_r11_c20_4 + p_12_19;
  assign t_r11_c20_9 = t_r11_c20_5 + t_r11_c20_6;
  assign t_r11_c20_10 = t_r11_c20_7 + t_r11_c20_8;
  assign t_r11_c20_11 = t_r11_c20_9 + t_r11_c20_10;
  assign t_r11_c20_12 = t_r11_c20_11 + p_12_21;
  assign out_11_20 = t_r11_c20_12 >> 4;

  assign t_r11_c21_0 = p_10_21 << 1;
  assign t_r11_c21_1 = p_11_20 << 1;
  assign t_r11_c21_2 = p_11_21 << 2;
  assign t_r11_c21_3 = p_11_22 << 1;
  assign t_r11_c21_4 = p_12_21 << 1;
  assign t_r11_c21_5 = t_r11_c21_0 + p_10_20;
  assign t_r11_c21_6 = t_r11_c21_1 + p_10_22;
  assign t_r11_c21_7 = t_r11_c21_2 + t_r11_c21_3;
  assign t_r11_c21_8 = t_r11_c21_4 + p_12_20;
  assign t_r11_c21_9 = t_r11_c21_5 + t_r11_c21_6;
  assign t_r11_c21_10 = t_r11_c21_7 + t_r11_c21_8;
  assign t_r11_c21_11 = t_r11_c21_9 + t_r11_c21_10;
  assign t_r11_c21_12 = t_r11_c21_11 + p_12_22;
  assign out_11_21 = t_r11_c21_12 >> 4;

  assign t_r11_c22_0 = p_10_22 << 1;
  assign t_r11_c22_1 = p_11_21 << 1;
  assign t_r11_c22_2 = p_11_22 << 2;
  assign t_r11_c22_3 = p_11_23 << 1;
  assign t_r11_c22_4 = p_12_22 << 1;
  assign t_r11_c22_5 = t_r11_c22_0 + p_10_21;
  assign t_r11_c22_6 = t_r11_c22_1 + p_10_23;
  assign t_r11_c22_7 = t_r11_c22_2 + t_r11_c22_3;
  assign t_r11_c22_8 = t_r11_c22_4 + p_12_21;
  assign t_r11_c22_9 = t_r11_c22_5 + t_r11_c22_6;
  assign t_r11_c22_10 = t_r11_c22_7 + t_r11_c22_8;
  assign t_r11_c22_11 = t_r11_c22_9 + t_r11_c22_10;
  assign t_r11_c22_12 = t_r11_c22_11 + p_12_23;
  assign out_11_22 = t_r11_c22_12 >> 4;

  assign t_r11_c23_0 = p_10_23 << 1;
  assign t_r11_c23_1 = p_11_22 << 1;
  assign t_r11_c23_2 = p_11_23 << 2;
  assign t_r11_c23_3 = p_11_24 << 1;
  assign t_r11_c23_4 = p_12_23 << 1;
  assign t_r11_c23_5 = t_r11_c23_0 + p_10_22;
  assign t_r11_c23_6 = t_r11_c23_1 + p_10_24;
  assign t_r11_c23_7 = t_r11_c23_2 + t_r11_c23_3;
  assign t_r11_c23_8 = t_r11_c23_4 + p_12_22;
  assign t_r11_c23_9 = t_r11_c23_5 + t_r11_c23_6;
  assign t_r11_c23_10 = t_r11_c23_7 + t_r11_c23_8;
  assign t_r11_c23_11 = t_r11_c23_9 + t_r11_c23_10;
  assign t_r11_c23_12 = t_r11_c23_11 + p_12_24;
  assign out_11_23 = t_r11_c23_12 >> 4;

  assign t_r11_c24_0 = p_10_24 << 1;
  assign t_r11_c24_1 = p_11_23 << 1;
  assign t_r11_c24_2 = p_11_24 << 2;
  assign t_r11_c24_3 = p_11_25 << 1;
  assign t_r11_c24_4 = p_12_24 << 1;
  assign t_r11_c24_5 = t_r11_c24_0 + p_10_23;
  assign t_r11_c24_6 = t_r11_c24_1 + p_10_25;
  assign t_r11_c24_7 = t_r11_c24_2 + t_r11_c24_3;
  assign t_r11_c24_8 = t_r11_c24_4 + p_12_23;
  assign t_r11_c24_9 = t_r11_c24_5 + t_r11_c24_6;
  assign t_r11_c24_10 = t_r11_c24_7 + t_r11_c24_8;
  assign t_r11_c24_11 = t_r11_c24_9 + t_r11_c24_10;
  assign t_r11_c24_12 = t_r11_c24_11 + p_12_25;
  assign out_11_24 = t_r11_c24_12 >> 4;

  assign t_r11_c25_0 = p_10_25 << 1;
  assign t_r11_c25_1 = p_11_24 << 1;
  assign t_r11_c25_2 = p_11_25 << 2;
  assign t_r11_c25_3 = p_11_26 << 1;
  assign t_r11_c25_4 = p_12_25 << 1;
  assign t_r11_c25_5 = t_r11_c25_0 + p_10_24;
  assign t_r11_c25_6 = t_r11_c25_1 + p_10_26;
  assign t_r11_c25_7 = t_r11_c25_2 + t_r11_c25_3;
  assign t_r11_c25_8 = t_r11_c25_4 + p_12_24;
  assign t_r11_c25_9 = t_r11_c25_5 + t_r11_c25_6;
  assign t_r11_c25_10 = t_r11_c25_7 + t_r11_c25_8;
  assign t_r11_c25_11 = t_r11_c25_9 + t_r11_c25_10;
  assign t_r11_c25_12 = t_r11_c25_11 + p_12_26;
  assign out_11_25 = t_r11_c25_12 >> 4;

  assign t_r11_c26_0 = p_10_26 << 1;
  assign t_r11_c26_1 = p_11_25 << 1;
  assign t_r11_c26_2 = p_11_26 << 2;
  assign t_r11_c26_3 = p_11_27 << 1;
  assign t_r11_c26_4 = p_12_26 << 1;
  assign t_r11_c26_5 = t_r11_c26_0 + p_10_25;
  assign t_r11_c26_6 = t_r11_c26_1 + p_10_27;
  assign t_r11_c26_7 = t_r11_c26_2 + t_r11_c26_3;
  assign t_r11_c26_8 = t_r11_c26_4 + p_12_25;
  assign t_r11_c26_9 = t_r11_c26_5 + t_r11_c26_6;
  assign t_r11_c26_10 = t_r11_c26_7 + t_r11_c26_8;
  assign t_r11_c26_11 = t_r11_c26_9 + t_r11_c26_10;
  assign t_r11_c26_12 = t_r11_c26_11 + p_12_27;
  assign out_11_26 = t_r11_c26_12 >> 4;

  assign t_r11_c27_0 = p_10_27 << 1;
  assign t_r11_c27_1 = p_11_26 << 1;
  assign t_r11_c27_2 = p_11_27 << 2;
  assign t_r11_c27_3 = p_11_28 << 1;
  assign t_r11_c27_4 = p_12_27 << 1;
  assign t_r11_c27_5 = t_r11_c27_0 + p_10_26;
  assign t_r11_c27_6 = t_r11_c27_1 + p_10_28;
  assign t_r11_c27_7 = t_r11_c27_2 + t_r11_c27_3;
  assign t_r11_c27_8 = t_r11_c27_4 + p_12_26;
  assign t_r11_c27_9 = t_r11_c27_5 + t_r11_c27_6;
  assign t_r11_c27_10 = t_r11_c27_7 + t_r11_c27_8;
  assign t_r11_c27_11 = t_r11_c27_9 + t_r11_c27_10;
  assign t_r11_c27_12 = t_r11_c27_11 + p_12_28;
  assign out_11_27 = t_r11_c27_12 >> 4;

  assign t_r11_c28_0 = p_10_28 << 1;
  assign t_r11_c28_1 = p_11_27 << 1;
  assign t_r11_c28_2 = p_11_28 << 2;
  assign t_r11_c28_3 = p_11_29 << 1;
  assign t_r11_c28_4 = p_12_28 << 1;
  assign t_r11_c28_5 = t_r11_c28_0 + p_10_27;
  assign t_r11_c28_6 = t_r11_c28_1 + p_10_29;
  assign t_r11_c28_7 = t_r11_c28_2 + t_r11_c28_3;
  assign t_r11_c28_8 = t_r11_c28_4 + p_12_27;
  assign t_r11_c28_9 = t_r11_c28_5 + t_r11_c28_6;
  assign t_r11_c28_10 = t_r11_c28_7 + t_r11_c28_8;
  assign t_r11_c28_11 = t_r11_c28_9 + t_r11_c28_10;
  assign t_r11_c28_12 = t_r11_c28_11 + p_12_29;
  assign out_11_28 = t_r11_c28_12 >> 4;

  assign t_r11_c29_0 = p_10_29 << 1;
  assign t_r11_c29_1 = p_11_28 << 1;
  assign t_r11_c29_2 = p_11_29 << 2;
  assign t_r11_c29_3 = p_11_30 << 1;
  assign t_r11_c29_4 = p_12_29 << 1;
  assign t_r11_c29_5 = t_r11_c29_0 + p_10_28;
  assign t_r11_c29_6 = t_r11_c29_1 + p_10_30;
  assign t_r11_c29_7 = t_r11_c29_2 + t_r11_c29_3;
  assign t_r11_c29_8 = t_r11_c29_4 + p_12_28;
  assign t_r11_c29_9 = t_r11_c29_5 + t_r11_c29_6;
  assign t_r11_c29_10 = t_r11_c29_7 + t_r11_c29_8;
  assign t_r11_c29_11 = t_r11_c29_9 + t_r11_c29_10;
  assign t_r11_c29_12 = t_r11_c29_11 + p_12_30;
  assign out_11_29 = t_r11_c29_12 >> 4;

  assign t_r11_c30_0 = p_10_30 << 1;
  assign t_r11_c30_1 = p_11_29 << 1;
  assign t_r11_c30_2 = p_11_30 << 2;
  assign t_r11_c30_3 = p_11_31 << 1;
  assign t_r11_c30_4 = p_12_30 << 1;
  assign t_r11_c30_5 = t_r11_c30_0 + p_10_29;
  assign t_r11_c30_6 = t_r11_c30_1 + p_10_31;
  assign t_r11_c30_7 = t_r11_c30_2 + t_r11_c30_3;
  assign t_r11_c30_8 = t_r11_c30_4 + p_12_29;
  assign t_r11_c30_9 = t_r11_c30_5 + t_r11_c30_6;
  assign t_r11_c30_10 = t_r11_c30_7 + t_r11_c30_8;
  assign t_r11_c30_11 = t_r11_c30_9 + t_r11_c30_10;
  assign t_r11_c30_12 = t_r11_c30_11 + p_12_31;
  assign out_11_30 = t_r11_c30_12 >> 4;

  assign t_r11_c31_0 = p_10_31 << 1;
  assign t_r11_c31_1 = p_11_30 << 1;
  assign t_r11_c31_2 = p_11_31 << 2;
  assign t_r11_c31_3 = p_11_32 << 1;
  assign t_r11_c31_4 = p_12_31 << 1;
  assign t_r11_c31_5 = t_r11_c31_0 + p_10_30;
  assign t_r11_c31_6 = t_r11_c31_1 + p_10_32;
  assign t_r11_c31_7 = t_r11_c31_2 + t_r11_c31_3;
  assign t_r11_c31_8 = t_r11_c31_4 + p_12_30;
  assign t_r11_c31_9 = t_r11_c31_5 + t_r11_c31_6;
  assign t_r11_c31_10 = t_r11_c31_7 + t_r11_c31_8;
  assign t_r11_c31_11 = t_r11_c31_9 + t_r11_c31_10;
  assign t_r11_c31_12 = t_r11_c31_11 + p_12_32;
  assign out_11_31 = t_r11_c31_12 >> 4;

  assign t_r11_c32_0 = p_10_32 << 1;
  assign t_r11_c32_1 = p_11_31 << 1;
  assign t_r11_c32_2 = p_11_32 << 2;
  assign t_r11_c32_3 = p_11_33 << 1;
  assign t_r11_c32_4 = p_12_32 << 1;
  assign t_r11_c32_5 = t_r11_c32_0 + p_10_31;
  assign t_r11_c32_6 = t_r11_c32_1 + p_10_33;
  assign t_r11_c32_7 = t_r11_c32_2 + t_r11_c32_3;
  assign t_r11_c32_8 = t_r11_c32_4 + p_12_31;
  assign t_r11_c32_9 = t_r11_c32_5 + t_r11_c32_6;
  assign t_r11_c32_10 = t_r11_c32_7 + t_r11_c32_8;
  assign t_r11_c32_11 = t_r11_c32_9 + t_r11_c32_10;
  assign t_r11_c32_12 = t_r11_c32_11 + p_12_33;
  assign out_11_32 = t_r11_c32_12 >> 4;

  assign t_r11_c33_0 = p_10_33 << 1;
  assign t_r11_c33_1 = p_11_32 << 1;
  assign t_r11_c33_2 = p_11_33 << 2;
  assign t_r11_c33_3 = p_11_34 << 1;
  assign t_r11_c33_4 = p_12_33 << 1;
  assign t_r11_c33_5 = t_r11_c33_0 + p_10_32;
  assign t_r11_c33_6 = t_r11_c33_1 + p_10_34;
  assign t_r11_c33_7 = t_r11_c33_2 + t_r11_c33_3;
  assign t_r11_c33_8 = t_r11_c33_4 + p_12_32;
  assign t_r11_c33_9 = t_r11_c33_5 + t_r11_c33_6;
  assign t_r11_c33_10 = t_r11_c33_7 + t_r11_c33_8;
  assign t_r11_c33_11 = t_r11_c33_9 + t_r11_c33_10;
  assign t_r11_c33_12 = t_r11_c33_11 + p_12_34;
  assign out_11_33 = t_r11_c33_12 >> 4;

  assign t_r11_c34_0 = p_10_34 << 1;
  assign t_r11_c34_1 = p_11_33 << 1;
  assign t_r11_c34_2 = p_11_34 << 2;
  assign t_r11_c34_3 = p_11_35 << 1;
  assign t_r11_c34_4 = p_12_34 << 1;
  assign t_r11_c34_5 = t_r11_c34_0 + p_10_33;
  assign t_r11_c34_6 = t_r11_c34_1 + p_10_35;
  assign t_r11_c34_7 = t_r11_c34_2 + t_r11_c34_3;
  assign t_r11_c34_8 = t_r11_c34_4 + p_12_33;
  assign t_r11_c34_9 = t_r11_c34_5 + t_r11_c34_6;
  assign t_r11_c34_10 = t_r11_c34_7 + t_r11_c34_8;
  assign t_r11_c34_11 = t_r11_c34_9 + t_r11_c34_10;
  assign t_r11_c34_12 = t_r11_c34_11 + p_12_35;
  assign out_11_34 = t_r11_c34_12 >> 4;

  assign t_r11_c35_0 = p_10_35 << 1;
  assign t_r11_c35_1 = p_11_34 << 1;
  assign t_r11_c35_2 = p_11_35 << 2;
  assign t_r11_c35_3 = p_11_36 << 1;
  assign t_r11_c35_4 = p_12_35 << 1;
  assign t_r11_c35_5 = t_r11_c35_0 + p_10_34;
  assign t_r11_c35_6 = t_r11_c35_1 + p_10_36;
  assign t_r11_c35_7 = t_r11_c35_2 + t_r11_c35_3;
  assign t_r11_c35_8 = t_r11_c35_4 + p_12_34;
  assign t_r11_c35_9 = t_r11_c35_5 + t_r11_c35_6;
  assign t_r11_c35_10 = t_r11_c35_7 + t_r11_c35_8;
  assign t_r11_c35_11 = t_r11_c35_9 + t_r11_c35_10;
  assign t_r11_c35_12 = t_r11_c35_11 + p_12_36;
  assign out_11_35 = t_r11_c35_12 >> 4;

  assign t_r11_c36_0 = p_10_36 << 1;
  assign t_r11_c36_1 = p_11_35 << 1;
  assign t_r11_c36_2 = p_11_36 << 2;
  assign t_r11_c36_3 = p_11_37 << 1;
  assign t_r11_c36_4 = p_12_36 << 1;
  assign t_r11_c36_5 = t_r11_c36_0 + p_10_35;
  assign t_r11_c36_6 = t_r11_c36_1 + p_10_37;
  assign t_r11_c36_7 = t_r11_c36_2 + t_r11_c36_3;
  assign t_r11_c36_8 = t_r11_c36_4 + p_12_35;
  assign t_r11_c36_9 = t_r11_c36_5 + t_r11_c36_6;
  assign t_r11_c36_10 = t_r11_c36_7 + t_r11_c36_8;
  assign t_r11_c36_11 = t_r11_c36_9 + t_r11_c36_10;
  assign t_r11_c36_12 = t_r11_c36_11 + p_12_37;
  assign out_11_36 = t_r11_c36_12 >> 4;

  assign t_r11_c37_0 = p_10_37 << 1;
  assign t_r11_c37_1 = p_11_36 << 1;
  assign t_r11_c37_2 = p_11_37 << 2;
  assign t_r11_c37_3 = p_11_38 << 1;
  assign t_r11_c37_4 = p_12_37 << 1;
  assign t_r11_c37_5 = t_r11_c37_0 + p_10_36;
  assign t_r11_c37_6 = t_r11_c37_1 + p_10_38;
  assign t_r11_c37_7 = t_r11_c37_2 + t_r11_c37_3;
  assign t_r11_c37_8 = t_r11_c37_4 + p_12_36;
  assign t_r11_c37_9 = t_r11_c37_5 + t_r11_c37_6;
  assign t_r11_c37_10 = t_r11_c37_7 + t_r11_c37_8;
  assign t_r11_c37_11 = t_r11_c37_9 + t_r11_c37_10;
  assign t_r11_c37_12 = t_r11_c37_11 + p_12_38;
  assign out_11_37 = t_r11_c37_12 >> 4;

  assign t_r11_c38_0 = p_10_38 << 1;
  assign t_r11_c38_1 = p_11_37 << 1;
  assign t_r11_c38_2 = p_11_38 << 2;
  assign t_r11_c38_3 = p_11_39 << 1;
  assign t_r11_c38_4 = p_12_38 << 1;
  assign t_r11_c38_5 = t_r11_c38_0 + p_10_37;
  assign t_r11_c38_6 = t_r11_c38_1 + p_10_39;
  assign t_r11_c38_7 = t_r11_c38_2 + t_r11_c38_3;
  assign t_r11_c38_8 = t_r11_c38_4 + p_12_37;
  assign t_r11_c38_9 = t_r11_c38_5 + t_r11_c38_6;
  assign t_r11_c38_10 = t_r11_c38_7 + t_r11_c38_8;
  assign t_r11_c38_11 = t_r11_c38_9 + t_r11_c38_10;
  assign t_r11_c38_12 = t_r11_c38_11 + p_12_39;
  assign out_11_38 = t_r11_c38_12 >> 4;

  assign t_r11_c39_0 = p_10_39 << 1;
  assign t_r11_c39_1 = p_11_38 << 1;
  assign t_r11_c39_2 = p_11_39 << 2;
  assign t_r11_c39_3 = p_11_40 << 1;
  assign t_r11_c39_4 = p_12_39 << 1;
  assign t_r11_c39_5 = t_r11_c39_0 + p_10_38;
  assign t_r11_c39_6 = t_r11_c39_1 + p_10_40;
  assign t_r11_c39_7 = t_r11_c39_2 + t_r11_c39_3;
  assign t_r11_c39_8 = t_r11_c39_4 + p_12_38;
  assign t_r11_c39_9 = t_r11_c39_5 + t_r11_c39_6;
  assign t_r11_c39_10 = t_r11_c39_7 + t_r11_c39_8;
  assign t_r11_c39_11 = t_r11_c39_9 + t_r11_c39_10;
  assign t_r11_c39_12 = t_r11_c39_11 + p_12_40;
  assign out_11_39 = t_r11_c39_12 >> 4;

  assign t_r11_c40_0 = p_10_40 << 1;
  assign t_r11_c40_1 = p_11_39 << 1;
  assign t_r11_c40_2 = p_11_40 << 2;
  assign t_r11_c40_3 = p_11_41 << 1;
  assign t_r11_c40_4 = p_12_40 << 1;
  assign t_r11_c40_5 = t_r11_c40_0 + p_10_39;
  assign t_r11_c40_6 = t_r11_c40_1 + p_10_41;
  assign t_r11_c40_7 = t_r11_c40_2 + t_r11_c40_3;
  assign t_r11_c40_8 = t_r11_c40_4 + p_12_39;
  assign t_r11_c40_9 = t_r11_c40_5 + t_r11_c40_6;
  assign t_r11_c40_10 = t_r11_c40_7 + t_r11_c40_8;
  assign t_r11_c40_11 = t_r11_c40_9 + t_r11_c40_10;
  assign t_r11_c40_12 = t_r11_c40_11 + p_12_41;
  assign out_11_40 = t_r11_c40_12 >> 4;

  assign t_r11_c41_0 = p_10_41 << 1;
  assign t_r11_c41_1 = p_11_40 << 1;
  assign t_r11_c41_2 = p_11_41 << 2;
  assign t_r11_c41_3 = p_11_42 << 1;
  assign t_r11_c41_4 = p_12_41 << 1;
  assign t_r11_c41_5 = t_r11_c41_0 + p_10_40;
  assign t_r11_c41_6 = t_r11_c41_1 + p_10_42;
  assign t_r11_c41_7 = t_r11_c41_2 + t_r11_c41_3;
  assign t_r11_c41_8 = t_r11_c41_4 + p_12_40;
  assign t_r11_c41_9 = t_r11_c41_5 + t_r11_c41_6;
  assign t_r11_c41_10 = t_r11_c41_7 + t_r11_c41_8;
  assign t_r11_c41_11 = t_r11_c41_9 + t_r11_c41_10;
  assign t_r11_c41_12 = t_r11_c41_11 + p_12_42;
  assign out_11_41 = t_r11_c41_12 >> 4;

  assign t_r11_c42_0 = p_10_42 << 1;
  assign t_r11_c42_1 = p_11_41 << 1;
  assign t_r11_c42_2 = p_11_42 << 2;
  assign t_r11_c42_3 = p_11_43 << 1;
  assign t_r11_c42_4 = p_12_42 << 1;
  assign t_r11_c42_5 = t_r11_c42_0 + p_10_41;
  assign t_r11_c42_6 = t_r11_c42_1 + p_10_43;
  assign t_r11_c42_7 = t_r11_c42_2 + t_r11_c42_3;
  assign t_r11_c42_8 = t_r11_c42_4 + p_12_41;
  assign t_r11_c42_9 = t_r11_c42_5 + t_r11_c42_6;
  assign t_r11_c42_10 = t_r11_c42_7 + t_r11_c42_8;
  assign t_r11_c42_11 = t_r11_c42_9 + t_r11_c42_10;
  assign t_r11_c42_12 = t_r11_c42_11 + p_12_43;
  assign out_11_42 = t_r11_c42_12 >> 4;

  assign t_r11_c43_0 = p_10_43 << 1;
  assign t_r11_c43_1 = p_11_42 << 1;
  assign t_r11_c43_2 = p_11_43 << 2;
  assign t_r11_c43_3 = p_11_44 << 1;
  assign t_r11_c43_4 = p_12_43 << 1;
  assign t_r11_c43_5 = t_r11_c43_0 + p_10_42;
  assign t_r11_c43_6 = t_r11_c43_1 + p_10_44;
  assign t_r11_c43_7 = t_r11_c43_2 + t_r11_c43_3;
  assign t_r11_c43_8 = t_r11_c43_4 + p_12_42;
  assign t_r11_c43_9 = t_r11_c43_5 + t_r11_c43_6;
  assign t_r11_c43_10 = t_r11_c43_7 + t_r11_c43_8;
  assign t_r11_c43_11 = t_r11_c43_9 + t_r11_c43_10;
  assign t_r11_c43_12 = t_r11_c43_11 + p_12_44;
  assign out_11_43 = t_r11_c43_12 >> 4;

  assign t_r11_c44_0 = p_10_44 << 1;
  assign t_r11_c44_1 = p_11_43 << 1;
  assign t_r11_c44_2 = p_11_44 << 2;
  assign t_r11_c44_3 = p_11_45 << 1;
  assign t_r11_c44_4 = p_12_44 << 1;
  assign t_r11_c44_5 = t_r11_c44_0 + p_10_43;
  assign t_r11_c44_6 = t_r11_c44_1 + p_10_45;
  assign t_r11_c44_7 = t_r11_c44_2 + t_r11_c44_3;
  assign t_r11_c44_8 = t_r11_c44_4 + p_12_43;
  assign t_r11_c44_9 = t_r11_c44_5 + t_r11_c44_6;
  assign t_r11_c44_10 = t_r11_c44_7 + t_r11_c44_8;
  assign t_r11_c44_11 = t_r11_c44_9 + t_r11_c44_10;
  assign t_r11_c44_12 = t_r11_c44_11 + p_12_45;
  assign out_11_44 = t_r11_c44_12 >> 4;

  assign t_r11_c45_0 = p_10_45 << 1;
  assign t_r11_c45_1 = p_11_44 << 1;
  assign t_r11_c45_2 = p_11_45 << 2;
  assign t_r11_c45_3 = p_11_46 << 1;
  assign t_r11_c45_4 = p_12_45 << 1;
  assign t_r11_c45_5 = t_r11_c45_0 + p_10_44;
  assign t_r11_c45_6 = t_r11_c45_1 + p_10_46;
  assign t_r11_c45_7 = t_r11_c45_2 + t_r11_c45_3;
  assign t_r11_c45_8 = t_r11_c45_4 + p_12_44;
  assign t_r11_c45_9 = t_r11_c45_5 + t_r11_c45_6;
  assign t_r11_c45_10 = t_r11_c45_7 + t_r11_c45_8;
  assign t_r11_c45_11 = t_r11_c45_9 + t_r11_c45_10;
  assign t_r11_c45_12 = t_r11_c45_11 + p_12_46;
  assign out_11_45 = t_r11_c45_12 >> 4;

  assign t_r11_c46_0 = p_10_46 << 1;
  assign t_r11_c46_1 = p_11_45 << 1;
  assign t_r11_c46_2 = p_11_46 << 2;
  assign t_r11_c46_3 = p_11_47 << 1;
  assign t_r11_c46_4 = p_12_46 << 1;
  assign t_r11_c46_5 = t_r11_c46_0 + p_10_45;
  assign t_r11_c46_6 = t_r11_c46_1 + p_10_47;
  assign t_r11_c46_7 = t_r11_c46_2 + t_r11_c46_3;
  assign t_r11_c46_8 = t_r11_c46_4 + p_12_45;
  assign t_r11_c46_9 = t_r11_c46_5 + t_r11_c46_6;
  assign t_r11_c46_10 = t_r11_c46_7 + t_r11_c46_8;
  assign t_r11_c46_11 = t_r11_c46_9 + t_r11_c46_10;
  assign t_r11_c46_12 = t_r11_c46_11 + p_12_47;
  assign out_11_46 = t_r11_c46_12 >> 4;

  assign t_r11_c47_0 = p_10_47 << 1;
  assign t_r11_c47_1 = p_11_46 << 1;
  assign t_r11_c47_2 = p_11_47 << 2;
  assign t_r11_c47_3 = p_11_48 << 1;
  assign t_r11_c47_4 = p_12_47 << 1;
  assign t_r11_c47_5 = t_r11_c47_0 + p_10_46;
  assign t_r11_c47_6 = t_r11_c47_1 + p_10_48;
  assign t_r11_c47_7 = t_r11_c47_2 + t_r11_c47_3;
  assign t_r11_c47_8 = t_r11_c47_4 + p_12_46;
  assign t_r11_c47_9 = t_r11_c47_5 + t_r11_c47_6;
  assign t_r11_c47_10 = t_r11_c47_7 + t_r11_c47_8;
  assign t_r11_c47_11 = t_r11_c47_9 + t_r11_c47_10;
  assign t_r11_c47_12 = t_r11_c47_11 + p_12_48;
  assign out_11_47 = t_r11_c47_12 >> 4;

  assign t_r11_c48_0 = p_10_48 << 1;
  assign t_r11_c48_1 = p_11_47 << 1;
  assign t_r11_c48_2 = p_11_48 << 2;
  assign t_r11_c48_3 = p_11_49 << 1;
  assign t_r11_c48_4 = p_12_48 << 1;
  assign t_r11_c48_5 = t_r11_c48_0 + p_10_47;
  assign t_r11_c48_6 = t_r11_c48_1 + p_10_49;
  assign t_r11_c48_7 = t_r11_c48_2 + t_r11_c48_3;
  assign t_r11_c48_8 = t_r11_c48_4 + p_12_47;
  assign t_r11_c48_9 = t_r11_c48_5 + t_r11_c48_6;
  assign t_r11_c48_10 = t_r11_c48_7 + t_r11_c48_8;
  assign t_r11_c48_11 = t_r11_c48_9 + t_r11_c48_10;
  assign t_r11_c48_12 = t_r11_c48_11 + p_12_49;
  assign out_11_48 = t_r11_c48_12 >> 4;

  assign t_r11_c49_0 = p_10_49 << 1;
  assign t_r11_c49_1 = p_11_48 << 1;
  assign t_r11_c49_2 = p_11_49 << 2;
  assign t_r11_c49_3 = p_11_50 << 1;
  assign t_r11_c49_4 = p_12_49 << 1;
  assign t_r11_c49_5 = t_r11_c49_0 + p_10_48;
  assign t_r11_c49_6 = t_r11_c49_1 + p_10_50;
  assign t_r11_c49_7 = t_r11_c49_2 + t_r11_c49_3;
  assign t_r11_c49_8 = t_r11_c49_4 + p_12_48;
  assign t_r11_c49_9 = t_r11_c49_5 + t_r11_c49_6;
  assign t_r11_c49_10 = t_r11_c49_7 + t_r11_c49_8;
  assign t_r11_c49_11 = t_r11_c49_9 + t_r11_c49_10;
  assign t_r11_c49_12 = t_r11_c49_11 + p_12_50;
  assign out_11_49 = t_r11_c49_12 >> 4;

  assign t_r11_c50_0 = p_10_50 << 1;
  assign t_r11_c50_1 = p_11_49 << 1;
  assign t_r11_c50_2 = p_11_50 << 2;
  assign t_r11_c50_3 = p_11_51 << 1;
  assign t_r11_c50_4 = p_12_50 << 1;
  assign t_r11_c50_5 = t_r11_c50_0 + p_10_49;
  assign t_r11_c50_6 = t_r11_c50_1 + p_10_51;
  assign t_r11_c50_7 = t_r11_c50_2 + t_r11_c50_3;
  assign t_r11_c50_8 = t_r11_c50_4 + p_12_49;
  assign t_r11_c50_9 = t_r11_c50_5 + t_r11_c50_6;
  assign t_r11_c50_10 = t_r11_c50_7 + t_r11_c50_8;
  assign t_r11_c50_11 = t_r11_c50_9 + t_r11_c50_10;
  assign t_r11_c50_12 = t_r11_c50_11 + p_12_51;
  assign out_11_50 = t_r11_c50_12 >> 4;

  assign t_r11_c51_0 = p_10_51 << 1;
  assign t_r11_c51_1 = p_11_50 << 1;
  assign t_r11_c51_2 = p_11_51 << 2;
  assign t_r11_c51_3 = p_11_52 << 1;
  assign t_r11_c51_4 = p_12_51 << 1;
  assign t_r11_c51_5 = t_r11_c51_0 + p_10_50;
  assign t_r11_c51_6 = t_r11_c51_1 + p_10_52;
  assign t_r11_c51_7 = t_r11_c51_2 + t_r11_c51_3;
  assign t_r11_c51_8 = t_r11_c51_4 + p_12_50;
  assign t_r11_c51_9 = t_r11_c51_5 + t_r11_c51_6;
  assign t_r11_c51_10 = t_r11_c51_7 + t_r11_c51_8;
  assign t_r11_c51_11 = t_r11_c51_9 + t_r11_c51_10;
  assign t_r11_c51_12 = t_r11_c51_11 + p_12_52;
  assign out_11_51 = t_r11_c51_12 >> 4;

  assign t_r11_c52_0 = p_10_52 << 1;
  assign t_r11_c52_1 = p_11_51 << 1;
  assign t_r11_c52_2 = p_11_52 << 2;
  assign t_r11_c52_3 = p_11_53 << 1;
  assign t_r11_c52_4 = p_12_52 << 1;
  assign t_r11_c52_5 = t_r11_c52_0 + p_10_51;
  assign t_r11_c52_6 = t_r11_c52_1 + p_10_53;
  assign t_r11_c52_7 = t_r11_c52_2 + t_r11_c52_3;
  assign t_r11_c52_8 = t_r11_c52_4 + p_12_51;
  assign t_r11_c52_9 = t_r11_c52_5 + t_r11_c52_6;
  assign t_r11_c52_10 = t_r11_c52_7 + t_r11_c52_8;
  assign t_r11_c52_11 = t_r11_c52_9 + t_r11_c52_10;
  assign t_r11_c52_12 = t_r11_c52_11 + p_12_53;
  assign out_11_52 = t_r11_c52_12 >> 4;

  assign t_r11_c53_0 = p_10_53 << 1;
  assign t_r11_c53_1 = p_11_52 << 1;
  assign t_r11_c53_2 = p_11_53 << 2;
  assign t_r11_c53_3 = p_11_54 << 1;
  assign t_r11_c53_4 = p_12_53 << 1;
  assign t_r11_c53_5 = t_r11_c53_0 + p_10_52;
  assign t_r11_c53_6 = t_r11_c53_1 + p_10_54;
  assign t_r11_c53_7 = t_r11_c53_2 + t_r11_c53_3;
  assign t_r11_c53_8 = t_r11_c53_4 + p_12_52;
  assign t_r11_c53_9 = t_r11_c53_5 + t_r11_c53_6;
  assign t_r11_c53_10 = t_r11_c53_7 + t_r11_c53_8;
  assign t_r11_c53_11 = t_r11_c53_9 + t_r11_c53_10;
  assign t_r11_c53_12 = t_r11_c53_11 + p_12_54;
  assign out_11_53 = t_r11_c53_12 >> 4;

  assign t_r11_c54_0 = p_10_54 << 1;
  assign t_r11_c54_1 = p_11_53 << 1;
  assign t_r11_c54_2 = p_11_54 << 2;
  assign t_r11_c54_3 = p_11_55 << 1;
  assign t_r11_c54_4 = p_12_54 << 1;
  assign t_r11_c54_5 = t_r11_c54_0 + p_10_53;
  assign t_r11_c54_6 = t_r11_c54_1 + p_10_55;
  assign t_r11_c54_7 = t_r11_c54_2 + t_r11_c54_3;
  assign t_r11_c54_8 = t_r11_c54_4 + p_12_53;
  assign t_r11_c54_9 = t_r11_c54_5 + t_r11_c54_6;
  assign t_r11_c54_10 = t_r11_c54_7 + t_r11_c54_8;
  assign t_r11_c54_11 = t_r11_c54_9 + t_r11_c54_10;
  assign t_r11_c54_12 = t_r11_c54_11 + p_12_55;
  assign out_11_54 = t_r11_c54_12 >> 4;

  assign t_r11_c55_0 = p_10_55 << 1;
  assign t_r11_c55_1 = p_11_54 << 1;
  assign t_r11_c55_2 = p_11_55 << 2;
  assign t_r11_c55_3 = p_11_56 << 1;
  assign t_r11_c55_4 = p_12_55 << 1;
  assign t_r11_c55_5 = t_r11_c55_0 + p_10_54;
  assign t_r11_c55_6 = t_r11_c55_1 + p_10_56;
  assign t_r11_c55_7 = t_r11_c55_2 + t_r11_c55_3;
  assign t_r11_c55_8 = t_r11_c55_4 + p_12_54;
  assign t_r11_c55_9 = t_r11_c55_5 + t_r11_c55_6;
  assign t_r11_c55_10 = t_r11_c55_7 + t_r11_c55_8;
  assign t_r11_c55_11 = t_r11_c55_9 + t_r11_c55_10;
  assign t_r11_c55_12 = t_r11_c55_11 + p_12_56;
  assign out_11_55 = t_r11_c55_12 >> 4;

  assign t_r11_c56_0 = p_10_56 << 1;
  assign t_r11_c56_1 = p_11_55 << 1;
  assign t_r11_c56_2 = p_11_56 << 2;
  assign t_r11_c56_3 = p_11_57 << 1;
  assign t_r11_c56_4 = p_12_56 << 1;
  assign t_r11_c56_5 = t_r11_c56_0 + p_10_55;
  assign t_r11_c56_6 = t_r11_c56_1 + p_10_57;
  assign t_r11_c56_7 = t_r11_c56_2 + t_r11_c56_3;
  assign t_r11_c56_8 = t_r11_c56_4 + p_12_55;
  assign t_r11_c56_9 = t_r11_c56_5 + t_r11_c56_6;
  assign t_r11_c56_10 = t_r11_c56_7 + t_r11_c56_8;
  assign t_r11_c56_11 = t_r11_c56_9 + t_r11_c56_10;
  assign t_r11_c56_12 = t_r11_c56_11 + p_12_57;
  assign out_11_56 = t_r11_c56_12 >> 4;

  assign t_r11_c57_0 = p_10_57 << 1;
  assign t_r11_c57_1 = p_11_56 << 1;
  assign t_r11_c57_2 = p_11_57 << 2;
  assign t_r11_c57_3 = p_11_58 << 1;
  assign t_r11_c57_4 = p_12_57 << 1;
  assign t_r11_c57_5 = t_r11_c57_0 + p_10_56;
  assign t_r11_c57_6 = t_r11_c57_1 + p_10_58;
  assign t_r11_c57_7 = t_r11_c57_2 + t_r11_c57_3;
  assign t_r11_c57_8 = t_r11_c57_4 + p_12_56;
  assign t_r11_c57_9 = t_r11_c57_5 + t_r11_c57_6;
  assign t_r11_c57_10 = t_r11_c57_7 + t_r11_c57_8;
  assign t_r11_c57_11 = t_r11_c57_9 + t_r11_c57_10;
  assign t_r11_c57_12 = t_r11_c57_11 + p_12_58;
  assign out_11_57 = t_r11_c57_12 >> 4;

  assign t_r11_c58_0 = p_10_58 << 1;
  assign t_r11_c58_1 = p_11_57 << 1;
  assign t_r11_c58_2 = p_11_58 << 2;
  assign t_r11_c58_3 = p_11_59 << 1;
  assign t_r11_c58_4 = p_12_58 << 1;
  assign t_r11_c58_5 = t_r11_c58_0 + p_10_57;
  assign t_r11_c58_6 = t_r11_c58_1 + p_10_59;
  assign t_r11_c58_7 = t_r11_c58_2 + t_r11_c58_3;
  assign t_r11_c58_8 = t_r11_c58_4 + p_12_57;
  assign t_r11_c58_9 = t_r11_c58_5 + t_r11_c58_6;
  assign t_r11_c58_10 = t_r11_c58_7 + t_r11_c58_8;
  assign t_r11_c58_11 = t_r11_c58_9 + t_r11_c58_10;
  assign t_r11_c58_12 = t_r11_c58_11 + p_12_59;
  assign out_11_58 = t_r11_c58_12 >> 4;

  assign t_r11_c59_0 = p_10_59 << 1;
  assign t_r11_c59_1 = p_11_58 << 1;
  assign t_r11_c59_2 = p_11_59 << 2;
  assign t_r11_c59_3 = p_11_60 << 1;
  assign t_r11_c59_4 = p_12_59 << 1;
  assign t_r11_c59_5 = t_r11_c59_0 + p_10_58;
  assign t_r11_c59_6 = t_r11_c59_1 + p_10_60;
  assign t_r11_c59_7 = t_r11_c59_2 + t_r11_c59_3;
  assign t_r11_c59_8 = t_r11_c59_4 + p_12_58;
  assign t_r11_c59_9 = t_r11_c59_5 + t_r11_c59_6;
  assign t_r11_c59_10 = t_r11_c59_7 + t_r11_c59_8;
  assign t_r11_c59_11 = t_r11_c59_9 + t_r11_c59_10;
  assign t_r11_c59_12 = t_r11_c59_11 + p_12_60;
  assign out_11_59 = t_r11_c59_12 >> 4;

  assign t_r11_c60_0 = p_10_60 << 1;
  assign t_r11_c60_1 = p_11_59 << 1;
  assign t_r11_c60_2 = p_11_60 << 2;
  assign t_r11_c60_3 = p_11_61 << 1;
  assign t_r11_c60_4 = p_12_60 << 1;
  assign t_r11_c60_5 = t_r11_c60_0 + p_10_59;
  assign t_r11_c60_6 = t_r11_c60_1 + p_10_61;
  assign t_r11_c60_7 = t_r11_c60_2 + t_r11_c60_3;
  assign t_r11_c60_8 = t_r11_c60_4 + p_12_59;
  assign t_r11_c60_9 = t_r11_c60_5 + t_r11_c60_6;
  assign t_r11_c60_10 = t_r11_c60_7 + t_r11_c60_8;
  assign t_r11_c60_11 = t_r11_c60_9 + t_r11_c60_10;
  assign t_r11_c60_12 = t_r11_c60_11 + p_12_61;
  assign out_11_60 = t_r11_c60_12 >> 4;

  assign t_r11_c61_0 = p_10_61 << 1;
  assign t_r11_c61_1 = p_11_60 << 1;
  assign t_r11_c61_2 = p_11_61 << 2;
  assign t_r11_c61_3 = p_11_62 << 1;
  assign t_r11_c61_4 = p_12_61 << 1;
  assign t_r11_c61_5 = t_r11_c61_0 + p_10_60;
  assign t_r11_c61_6 = t_r11_c61_1 + p_10_62;
  assign t_r11_c61_7 = t_r11_c61_2 + t_r11_c61_3;
  assign t_r11_c61_8 = t_r11_c61_4 + p_12_60;
  assign t_r11_c61_9 = t_r11_c61_5 + t_r11_c61_6;
  assign t_r11_c61_10 = t_r11_c61_7 + t_r11_c61_8;
  assign t_r11_c61_11 = t_r11_c61_9 + t_r11_c61_10;
  assign t_r11_c61_12 = t_r11_c61_11 + p_12_62;
  assign out_11_61 = t_r11_c61_12 >> 4;

  assign t_r11_c62_0 = p_10_62 << 1;
  assign t_r11_c62_1 = p_11_61 << 1;
  assign t_r11_c62_2 = p_11_62 << 2;
  assign t_r11_c62_3 = p_11_63 << 1;
  assign t_r11_c62_4 = p_12_62 << 1;
  assign t_r11_c62_5 = t_r11_c62_0 + p_10_61;
  assign t_r11_c62_6 = t_r11_c62_1 + p_10_63;
  assign t_r11_c62_7 = t_r11_c62_2 + t_r11_c62_3;
  assign t_r11_c62_8 = t_r11_c62_4 + p_12_61;
  assign t_r11_c62_9 = t_r11_c62_5 + t_r11_c62_6;
  assign t_r11_c62_10 = t_r11_c62_7 + t_r11_c62_8;
  assign t_r11_c62_11 = t_r11_c62_9 + t_r11_c62_10;
  assign t_r11_c62_12 = t_r11_c62_11 + p_12_63;
  assign out_11_62 = t_r11_c62_12 >> 4;

  assign t_r11_c63_0 = p_10_63 << 1;
  assign t_r11_c63_1 = p_11_62 << 1;
  assign t_r11_c63_2 = p_11_63 << 2;
  assign t_r11_c63_3 = p_11_64 << 1;
  assign t_r11_c63_4 = p_12_63 << 1;
  assign t_r11_c63_5 = t_r11_c63_0 + p_10_62;
  assign t_r11_c63_6 = t_r11_c63_1 + p_10_64;
  assign t_r11_c63_7 = t_r11_c63_2 + t_r11_c63_3;
  assign t_r11_c63_8 = t_r11_c63_4 + p_12_62;
  assign t_r11_c63_9 = t_r11_c63_5 + t_r11_c63_6;
  assign t_r11_c63_10 = t_r11_c63_7 + t_r11_c63_8;
  assign t_r11_c63_11 = t_r11_c63_9 + t_r11_c63_10;
  assign t_r11_c63_12 = t_r11_c63_11 + p_12_64;
  assign out_11_63 = t_r11_c63_12 >> 4;

  assign t_r11_c64_0 = p_10_64 << 1;
  assign t_r11_c64_1 = p_11_63 << 1;
  assign t_r11_c64_2 = p_11_64 << 2;
  assign t_r11_c64_3 = p_11_65 << 1;
  assign t_r11_c64_4 = p_12_64 << 1;
  assign t_r11_c64_5 = t_r11_c64_0 + p_10_63;
  assign t_r11_c64_6 = t_r11_c64_1 + p_10_65;
  assign t_r11_c64_7 = t_r11_c64_2 + t_r11_c64_3;
  assign t_r11_c64_8 = t_r11_c64_4 + p_12_63;
  assign t_r11_c64_9 = t_r11_c64_5 + t_r11_c64_6;
  assign t_r11_c64_10 = t_r11_c64_7 + t_r11_c64_8;
  assign t_r11_c64_11 = t_r11_c64_9 + t_r11_c64_10;
  assign t_r11_c64_12 = t_r11_c64_11 + p_12_65;
  assign out_11_64 = t_r11_c64_12 >> 4;

  assign t_r12_c1_0 = p_11_1 << 1;
  assign t_r12_c1_1 = p_12_0 << 1;
  assign t_r12_c1_2 = p_12_1 << 2;
  assign t_r12_c1_3 = p_12_2 << 1;
  assign t_r12_c1_4 = p_13_1 << 1;
  assign t_r12_c1_5 = t_r12_c1_0 + p_11_0;
  assign t_r12_c1_6 = t_r12_c1_1 + p_11_2;
  assign t_r12_c1_7 = t_r12_c1_2 + t_r12_c1_3;
  assign t_r12_c1_8 = t_r12_c1_4 + p_13_0;
  assign t_r12_c1_9 = t_r12_c1_5 + t_r12_c1_6;
  assign t_r12_c1_10 = t_r12_c1_7 + t_r12_c1_8;
  assign t_r12_c1_11 = t_r12_c1_9 + t_r12_c1_10;
  assign t_r12_c1_12 = t_r12_c1_11 + p_13_2;
  assign out_12_1 = t_r12_c1_12 >> 4;

  assign t_r12_c2_0 = p_11_2 << 1;
  assign t_r12_c2_1 = p_12_1 << 1;
  assign t_r12_c2_2 = p_12_2 << 2;
  assign t_r12_c2_3 = p_12_3 << 1;
  assign t_r12_c2_4 = p_13_2 << 1;
  assign t_r12_c2_5 = t_r12_c2_0 + p_11_1;
  assign t_r12_c2_6 = t_r12_c2_1 + p_11_3;
  assign t_r12_c2_7 = t_r12_c2_2 + t_r12_c2_3;
  assign t_r12_c2_8 = t_r12_c2_4 + p_13_1;
  assign t_r12_c2_9 = t_r12_c2_5 + t_r12_c2_6;
  assign t_r12_c2_10 = t_r12_c2_7 + t_r12_c2_8;
  assign t_r12_c2_11 = t_r12_c2_9 + t_r12_c2_10;
  assign t_r12_c2_12 = t_r12_c2_11 + p_13_3;
  assign out_12_2 = t_r12_c2_12 >> 4;

  assign t_r12_c3_0 = p_11_3 << 1;
  assign t_r12_c3_1 = p_12_2 << 1;
  assign t_r12_c3_2 = p_12_3 << 2;
  assign t_r12_c3_3 = p_12_4 << 1;
  assign t_r12_c3_4 = p_13_3 << 1;
  assign t_r12_c3_5 = t_r12_c3_0 + p_11_2;
  assign t_r12_c3_6 = t_r12_c3_1 + p_11_4;
  assign t_r12_c3_7 = t_r12_c3_2 + t_r12_c3_3;
  assign t_r12_c3_8 = t_r12_c3_4 + p_13_2;
  assign t_r12_c3_9 = t_r12_c3_5 + t_r12_c3_6;
  assign t_r12_c3_10 = t_r12_c3_7 + t_r12_c3_8;
  assign t_r12_c3_11 = t_r12_c3_9 + t_r12_c3_10;
  assign t_r12_c3_12 = t_r12_c3_11 + p_13_4;
  assign out_12_3 = t_r12_c3_12 >> 4;

  assign t_r12_c4_0 = p_11_4 << 1;
  assign t_r12_c4_1 = p_12_3 << 1;
  assign t_r12_c4_2 = p_12_4 << 2;
  assign t_r12_c4_3 = p_12_5 << 1;
  assign t_r12_c4_4 = p_13_4 << 1;
  assign t_r12_c4_5 = t_r12_c4_0 + p_11_3;
  assign t_r12_c4_6 = t_r12_c4_1 + p_11_5;
  assign t_r12_c4_7 = t_r12_c4_2 + t_r12_c4_3;
  assign t_r12_c4_8 = t_r12_c4_4 + p_13_3;
  assign t_r12_c4_9 = t_r12_c4_5 + t_r12_c4_6;
  assign t_r12_c4_10 = t_r12_c4_7 + t_r12_c4_8;
  assign t_r12_c4_11 = t_r12_c4_9 + t_r12_c4_10;
  assign t_r12_c4_12 = t_r12_c4_11 + p_13_5;
  assign out_12_4 = t_r12_c4_12 >> 4;

  assign t_r12_c5_0 = p_11_5 << 1;
  assign t_r12_c5_1 = p_12_4 << 1;
  assign t_r12_c5_2 = p_12_5 << 2;
  assign t_r12_c5_3 = p_12_6 << 1;
  assign t_r12_c5_4 = p_13_5 << 1;
  assign t_r12_c5_5 = t_r12_c5_0 + p_11_4;
  assign t_r12_c5_6 = t_r12_c5_1 + p_11_6;
  assign t_r12_c5_7 = t_r12_c5_2 + t_r12_c5_3;
  assign t_r12_c5_8 = t_r12_c5_4 + p_13_4;
  assign t_r12_c5_9 = t_r12_c5_5 + t_r12_c5_6;
  assign t_r12_c5_10 = t_r12_c5_7 + t_r12_c5_8;
  assign t_r12_c5_11 = t_r12_c5_9 + t_r12_c5_10;
  assign t_r12_c5_12 = t_r12_c5_11 + p_13_6;
  assign out_12_5 = t_r12_c5_12 >> 4;

  assign t_r12_c6_0 = p_11_6 << 1;
  assign t_r12_c6_1 = p_12_5 << 1;
  assign t_r12_c6_2 = p_12_6 << 2;
  assign t_r12_c6_3 = p_12_7 << 1;
  assign t_r12_c6_4 = p_13_6 << 1;
  assign t_r12_c6_5 = t_r12_c6_0 + p_11_5;
  assign t_r12_c6_6 = t_r12_c6_1 + p_11_7;
  assign t_r12_c6_7 = t_r12_c6_2 + t_r12_c6_3;
  assign t_r12_c6_8 = t_r12_c6_4 + p_13_5;
  assign t_r12_c6_9 = t_r12_c6_5 + t_r12_c6_6;
  assign t_r12_c6_10 = t_r12_c6_7 + t_r12_c6_8;
  assign t_r12_c6_11 = t_r12_c6_9 + t_r12_c6_10;
  assign t_r12_c6_12 = t_r12_c6_11 + p_13_7;
  assign out_12_6 = t_r12_c6_12 >> 4;

  assign t_r12_c7_0 = p_11_7 << 1;
  assign t_r12_c7_1 = p_12_6 << 1;
  assign t_r12_c7_2 = p_12_7 << 2;
  assign t_r12_c7_3 = p_12_8 << 1;
  assign t_r12_c7_4 = p_13_7 << 1;
  assign t_r12_c7_5 = t_r12_c7_0 + p_11_6;
  assign t_r12_c7_6 = t_r12_c7_1 + p_11_8;
  assign t_r12_c7_7 = t_r12_c7_2 + t_r12_c7_3;
  assign t_r12_c7_8 = t_r12_c7_4 + p_13_6;
  assign t_r12_c7_9 = t_r12_c7_5 + t_r12_c7_6;
  assign t_r12_c7_10 = t_r12_c7_7 + t_r12_c7_8;
  assign t_r12_c7_11 = t_r12_c7_9 + t_r12_c7_10;
  assign t_r12_c7_12 = t_r12_c7_11 + p_13_8;
  assign out_12_7 = t_r12_c7_12 >> 4;

  assign t_r12_c8_0 = p_11_8 << 1;
  assign t_r12_c8_1 = p_12_7 << 1;
  assign t_r12_c8_2 = p_12_8 << 2;
  assign t_r12_c8_3 = p_12_9 << 1;
  assign t_r12_c8_4 = p_13_8 << 1;
  assign t_r12_c8_5 = t_r12_c8_0 + p_11_7;
  assign t_r12_c8_6 = t_r12_c8_1 + p_11_9;
  assign t_r12_c8_7 = t_r12_c8_2 + t_r12_c8_3;
  assign t_r12_c8_8 = t_r12_c8_4 + p_13_7;
  assign t_r12_c8_9 = t_r12_c8_5 + t_r12_c8_6;
  assign t_r12_c8_10 = t_r12_c8_7 + t_r12_c8_8;
  assign t_r12_c8_11 = t_r12_c8_9 + t_r12_c8_10;
  assign t_r12_c8_12 = t_r12_c8_11 + p_13_9;
  assign out_12_8 = t_r12_c8_12 >> 4;

  assign t_r12_c9_0 = p_11_9 << 1;
  assign t_r12_c9_1 = p_12_8 << 1;
  assign t_r12_c9_2 = p_12_9 << 2;
  assign t_r12_c9_3 = p_12_10 << 1;
  assign t_r12_c9_4 = p_13_9 << 1;
  assign t_r12_c9_5 = t_r12_c9_0 + p_11_8;
  assign t_r12_c9_6 = t_r12_c9_1 + p_11_10;
  assign t_r12_c9_7 = t_r12_c9_2 + t_r12_c9_3;
  assign t_r12_c9_8 = t_r12_c9_4 + p_13_8;
  assign t_r12_c9_9 = t_r12_c9_5 + t_r12_c9_6;
  assign t_r12_c9_10 = t_r12_c9_7 + t_r12_c9_8;
  assign t_r12_c9_11 = t_r12_c9_9 + t_r12_c9_10;
  assign t_r12_c9_12 = t_r12_c9_11 + p_13_10;
  assign out_12_9 = t_r12_c9_12 >> 4;

  assign t_r12_c10_0 = p_11_10 << 1;
  assign t_r12_c10_1 = p_12_9 << 1;
  assign t_r12_c10_2 = p_12_10 << 2;
  assign t_r12_c10_3 = p_12_11 << 1;
  assign t_r12_c10_4 = p_13_10 << 1;
  assign t_r12_c10_5 = t_r12_c10_0 + p_11_9;
  assign t_r12_c10_6 = t_r12_c10_1 + p_11_11;
  assign t_r12_c10_7 = t_r12_c10_2 + t_r12_c10_3;
  assign t_r12_c10_8 = t_r12_c10_4 + p_13_9;
  assign t_r12_c10_9 = t_r12_c10_5 + t_r12_c10_6;
  assign t_r12_c10_10 = t_r12_c10_7 + t_r12_c10_8;
  assign t_r12_c10_11 = t_r12_c10_9 + t_r12_c10_10;
  assign t_r12_c10_12 = t_r12_c10_11 + p_13_11;
  assign out_12_10 = t_r12_c10_12 >> 4;

  assign t_r12_c11_0 = p_11_11 << 1;
  assign t_r12_c11_1 = p_12_10 << 1;
  assign t_r12_c11_2 = p_12_11 << 2;
  assign t_r12_c11_3 = p_12_12 << 1;
  assign t_r12_c11_4 = p_13_11 << 1;
  assign t_r12_c11_5 = t_r12_c11_0 + p_11_10;
  assign t_r12_c11_6 = t_r12_c11_1 + p_11_12;
  assign t_r12_c11_7 = t_r12_c11_2 + t_r12_c11_3;
  assign t_r12_c11_8 = t_r12_c11_4 + p_13_10;
  assign t_r12_c11_9 = t_r12_c11_5 + t_r12_c11_6;
  assign t_r12_c11_10 = t_r12_c11_7 + t_r12_c11_8;
  assign t_r12_c11_11 = t_r12_c11_9 + t_r12_c11_10;
  assign t_r12_c11_12 = t_r12_c11_11 + p_13_12;
  assign out_12_11 = t_r12_c11_12 >> 4;

  assign t_r12_c12_0 = p_11_12 << 1;
  assign t_r12_c12_1 = p_12_11 << 1;
  assign t_r12_c12_2 = p_12_12 << 2;
  assign t_r12_c12_3 = p_12_13 << 1;
  assign t_r12_c12_4 = p_13_12 << 1;
  assign t_r12_c12_5 = t_r12_c12_0 + p_11_11;
  assign t_r12_c12_6 = t_r12_c12_1 + p_11_13;
  assign t_r12_c12_7 = t_r12_c12_2 + t_r12_c12_3;
  assign t_r12_c12_8 = t_r12_c12_4 + p_13_11;
  assign t_r12_c12_9 = t_r12_c12_5 + t_r12_c12_6;
  assign t_r12_c12_10 = t_r12_c12_7 + t_r12_c12_8;
  assign t_r12_c12_11 = t_r12_c12_9 + t_r12_c12_10;
  assign t_r12_c12_12 = t_r12_c12_11 + p_13_13;
  assign out_12_12 = t_r12_c12_12 >> 4;

  assign t_r12_c13_0 = p_11_13 << 1;
  assign t_r12_c13_1 = p_12_12 << 1;
  assign t_r12_c13_2 = p_12_13 << 2;
  assign t_r12_c13_3 = p_12_14 << 1;
  assign t_r12_c13_4 = p_13_13 << 1;
  assign t_r12_c13_5 = t_r12_c13_0 + p_11_12;
  assign t_r12_c13_6 = t_r12_c13_1 + p_11_14;
  assign t_r12_c13_7 = t_r12_c13_2 + t_r12_c13_3;
  assign t_r12_c13_8 = t_r12_c13_4 + p_13_12;
  assign t_r12_c13_9 = t_r12_c13_5 + t_r12_c13_6;
  assign t_r12_c13_10 = t_r12_c13_7 + t_r12_c13_8;
  assign t_r12_c13_11 = t_r12_c13_9 + t_r12_c13_10;
  assign t_r12_c13_12 = t_r12_c13_11 + p_13_14;
  assign out_12_13 = t_r12_c13_12 >> 4;

  assign t_r12_c14_0 = p_11_14 << 1;
  assign t_r12_c14_1 = p_12_13 << 1;
  assign t_r12_c14_2 = p_12_14 << 2;
  assign t_r12_c14_3 = p_12_15 << 1;
  assign t_r12_c14_4 = p_13_14 << 1;
  assign t_r12_c14_5 = t_r12_c14_0 + p_11_13;
  assign t_r12_c14_6 = t_r12_c14_1 + p_11_15;
  assign t_r12_c14_7 = t_r12_c14_2 + t_r12_c14_3;
  assign t_r12_c14_8 = t_r12_c14_4 + p_13_13;
  assign t_r12_c14_9 = t_r12_c14_5 + t_r12_c14_6;
  assign t_r12_c14_10 = t_r12_c14_7 + t_r12_c14_8;
  assign t_r12_c14_11 = t_r12_c14_9 + t_r12_c14_10;
  assign t_r12_c14_12 = t_r12_c14_11 + p_13_15;
  assign out_12_14 = t_r12_c14_12 >> 4;

  assign t_r12_c15_0 = p_11_15 << 1;
  assign t_r12_c15_1 = p_12_14 << 1;
  assign t_r12_c15_2 = p_12_15 << 2;
  assign t_r12_c15_3 = p_12_16 << 1;
  assign t_r12_c15_4 = p_13_15 << 1;
  assign t_r12_c15_5 = t_r12_c15_0 + p_11_14;
  assign t_r12_c15_6 = t_r12_c15_1 + p_11_16;
  assign t_r12_c15_7 = t_r12_c15_2 + t_r12_c15_3;
  assign t_r12_c15_8 = t_r12_c15_4 + p_13_14;
  assign t_r12_c15_9 = t_r12_c15_5 + t_r12_c15_6;
  assign t_r12_c15_10 = t_r12_c15_7 + t_r12_c15_8;
  assign t_r12_c15_11 = t_r12_c15_9 + t_r12_c15_10;
  assign t_r12_c15_12 = t_r12_c15_11 + p_13_16;
  assign out_12_15 = t_r12_c15_12 >> 4;

  assign t_r12_c16_0 = p_11_16 << 1;
  assign t_r12_c16_1 = p_12_15 << 1;
  assign t_r12_c16_2 = p_12_16 << 2;
  assign t_r12_c16_3 = p_12_17 << 1;
  assign t_r12_c16_4 = p_13_16 << 1;
  assign t_r12_c16_5 = t_r12_c16_0 + p_11_15;
  assign t_r12_c16_6 = t_r12_c16_1 + p_11_17;
  assign t_r12_c16_7 = t_r12_c16_2 + t_r12_c16_3;
  assign t_r12_c16_8 = t_r12_c16_4 + p_13_15;
  assign t_r12_c16_9 = t_r12_c16_5 + t_r12_c16_6;
  assign t_r12_c16_10 = t_r12_c16_7 + t_r12_c16_8;
  assign t_r12_c16_11 = t_r12_c16_9 + t_r12_c16_10;
  assign t_r12_c16_12 = t_r12_c16_11 + p_13_17;
  assign out_12_16 = t_r12_c16_12 >> 4;

  assign t_r12_c17_0 = p_11_17 << 1;
  assign t_r12_c17_1 = p_12_16 << 1;
  assign t_r12_c17_2 = p_12_17 << 2;
  assign t_r12_c17_3 = p_12_18 << 1;
  assign t_r12_c17_4 = p_13_17 << 1;
  assign t_r12_c17_5 = t_r12_c17_0 + p_11_16;
  assign t_r12_c17_6 = t_r12_c17_1 + p_11_18;
  assign t_r12_c17_7 = t_r12_c17_2 + t_r12_c17_3;
  assign t_r12_c17_8 = t_r12_c17_4 + p_13_16;
  assign t_r12_c17_9 = t_r12_c17_5 + t_r12_c17_6;
  assign t_r12_c17_10 = t_r12_c17_7 + t_r12_c17_8;
  assign t_r12_c17_11 = t_r12_c17_9 + t_r12_c17_10;
  assign t_r12_c17_12 = t_r12_c17_11 + p_13_18;
  assign out_12_17 = t_r12_c17_12 >> 4;

  assign t_r12_c18_0 = p_11_18 << 1;
  assign t_r12_c18_1 = p_12_17 << 1;
  assign t_r12_c18_2 = p_12_18 << 2;
  assign t_r12_c18_3 = p_12_19 << 1;
  assign t_r12_c18_4 = p_13_18 << 1;
  assign t_r12_c18_5 = t_r12_c18_0 + p_11_17;
  assign t_r12_c18_6 = t_r12_c18_1 + p_11_19;
  assign t_r12_c18_7 = t_r12_c18_2 + t_r12_c18_3;
  assign t_r12_c18_8 = t_r12_c18_4 + p_13_17;
  assign t_r12_c18_9 = t_r12_c18_5 + t_r12_c18_6;
  assign t_r12_c18_10 = t_r12_c18_7 + t_r12_c18_8;
  assign t_r12_c18_11 = t_r12_c18_9 + t_r12_c18_10;
  assign t_r12_c18_12 = t_r12_c18_11 + p_13_19;
  assign out_12_18 = t_r12_c18_12 >> 4;

  assign t_r12_c19_0 = p_11_19 << 1;
  assign t_r12_c19_1 = p_12_18 << 1;
  assign t_r12_c19_2 = p_12_19 << 2;
  assign t_r12_c19_3 = p_12_20 << 1;
  assign t_r12_c19_4 = p_13_19 << 1;
  assign t_r12_c19_5 = t_r12_c19_0 + p_11_18;
  assign t_r12_c19_6 = t_r12_c19_1 + p_11_20;
  assign t_r12_c19_7 = t_r12_c19_2 + t_r12_c19_3;
  assign t_r12_c19_8 = t_r12_c19_4 + p_13_18;
  assign t_r12_c19_9 = t_r12_c19_5 + t_r12_c19_6;
  assign t_r12_c19_10 = t_r12_c19_7 + t_r12_c19_8;
  assign t_r12_c19_11 = t_r12_c19_9 + t_r12_c19_10;
  assign t_r12_c19_12 = t_r12_c19_11 + p_13_20;
  assign out_12_19 = t_r12_c19_12 >> 4;

  assign t_r12_c20_0 = p_11_20 << 1;
  assign t_r12_c20_1 = p_12_19 << 1;
  assign t_r12_c20_2 = p_12_20 << 2;
  assign t_r12_c20_3 = p_12_21 << 1;
  assign t_r12_c20_4 = p_13_20 << 1;
  assign t_r12_c20_5 = t_r12_c20_0 + p_11_19;
  assign t_r12_c20_6 = t_r12_c20_1 + p_11_21;
  assign t_r12_c20_7 = t_r12_c20_2 + t_r12_c20_3;
  assign t_r12_c20_8 = t_r12_c20_4 + p_13_19;
  assign t_r12_c20_9 = t_r12_c20_5 + t_r12_c20_6;
  assign t_r12_c20_10 = t_r12_c20_7 + t_r12_c20_8;
  assign t_r12_c20_11 = t_r12_c20_9 + t_r12_c20_10;
  assign t_r12_c20_12 = t_r12_c20_11 + p_13_21;
  assign out_12_20 = t_r12_c20_12 >> 4;

  assign t_r12_c21_0 = p_11_21 << 1;
  assign t_r12_c21_1 = p_12_20 << 1;
  assign t_r12_c21_2 = p_12_21 << 2;
  assign t_r12_c21_3 = p_12_22 << 1;
  assign t_r12_c21_4 = p_13_21 << 1;
  assign t_r12_c21_5 = t_r12_c21_0 + p_11_20;
  assign t_r12_c21_6 = t_r12_c21_1 + p_11_22;
  assign t_r12_c21_7 = t_r12_c21_2 + t_r12_c21_3;
  assign t_r12_c21_8 = t_r12_c21_4 + p_13_20;
  assign t_r12_c21_9 = t_r12_c21_5 + t_r12_c21_6;
  assign t_r12_c21_10 = t_r12_c21_7 + t_r12_c21_8;
  assign t_r12_c21_11 = t_r12_c21_9 + t_r12_c21_10;
  assign t_r12_c21_12 = t_r12_c21_11 + p_13_22;
  assign out_12_21 = t_r12_c21_12 >> 4;

  assign t_r12_c22_0 = p_11_22 << 1;
  assign t_r12_c22_1 = p_12_21 << 1;
  assign t_r12_c22_2 = p_12_22 << 2;
  assign t_r12_c22_3 = p_12_23 << 1;
  assign t_r12_c22_4 = p_13_22 << 1;
  assign t_r12_c22_5 = t_r12_c22_0 + p_11_21;
  assign t_r12_c22_6 = t_r12_c22_1 + p_11_23;
  assign t_r12_c22_7 = t_r12_c22_2 + t_r12_c22_3;
  assign t_r12_c22_8 = t_r12_c22_4 + p_13_21;
  assign t_r12_c22_9 = t_r12_c22_5 + t_r12_c22_6;
  assign t_r12_c22_10 = t_r12_c22_7 + t_r12_c22_8;
  assign t_r12_c22_11 = t_r12_c22_9 + t_r12_c22_10;
  assign t_r12_c22_12 = t_r12_c22_11 + p_13_23;
  assign out_12_22 = t_r12_c22_12 >> 4;

  assign t_r12_c23_0 = p_11_23 << 1;
  assign t_r12_c23_1 = p_12_22 << 1;
  assign t_r12_c23_2 = p_12_23 << 2;
  assign t_r12_c23_3 = p_12_24 << 1;
  assign t_r12_c23_4 = p_13_23 << 1;
  assign t_r12_c23_5 = t_r12_c23_0 + p_11_22;
  assign t_r12_c23_6 = t_r12_c23_1 + p_11_24;
  assign t_r12_c23_7 = t_r12_c23_2 + t_r12_c23_3;
  assign t_r12_c23_8 = t_r12_c23_4 + p_13_22;
  assign t_r12_c23_9 = t_r12_c23_5 + t_r12_c23_6;
  assign t_r12_c23_10 = t_r12_c23_7 + t_r12_c23_8;
  assign t_r12_c23_11 = t_r12_c23_9 + t_r12_c23_10;
  assign t_r12_c23_12 = t_r12_c23_11 + p_13_24;
  assign out_12_23 = t_r12_c23_12 >> 4;

  assign t_r12_c24_0 = p_11_24 << 1;
  assign t_r12_c24_1 = p_12_23 << 1;
  assign t_r12_c24_2 = p_12_24 << 2;
  assign t_r12_c24_3 = p_12_25 << 1;
  assign t_r12_c24_4 = p_13_24 << 1;
  assign t_r12_c24_5 = t_r12_c24_0 + p_11_23;
  assign t_r12_c24_6 = t_r12_c24_1 + p_11_25;
  assign t_r12_c24_7 = t_r12_c24_2 + t_r12_c24_3;
  assign t_r12_c24_8 = t_r12_c24_4 + p_13_23;
  assign t_r12_c24_9 = t_r12_c24_5 + t_r12_c24_6;
  assign t_r12_c24_10 = t_r12_c24_7 + t_r12_c24_8;
  assign t_r12_c24_11 = t_r12_c24_9 + t_r12_c24_10;
  assign t_r12_c24_12 = t_r12_c24_11 + p_13_25;
  assign out_12_24 = t_r12_c24_12 >> 4;

  assign t_r12_c25_0 = p_11_25 << 1;
  assign t_r12_c25_1 = p_12_24 << 1;
  assign t_r12_c25_2 = p_12_25 << 2;
  assign t_r12_c25_3 = p_12_26 << 1;
  assign t_r12_c25_4 = p_13_25 << 1;
  assign t_r12_c25_5 = t_r12_c25_0 + p_11_24;
  assign t_r12_c25_6 = t_r12_c25_1 + p_11_26;
  assign t_r12_c25_7 = t_r12_c25_2 + t_r12_c25_3;
  assign t_r12_c25_8 = t_r12_c25_4 + p_13_24;
  assign t_r12_c25_9 = t_r12_c25_5 + t_r12_c25_6;
  assign t_r12_c25_10 = t_r12_c25_7 + t_r12_c25_8;
  assign t_r12_c25_11 = t_r12_c25_9 + t_r12_c25_10;
  assign t_r12_c25_12 = t_r12_c25_11 + p_13_26;
  assign out_12_25 = t_r12_c25_12 >> 4;

  assign t_r12_c26_0 = p_11_26 << 1;
  assign t_r12_c26_1 = p_12_25 << 1;
  assign t_r12_c26_2 = p_12_26 << 2;
  assign t_r12_c26_3 = p_12_27 << 1;
  assign t_r12_c26_4 = p_13_26 << 1;
  assign t_r12_c26_5 = t_r12_c26_0 + p_11_25;
  assign t_r12_c26_6 = t_r12_c26_1 + p_11_27;
  assign t_r12_c26_7 = t_r12_c26_2 + t_r12_c26_3;
  assign t_r12_c26_8 = t_r12_c26_4 + p_13_25;
  assign t_r12_c26_9 = t_r12_c26_5 + t_r12_c26_6;
  assign t_r12_c26_10 = t_r12_c26_7 + t_r12_c26_8;
  assign t_r12_c26_11 = t_r12_c26_9 + t_r12_c26_10;
  assign t_r12_c26_12 = t_r12_c26_11 + p_13_27;
  assign out_12_26 = t_r12_c26_12 >> 4;

  assign t_r12_c27_0 = p_11_27 << 1;
  assign t_r12_c27_1 = p_12_26 << 1;
  assign t_r12_c27_2 = p_12_27 << 2;
  assign t_r12_c27_3 = p_12_28 << 1;
  assign t_r12_c27_4 = p_13_27 << 1;
  assign t_r12_c27_5 = t_r12_c27_0 + p_11_26;
  assign t_r12_c27_6 = t_r12_c27_1 + p_11_28;
  assign t_r12_c27_7 = t_r12_c27_2 + t_r12_c27_3;
  assign t_r12_c27_8 = t_r12_c27_4 + p_13_26;
  assign t_r12_c27_9 = t_r12_c27_5 + t_r12_c27_6;
  assign t_r12_c27_10 = t_r12_c27_7 + t_r12_c27_8;
  assign t_r12_c27_11 = t_r12_c27_9 + t_r12_c27_10;
  assign t_r12_c27_12 = t_r12_c27_11 + p_13_28;
  assign out_12_27 = t_r12_c27_12 >> 4;

  assign t_r12_c28_0 = p_11_28 << 1;
  assign t_r12_c28_1 = p_12_27 << 1;
  assign t_r12_c28_2 = p_12_28 << 2;
  assign t_r12_c28_3 = p_12_29 << 1;
  assign t_r12_c28_4 = p_13_28 << 1;
  assign t_r12_c28_5 = t_r12_c28_0 + p_11_27;
  assign t_r12_c28_6 = t_r12_c28_1 + p_11_29;
  assign t_r12_c28_7 = t_r12_c28_2 + t_r12_c28_3;
  assign t_r12_c28_8 = t_r12_c28_4 + p_13_27;
  assign t_r12_c28_9 = t_r12_c28_5 + t_r12_c28_6;
  assign t_r12_c28_10 = t_r12_c28_7 + t_r12_c28_8;
  assign t_r12_c28_11 = t_r12_c28_9 + t_r12_c28_10;
  assign t_r12_c28_12 = t_r12_c28_11 + p_13_29;
  assign out_12_28 = t_r12_c28_12 >> 4;

  assign t_r12_c29_0 = p_11_29 << 1;
  assign t_r12_c29_1 = p_12_28 << 1;
  assign t_r12_c29_2 = p_12_29 << 2;
  assign t_r12_c29_3 = p_12_30 << 1;
  assign t_r12_c29_4 = p_13_29 << 1;
  assign t_r12_c29_5 = t_r12_c29_0 + p_11_28;
  assign t_r12_c29_6 = t_r12_c29_1 + p_11_30;
  assign t_r12_c29_7 = t_r12_c29_2 + t_r12_c29_3;
  assign t_r12_c29_8 = t_r12_c29_4 + p_13_28;
  assign t_r12_c29_9 = t_r12_c29_5 + t_r12_c29_6;
  assign t_r12_c29_10 = t_r12_c29_7 + t_r12_c29_8;
  assign t_r12_c29_11 = t_r12_c29_9 + t_r12_c29_10;
  assign t_r12_c29_12 = t_r12_c29_11 + p_13_30;
  assign out_12_29 = t_r12_c29_12 >> 4;

  assign t_r12_c30_0 = p_11_30 << 1;
  assign t_r12_c30_1 = p_12_29 << 1;
  assign t_r12_c30_2 = p_12_30 << 2;
  assign t_r12_c30_3 = p_12_31 << 1;
  assign t_r12_c30_4 = p_13_30 << 1;
  assign t_r12_c30_5 = t_r12_c30_0 + p_11_29;
  assign t_r12_c30_6 = t_r12_c30_1 + p_11_31;
  assign t_r12_c30_7 = t_r12_c30_2 + t_r12_c30_3;
  assign t_r12_c30_8 = t_r12_c30_4 + p_13_29;
  assign t_r12_c30_9 = t_r12_c30_5 + t_r12_c30_6;
  assign t_r12_c30_10 = t_r12_c30_7 + t_r12_c30_8;
  assign t_r12_c30_11 = t_r12_c30_9 + t_r12_c30_10;
  assign t_r12_c30_12 = t_r12_c30_11 + p_13_31;
  assign out_12_30 = t_r12_c30_12 >> 4;

  assign t_r12_c31_0 = p_11_31 << 1;
  assign t_r12_c31_1 = p_12_30 << 1;
  assign t_r12_c31_2 = p_12_31 << 2;
  assign t_r12_c31_3 = p_12_32 << 1;
  assign t_r12_c31_4 = p_13_31 << 1;
  assign t_r12_c31_5 = t_r12_c31_0 + p_11_30;
  assign t_r12_c31_6 = t_r12_c31_1 + p_11_32;
  assign t_r12_c31_7 = t_r12_c31_2 + t_r12_c31_3;
  assign t_r12_c31_8 = t_r12_c31_4 + p_13_30;
  assign t_r12_c31_9 = t_r12_c31_5 + t_r12_c31_6;
  assign t_r12_c31_10 = t_r12_c31_7 + t_r12_c31_8;
  assign t_r12_c31_11 = t_r12_c31_9 + t_r12_c31_10;
  assign t_r12_c31_12 = t_r12_c31_11 + p_13_32;
  assign out_12_31 = t_r12_c31_12 >> 4;

  assign t_r12_c32_0 = p_11_32 << 1;
  assign t_r12_c32_1 = p_12_31 << 1;
  assign t_r12_c32_2 = p_12_32 << 2;
  assign t_r12_c32_3 = p_12_33 << 1;
  assign t_r12_c32_4 = p_13_32 << 1;
  assign t_r12_c32_5 = t_r12_c32_0 + p_11_31;
  assign t_r12_c32_6 = t_r12_c32_1 + p_11_33;
  assign t_r12_c32_7 = t_r12_c32_2 + t_r12_c32_3;
  assign t_r12_c32_8 = t_r12_c32_4 + p_13_31;
  assign t_r12_c32_9 = t_r12_c32_5 + t_r12_c32_6;
  assign t_r12_c32_10 = t_r12_c32_7 + t_r12_c32_8;
  assign t_r12_c32_11 = t_r12_c32_9 + t_r12_c32_10;
  assign t_r12_c32_12 = t_r12_c32_11 + p_13_33;
  assign out_12_32 = t_r12_c32_12 >> 4;

  assign t_r12_c33_0 = p_11_33 << 1;
  assign t_r12_c33_1 = p_12_32 << 1;
  assign t_r12_c33_2 = p_12_33 << 2;
  assign t_r12_c33_3 = p_12_34 << 1;
  assign t_r12_c33_4 = p_13_33 << 1;
  assign t_r12_c33_5 = t_r12_c33_0 + p_11_32;
  assign t_r12_c33_6 = t_r12_c33_1 + p_11_34;
  assign t_r12_c33_7 = t_r12_c33_2 + t_r12_c33_3;
  assign t_r12_c33_8 = t_r12_c33_4 + p_13_32;
  assign t_r12_c33_9 = t_r12_c33_5 + t_r12_c33_6;
  assign t_r12_c33_10 = t_r12_c33_7 + t_r12_c33_8;
  assign t_r12_c33_11 = t_r12_c33_9 + t_r12_c33_10;
  assign t_r12_c33_12 = t_r12_c33_11 + p_13_34;
  assign out_12_33 = t_r12_c33_12 >> 4;

  assign t_r12_c34_0 = p_11_34 << 1;
  assign t_r12_c34_1 = p_12_33 << 1;
  assign t_r12_c34_2 = p_12_34 << 2;
  assign t_r12_c34_3 = p_12_35 << 1;
  assign t_r12_c34_4 = p_13_34 << 1;
  assign t_r12_c34_5 = t_r12_c34_0 + p_11_33;
  assign t_r12_c34_6 = t_r12_c34_1 + p_11_35;
  assign t_r12_c34_7 = t_r12_c34_2 + t_r12_c34_3;
  assign t_r12_c34_8 = t_r12_c34_4 + p_13_33;
  assign t_r12_c34_9 = t_r12_c34_5 + t_r12_c34_6;
  assign t_r12_c34_10 = t_r12_c34_7 + t_r12_c34_8;
  assign t_r12_c34_11 = t_r12_c34_9 + t_r12_c34_10;
  assign t_r12_c34_12 = t_r12_c34_11 + p_13_35;
  assign out_12_34 = t_r12_c34_12 >> 4;

  assign t_r12_c35_0 = p_11_35 << 1;
  assign t_r12_c35_1 = p_12_34 << 1;
  assign t_r12_c35_2 = p_12_35 << 2;
  assign t_r12_c35_3 = p_12_36 << 1;
  assign t_r12_c35_4 = p_13_35 << 1;
  assign t_r12_c35_5 = t_r12_c35_0 + p_11_34;
  assign t_r12_c35_6 = t_r12_c35_1 + p_11_36;
  assign t_r12_c35_7 = t_r12_c35_2 + t_r12_c35_3;
  assign t_r12_c35_8 = t_r12_c35_4 + p_13_34;
  assign t_r12_c35_9 = t_r12_c35_5 + t_r12_c35_6;
  assign t_r12_c35_10 = t_r12_c35_7 + t_r12_c35_8;
  assign t_r12_c35_11 = t_r12_c35_9 + t_r12_c35_10;
  assign t_r12_c35_12 = t_r12_c35_11 + p_13_36;
  assign out_12_35 = t_r12_c35_12 >> 4;

  assign t_r12_c36_0 = p_11_36 << 1;
  assign t_r12_c36_1 = p_12_35 << 1;
  assign t_r12_c36_2 = p_12_36 << 2;
  assign t_r12_c36_3 = p_12_37 << 1;
  assign t_r12_c36_4 = p_13_36 << 1;
  assign t_r12_c36_5 = t_r12_c36_0 + p_11_35;
  assign t_r12_c36_6 = t_r12_c36_1 + p_11_37;
  assign t_r12_c36_7 = t_r12_c36_2 + t_r12_c36_3;
  assign t_r12_c36_8 = t_r12_c36_4 + p_13_35;
  assign t_r12_c36_9 = t_r12_c36_5 + t_r12_c36_6;
  assign t_r12_c36_10 = t_r12_c36_7 + t_r12_c36_8;
  assign t_r12_c36_11 = t_r12_c36_9 + t_r12_c36_10;
  assign t_r12_c36_12 = t_r12_c36_11 + p_13_37;
  assign out_12_36 = t_r12_c36_12 >> 4;

  assign t_r12_c37_0 = p_11_37 << 1;
  assign t_r12_c37_1 = p_12_36 << 1;
  assign t_r12_c37_2 = p_12_37 << 2;
  assign t_r12_c37_3 = p_12_38 << 1;
  assign t_r12_c37_4 = p_13_37 << 1;
  assign t_r12_c37_5 = t_r12_c37_0 + p_11_36;
  assign t_r12_c37_6 = t_r12_c37_1 + p_11_38;
  assign t_r12_c37_7 = t_r12_c37_2 + t_r12_c37_3;
  assign t_r12_c37_8 = t_r12_c37_4 + p_13_36;
  assign t_r12_c37_9 = t_r12_c37_5 + t_r12_c37_6;
  assign t_r12_c37_10 = t_r12_c37_7 + t_r12_c37_8;
  assign t_r12_c37_11 = t_r12_c37_9 + t_r12_c37_10;
  assign t_r12_c37_12 = t_r12_c37_11 + p_13_38;
  assign out_12_37 = t_r12_c37_12 >> 4;

  assign t_r12_c38_0 = p_11_38 << 1;
  assign t_r12_c38_1 = p_12_37 << 1;
  assign t_r12_c38_2 = p_12_38 << 2;
  assign t_r12_c38_3 = p_12_39 << 1;
  assign t_r12_c38_4 = p_13_38 << 1;
  assign t_r12_c38_5 = t_r12_c38_0 + p_11_37;
  assign t_r12_c38_6 = t_r12_c38_1 + p_11_39;
  assign t_r12_c38_7 = t_r12_c38_2 + t_r12_c38_3;
  assign t_r12_c38_8 = t_r12_c38_4 + p_13_37;
  assign t_r12_c38_9 = t_r12_c38_5 + t_r12_c38_6;
  assign t_r12_c38_10 = t_r12_c38_7 + t_r12_c38_8;
  assign t_r12_c38_11 = t_r12_c38_9 + t_r12_c38_10;
  assign t_r12_c38_12 = t_r12_c38_11 + p_13_39;
  assign out_12_38 = t_r12_c38_12 >> 4;

  assign t_r12_c39_0 = p_11_39 << 1;
  assign t_r12_c39_1 = p_12_38 << 1;
  assign t_r12_c39_2 = p_12_39 << 2;
  assign t_r12_c39_3 = p_12_40 << 1;
  assign t_r12_c39_4 = p_13_39 << 1;
  assign t_r12_c39_5 = t_r12_c39_0 + p_11_38;
  assign t_r12_c39_6 = t_r12_c39_1 + p_11_40;
  assign t_r12_c39_7 = t_r12_c39_2 + t_r12_c39_3;
  assign t_r12_c39_8 = t_r12_c39_4 + p_13_38;
  assign t_r12_c39_9 = t_r12_c39_5 + t_r12_c39_6;
  assign t_r12_c39_10 = t_r12_c39_7 + t_r12_c39_8;
  assign t_r12_c39_11 = t_r12_c39_9 + t_r12_c39_10;
  assign t_r12_c39_12 = t_r12_c39_11 + p_13_40;
  assign out_12_39 = t_r12_c39_12 >> 4;

  assign t_r12_c40_0 = p_11_40 << 1;
  assign t_r12_c40_1 = p_12_39 << 1;
  assign t_r12_c40_2 = p_12_40 << 2;
  assign t_r12_c40_3 = p_12_41 << 1;
  assign t_r12_c40_4 = p_13_40 << 1;
  assign t_r12_c40_5 = t_r12_c40_0 + p_11_39;
  assign t_r12_c40_6 = t_r12_c40_1 + p_11_41;
  assign t_r12_c40_7 = t_r12_c40_2 + t_r12_c40_3;
  assign t_r12_c40_8 = t_r12_c40_4 + p_13_39;
  assign t_r12_c40_9 = t_r12_c40_5 + t_r12_c40_6;
  assign t_r12_c40_10 = t_r12_c40_7 + t_r12_c40_8;
  assign t_r12_c40_11 = t_r12_c40_9 + t_r12_c40_10;
  assign t_r12_c40_12 = t_r12_c40_11 + p_13_41;
  assign out_12_40 = t_r12_c40_12 >> 4;

  assign t_r12_c41_0 = p_11_41 << 1;
  assign t_r12_c41_1 = p_12_40 << 1;
  assign t_r12_c41_2 = p_12_41 << 2;
  assign t_r12_c41_3 = p_12_42 << 1;
  assign t_r12_c41_4 = p_13_41 << 1;
  assign t_r12_c41_5 = t_r12_c41_0 + p_11_40;
  assign t_r12_c41_6 = t_r12_c41_1 + p_11_42;
  assign t_r12_c41_7 = t_r12_c41_2 + t_r12_c41_3;
  assign t_r12_c41_8 = t_r12_c41_4 + p_13_40;
  assign t_r12_c41_9 = t_r12_c41_5 + t_r12_c41_6;
  assign t_r12_c41_10 = t_r12_c41_7 + t_r12_c41_8;
  assign t_r12_c41_11 = t_r12_c41_9 + t_r12_c41_10;
  assign t_r12_c41_12 = t_r12_c41_11 + p_13_42;
  assign out_12_41 = t_r12_c41_12 >> 4;

  assign t_r12_c42_0 = p_11_42 << 1;
  assign t_r12_c42_1 = p_12_41 << 1;
  assign t_r12_c42_2 = p_12_42 << 2;
  assign t_r12_c42_3 = p_12_43 << 1;
  assign t_r12_c42_4 = p_13_42 << 1;
  assign t_r12_c42_5 = t_r12_c42_0 + p_11_41;
  assign t_r12_c42_6 = t_r12_c42_1 + p_11_43;
  assign t_r12_c42_7 = t_r12_c42_2 + t_r12_c42_3;
  assign t_r12_c42_8 = t_r12_c42_4 + p_13_41;
  assign t_r12_c42_9 = t_r12_c42_5 + t_r12_c42_6;
  assign t_r12_c42_10 = t_r12_c42_7 + t_r12_c42_8;
  assign t_r12_c42_11 = t_r12_c42_9 + t_r12_c42_10;
  assign t_r12_c42_12 = t_r12_c42_11 + p_13_43;
  assign out_12_42 = t_r12_c42_12 >> 4;

  assign t_r12_c43_0 = p_11_43 << 1;
  assign t_r12_c43_1 = p_12_42 << 1;
  assign t_r12_c43_2 = p_12_43 << 2;
  assign t_r12_c43_3 = p_12_44 << 1;
  assign t_r12_c43_4 = p_13_43 << 1;
  assign t_r12_c43_5 = t_r12_c43_0 + p_11_42;
  assign t_r12_c43_6 = t_r12_c43_1 + p_11_44;
  assign t_r12_c43_7 = t_r12_c43_2 + t_r12_c43_3;
  assign t_r12_c43_8 = t_r12_c43_4 + p_13_42;
  assign t_r12_c43_9 = t_r12_c43_5 + t_r12_c43_6;
  assign t_r12_c43_10 = t_r12_c43_7 + t_r12_c43_8;
  assign t_r12_c43_11 = t_r12_c43_9 + t_r12_c43_10;
  assign t_r12_c43_12 = t_r12_c43_11 + p_13_44;
  assign out_12_43 = t_r12_c43_12 >> 4;

  assign t_r12_c44_0 = p_11_44 << 1;
  assign t_r12_c44_1 = p_12_43 << 1;
  assign t_r12_c44_2 = p_12_44 << 2;
  assign t_r12_c44_3 = p_12_45 << 1;
  assign t_r12_c44_4 = p_13_44 << 1;
  assign t_r12_c44_5 = t_r12_c44_0 + p_11_43;
  assign t_r12_c44_6 = t_r12_c44_1 + p_11_45;
  assign t_r12_c44_7 = t_r12_c44_2 + t_r12_c44_3;
  assign t_r12_c44_8 = t_r12_c44_4 + p_13_43;
  assign t_r12_c44_9 = t_r12_c44_5 + t_r12_c44_6;
  assign t_r12_c44_10 = t_r12_c44_7 + t_r12_c44_8;
  assign t_r12_c44_11 = t_r12_c44_9 + t_r12_c44_10;
  assign t_r12_c44_12 = t_r12_c44_11 + p_13_45;
  assign out_12_44 = t_r12_c44_12 >> 4;

  assign t_r12_c45_0 = p_11_45 << 1;
  assign t_r12_c45_1 = p_12_44 << 1;
  assign t_r12_c45_2 = p_12_45 << 2;
  assign t_r12_c45_3 = p_12_46 << 1;
  assign t_r12_c45_4 = p_13_45 << 1;
  assign t_r12_c45_5 = t_r12_c45_0 + p_11_44;
  assign t_r12_c45_6 = t_r12_c45_1 + p_11_46;
  assign t_r12_c45_7 = t_r12_c45_2 + t_r12_c45_3;
  assign t_r12_c45_8 = t_r12_c45_4 + p_13_44;
  assign t_r12_c45_9 = t_r12_c45_5 + t_r12_c45_6;
  assign t_r12_c45_10 = t_r12_c45_7 + t_r12_c45_8;
  assign t_r12_c45_11 = t_r12_c45_9 + t_r12_c45_10;
  assign t_r12_c45_12 = t_r12_c45_11 + p_13_46;
  assign out_12_45 = t_r12_c45_12 >> 4;

  assign t_r12_c46_0 = p_11_46 << 1;
  assign t_r12_c46_1 = p_12_45 << 1;
  assign t_r12_c46_2 = p_12_46 << 2;
  assign t_r12_c46_3 = p_12_47 << 1;
  assign t_r12_c46_4 = p_13_46 << 1;
  assign t_r12_c46_5 = t_r12_c46_0 + p_11_45;
  assign t_r12_c46_6 = t_r12_c46_1 + p_11_47;
  assign t_r12_c46_7 = t_r12_c46_2 + t_r12_c46_3;
  assign t_r12_c46_8 = t_r12_c46_4 + p_13_45;
  assign t_r12_c46_9 = t_r12_c46_5 + t_r12_c46_6;
  assign t_r12_c46_10 = t_r12_c46_7 + t_r12_c46_8;
  assign t_r12_c46_11 = t_r12_c46_9 + t_r12_c46_10;
  assign t_r12_c46_12 = t_r12_c46_11 + p_13_47;
  assign out_12_46 = t_r12_c46_12 >> 4;

  assign t_r12_c47_0 = p_11_47 << 1;
  assign t_r12_c47_1 = p_12_46 << 1;
  assign t_r12_c47_2 = p_12_47 << 2;
  assign t_r12_c47_3 = p_12_48 << 1;
  assign t_r12_c47_4 = p_13_47 << 1;
  assign t_r12_c47_5 = t_r12_c47_0 + p_11_46;
  assign t_r12_c47_6 = t_r12_c47_1 + p_11_48;
  assign t_r12_c47_7 = t_r12_c47_2 + t_r12_c47_3;
  assign t_r12_c47_8 = t_r12_c47_4 + p_13_46;
  assign t_r12_c47_9 = t_r12_c47_5 + t_r12_c47_6;
  assign t_r12_c47_10 = t_r12_c47_7 + t_r12_c47_8;
  assign t_r12_c47_11 = t_r12_c47_9 + t_r12_c47_10;
  assign t_r12_c47_12 = t_r12_c47_11 + p_13_48;
  assign out_12_47 = t_r12_c47_12 >> 4;

  assign t_r12_c48_0 = p_11_48 << 1;
  assign t_r12_c48_1 = p_12_47 << 1;
  assign t_r12_c48_2 = p_12_48 << 2;
  assign t_r12_c48_3 = p_12_49 << 1;
  assign t_r12_c48_4 = p_13_48 << 1;
  assign t_r12_c48_5 = t_r12_c48_0 + p_11_47;
  assign t_r12_c48_6 = t_r12_c48_1 + p_11_49;
  assign t_r12_c48_7 = t_r12_c48_2 + t_r12_c48_3;
  assign t_r12_c48_8 = t_r12_c48_4 + p_13_47;
  assign t_r12_c48_9 = t_r12_c48_5 + t_r12_c48_6;
  assign t_r12_c48_10 = t_r12_c48_7 + t_r12_c48_8;
  assign t_r12_c48_11 = t_r12_c48_9 + t_r12_c48_10;
  assign t_r12_c48_12 = t_r12_c48_11 + p_13_49;
  assign out_12_48 = t_r12_c48_12 >> 4;

  assign t_r12_c49_0 = p_11_49 << 1;
  assign t_r12_c49_1 = p_12_48 << 1;
  assign t_r12_c49_2 = p_12_49 << 2;
  assign t_r12_c49_3 = p_12_50 << 1;
  assign t_r12_c49_4 = p_13_49 << 1;
  assign t_r12_c49_5 = t_r12_c49_0 + p_11_48;
  assign t_r12_c49_6 = t_r12_c49_1 + p_11_50;
  assign t_r12_c49_7 = t_r12_c49_2 + t_r12_c49_3;
  assign t_r12_c49_8 = t_r12_c49_4 + p_13_48;
  assign t_r12_c49_9 = t_r12_c49_5 + t_r12_c49_6;
  assign t_r12_c49_10 = t_r12_c49_7 + t_r12_c49_8;
  assign t_r12_c49_11 = t_r12_c49_9 + t_r12_c49_10;
  assign t_r12_c49_12 = t_r12_c49_11 + p_13_50;
  assign out_12_49 = t_r12_c49_12 >> 4;

  assign t_r12_c50_0 = p_11_50 << 1;
  assign t_r12_c50_1 = p_12_49 << 1;
  assign t_r12_c50_2 = p_12_50 << 2;
  assign t_r12_c50_3 = p_12_51 << 1;
  assign t_r12_c50_4 = p_13_50 << 1;
  assign t_r12_c50_5 = t_r12_c50_0 + p_11_49;
  assign t_r12_c50_6 = t_r12_c50_1 + p_11_51;
  assign t_r12_c50_7 = t_r12_c50_2 + t_r12_c50_3;
  assign t_r12_c50_8 = t_r12_c50_4 + p_13_49;
  assign t_r12_c50_9 = t_r12_c50_5 + t_r12_c50_6;
  assign t_r12_c50_10 = t_r12_c50_7 + t_r12_c50_8;
  assign t_r12_c50_11 = t_r12_c50_9 + t_r12_c50_10;
  assign t_r12_c50_12 = t_r12_c50_11 + p_13_51;
  assign out_12_50 = t_r12_c50_12 >> 4;

  assign t_r12_c51_0 = p_11_51 << 1;
  assign t_r12_c51_1 = p_12_50 << 1;
  assign t_r12_c51_2 = p_12_51 << 2;
  assign t_r12_c51_3 = p_12_52 << 1;
  assign t_r12_c51_4 = p_13_51 << 1;
  assign t_r12_c51_5 = t_r12_c51_0 + p_11_50;
  assign t_r12_c51_6 = t_r12_c51_1 + p_11_52;
  assign t_r12_c51_7 = t_r12_c51_2 + t_r12_c51_3;
  assign t_r12_c51_8 = t_r12_c51_4 + p_13_50;
  assign t_r12_c51_9 = t_r12_c51_5 + t_r12_c51_6;
  assign t_r12_c51_10 = t_r12_c51_7 + t_r12_c51_8;
  assign t_r12_c51_11 = t_r12_c51_9 + t_r12_c51_10;
  assign t_r12_c51_12 = t_r12_c51_11 + p_13_52;
  assign out_12_51 = t_r12_c51_12 >> 4;

  assign t_r12_c52_0 = p_11_52 << 1;
  assign t_r12_c52_1 = p_12_51 << 1;
  assign t_r12_c52_2 = p_12_52 << 2;
  assign t_r12_c52_3 = p_12_53 << 1;
  assign t_r12_c52_4 = p_13_52 << 1;
  assign t_r12_c52_5 = t_r12_c52_0 + p_11_51;
  assign t_r12_c52_6 = t_r12_c52_1 + p_11_53;
  assign t_r12_c52_7 = t_r12_c52_2 + t_r12_c52_3;
  assign t_r12_c52_8 = t_r12_c52_4 + p_13_51;
  assign t_r12_c52_9 = t_r12_c52_5 + t_r12_c52_6;
  assign t_r12_c52_10 = t_r12_c52_7 + t_r12_c52_8;
  assign t_r12_c52_11 = t_r12_c52_9 + t_r12_c52_10;
  assign t_r12_c52_12 = t_r12_c52_11 + p_13_53;
  assign out_12_52 = t_r12_c52_12 >> 4;

  assign t_r12_c53_0 = p_11_53 << 1;
  assign t_r12_c53_1 = p_12_52 << 1;
  assign t_r12_c53_2 = p_12_53 << 2;
  assign t_r12_c53_3 = p_12_54 << 1;
  assign t_r12_c53_4 = p_13_53 << 1;
  assign t_r12_c53_5 = t_r12_c53_0 + p_11_52;
  assign t_r12_c53_6 = t_r12_c53_1 + p_11_54;
  assign t_r12_c53_7 = t_r12_c53_2 + t_r12_c53_3;
  assign t_r12_c53_8 = t_r12_c53_4 + p_13_52;
  assign t_r12_c53_9 = t_r12_c53_5 + t_r12_c53_6;
  assign t_r12_c53_10 = t_r12_c53_7 + t_r12_c53_8;
  assign t_r12_c53_11 = t_r12_c53_9 + t_r12_c53_10;
  assign t_r12_c53_12 = t_r12_c53_11 + p_13_54;
  assign out_12_53 = t_r12_c53_12 >> 4;

  assign t_r12_c54_0 = p_11_54 << 1;
  assign t_r12_c54_1 = p_12_53 << 1;
  assign t_r12_c54_2 = p_12_54 << 2;
  assign t_r12_c54_3 = p_12_55 << 1;
  assign t_r12_c54_4 = p_13_54 << 1;
  assign t_r12_c54_5 = t_r12_c54_0 + p_11_53;
  assign t_r12_c54_6 = t_r12_c54_1 + p_11_55;
  assign t_r12_c54_7 = t_r12_c54_2 + t_r12_c54_3;
  assign t_r12_c54_8 = t_r12_c54_4 + p_13_53;
  assign t_r12_c54_9 = t_r12_c54_5 + t_r12_c54_6;
  assign t_r12_c54_10 = t_r12_c54_7 + t_r12_c54_8;
  assign t_r12_c54_11 = t_r12_c54_9 + t_r12_c54_10;
  assign t_r12_c54_12 = t_r12_c54_11 + p_13_55;
  assign out_12_54 = t_r12_c54_12 >> 4;

  assign t_r12_c55_0 = p_11_55 << 1;
  assign t_r12_c55_1 = p_12_54 << 1;
  assign t_r12_c55_2 = p_12_55 << 2;
  assign t_r12_c55_3 = p_12_56 << 1;
  assign t_r12_c55_4 = p_13_55 << 1;
  assign t_r12_c55_5 = t_r12_c55_0 + p_11_54;
  assign t_r12_c55_6 = t_r12_c55_1 + p_11_56;
  assign t_r12_c55_7 = t_r12_c55_2 + t_r12_c55_3;
  assign t_r12_c55_8 = t_r12_c55_4 + p_13_54;
  assign t_r12_c55_9 = t_r12_c55_5 + t_r12_c55_6;
  assign t_r12_c55_10 = t_r12_c55_7 + t_r12_c55_8;
  assign t_r12_c55_11 = t_r12_c55_9 + t_r12_c55_10;
  assign t_r12_c55_12 = t_r12_c55_11 + p_13_56;
  assign out_12_55 = t_r12_c55_12 >> 4;

  assign t_r12_c56_0 = p_11_56 << 1;
  assign t_r12_c56_1 = p_12_55 << 1;
  assign t_r12_c56_2 = p_12_56 << 2;
  assign t_r12_c56_3 = p_12_57 << 1;
  assign t_r12_c56_4 = p_13_56 << 1;
  assign t_r12_c56_5 = t_r12_c56_0 + p_11_55;
  assign t_r12_c56_6 = t_r12_c56_1 + p_11_57;
  assign t_r12_c56_7 = t_r12_c56_2 + t_r12_c56_3;
  assign t_r12_c56_8 = t_r12_c56_4 + p_13_55;
  assign t_r12_c56_9 = t_r12_c56_5 + t_r12_c56_6;
  assign t_r12_c56_10 = t_r12_c56_7 + t_r12_c56_8;
  assign t_r12_c56_11 = t_r12_c56_9 + t_r12_c56_10;
  assign t_r12_c56_12 = t_r12_c56_11 + p_13_57;
  assign out_12_56 = t_r12_c56_12 >> 4;

  assign t_r12_c57_0 = p_11_57 << 1;
  assign t_r12_c57_1 = p_12_56 << 1;
  assign t_r12_c57_2 = p_12_57 << 2;
  assign t_r12_c57_3 = p_12_58 << 1;
  assign t_r12_c57_4 = p_13_57 << 1;
  assign t_r12_c57_5 = t_r12_c57_0 + p_11_56;
  assign t_r12_c57_6 = t_r12_c57_1 + p_11_58;
  assign t_r12_c57_7 = t_r12_c57_2 + t_r12_c57_3;
  assign t_r12_c57_8 = t_r12_c57_4 + p_13_56;
  assign t_r12_c57_9 = t_r12_c57_5 + t_r12_c57_6;
  assign t_r12_c57_10 = t_r12_c57_7 + t_r12_c57_8;
  assign t_r12_c57_11 = t_r12_c57_9 + t_r12_c57_10;
  assign t_r12_c57_12 = t_r12_c57_11 + p_13_58;
  assign out_12_57 = t_r12_c57_12 >> 4;

  assign t_r12_c58_0 = p_11_58 << 1;
  assign t_r12_c58_1 = p_12_57 << 1;
  assign t_r12_c58_2 = p_12_58 << 2;
  assign t_r12_c58_3 = p_12_59 << 1;
  assign t_r12_c58_4 = p_13_58 << 1;
  assign t_r12_c58_5 = t_r12_c58_0 + p_11_57;
  assign t_r12_c58_6 = t_r12_c58_1 + p_11_59;
  assign t_r12_c58_7 = t_r12_c58_2 + t_r12_c58_3;
  assign t_r12_c58_8 = t_r12_c58_4 + p_13_57;
  assign t_r12_c58_9 = t_r12_c58_5 + t_r12_c58_6;
  assign t_r12_c58_10 = t_r12_c58_7 + t_r12_c58_8;
  assign t_r12_c58_11 = t_r12_c58_9 + t_r12_c58_10;
  assign t_r12_c58_12 = t_r12_c58_11 + p_13_59;
  assign out_12_58 = t_r12_c58_12 >> 4;

  assign t_r12_c59_0 = p_11_59 << 1;
  assign t_r12_c59_1 = p_12_58 << 1;
  assign t_r12_c59_2 = p_12_59 << 2;
  assign t_r12_c59_3 = p_12_60 << 1;
  assign t_r12_c59_4 = p_13_59 << 1;
  assign t_r12_c59_5 = t_r12_c59_0 + p_11_58;
  assign t_r12_c59_6 = t_r12_c59_1 + p_11_60;
  assign t_r12_c59_7 = t_r12_c59_2 + t_r12_c59_3;
  assign t_r12_c59_8 = t_r12_c59_4 + p_13_58;
  assign t_r12_c59_9 = t_r12_c59_5 + t_r12_c59_6;
  assign t_r12_c59_10 = t_r12_c59_7 + t_r12_c59_8;
  assign t_r12_c59_11 = t_r12_c59_9 + t_r12_c59_10;
  assign t_r12_c59_12 = t_r12_c59_11 + p_13_60;
  assign out_12_59 = t_r12_c59_12 >> 4;

  assign t_r12_c60_0 = p_11_60 << 1;
  assign t_r12_c60_1 = p_12_59 << 1;
  assign t_r12_c60_2 = p_12_60 << 2;
  assign t_r12_c60_3 = p_12_61 << 1;
  assign t_r12_c60_4 = p_13_60 << 1;
  assign t_r12_c60_5 = t_r12_c60_0 + p_11_59;
  assign t_r12_c60_6 = t_r12_c60_1 + p_11_61;
  assign t_r12_c60_7 = t_r12_c60_2 + t_r12_c60_3;
  assign t_r12_c60_8 = t_r12_c60_4 + p_13_59;
  assign t_r12_c60_9 = t_r12_c60_5 + t_r12_c60_6;
  assign t_r12_c60_10 = t_r12_c60_7 + t_r12_c60_8;
  assign t_r12_c60_11 = t_r12_c60_9 + t_r12_c60_10;
  assign t_r12_c60_12 = t_r12_c60_11 + p_13_61;
  assign out_12_60 = t_r12_c60_12 >> 4;

  assign t_r12_c61_0 = p_11_61 << 1;
  assign t_r12_c61_1 = p_12_60 << 1;
  assign t_r12_c61_2 = p_12_61 << 2;
  assign t_r12_c61_3 = p_12_62 << 1;
  assign t_r12_c61_4 = p_13_61 << 1;
  assign t_r12_c61_5 = t_r12_c61_0 + p_11_60;
  assign t_r12_c61_6 = t_r12_c61_1 + p_11_62;
  assign t_r12_c61_7 = t_r12_c61_2 + t_r12_c61_3;
  assign t_r12_c61_8 = t_r12_c61_4 + p_13_60;
  assign t_r12_c61_9 = t_r12_c61_5 + t_r12_c61_6;
  assign t_r12_c61_10 = t_r12_c61_7 + t_r12_c61_8;
  assign t_r12_c61_11 = t_r12_c61_9 + t_r12_c61_10;
  assign t_r12_c61_12 = t_r12_c61_11 + p_13_62;
  assign out_12_61 = t_r12_c61_12 >> 4;

  assign t_r12_c62_0 = p_11_62 << 1;
  assign t_r12_c62_1 = p_12_61 << 1;
  assign t_r12_c62_2 = p_12_62 << 2;
  assign t_r12_c62_3 = p_12_63 << 1;
  assign t_r12_c62_4 = p_13_62 << 1;
  assign t_r12_c62_5 = t_r12_c62_0 + p_11_61;
  assign t_r12_c62_6 = t_r12_c62_1 + p_11_63;
  assign t_r12_c62_7 = t_r12_c62_2 + t_r12_c62_3;
  assign t_r12_c62_8 = t_r12_c62_4 + p_13_61;
  assign t_r12_c62_9 = t_r12_c62_5 + t_r12_c62_6;
  assign t_r12_c62_10 = t_r12_c62_7 + t_r12_c62_8;
  assign t_r12_c62_11 = t_r12_c62_9 + t_r12_c62_10;
  assign t_r12_c62_12 = t_r12_c62_11 + p_13_63;
  assign out_12_62 = t_r12_c62_12 >> 4;

  assign t_r12_c63_0 = p_11_63 << 1;
  assign t_r12_c63_1 = p_12_62 << 1;
  assign t_r12_c63_2 = p_12_63 << 2;
  assign t_r12_c63_3 = p_12_64 << 1;
  assign t_r12_c63_4 = p_13_63 << 1;
  assign t_r12_c63_5 = t_r12_c63_0 + p_11_62;
  assign t_r12_c63_6 = t_r12_c63_1 + p_11_64;
  assign t_r12_c63_7 = t_r12_c63_2 + t_r12_c63_3;
  assign t_r12_c63_8 = t_r12_c63_4 + p_13_62;
  assign t_r12_c63_9 = t_r12_c63_5 + t_r12_c63_6;
  assign t_r12_c63_10 = t_r12_c63_7 + t_r12_c63_8;
  assign t_r12_c63_11 = t_r12_c63_9 + t_r12_c63_10;
  assign t_r12_c63_12 = t_r12_c63_11 + p_13_64;
  assign out_12_63 = t_r12_c63_12 >> 4;

  assign t_r12_c64_0 = p_11_64 << 1;
  assign t_r12_c64_1 = p_12_63 << 1;
  assign t_r12_c64_2 = p_12_64 << 2;
  assign t_r12_c64_3 = p_12_65 << 1;
  assign t_r12_c64_4 = p_13_64 << 1;
  assign t_r12_c64_5 = t_r12_c64_0 + p_11_63;
  assign t_r12_c64_6 = t_r12_c64_1 + p_11_65;
  assign t_r12_c64_7 = t_r12_c64_2 + t_r12_c64_3;
  assign t_r12_c64_8 = t_r12_c64_4 + p_13_63;
  assign t_r12_c64_9 = t_r12_c64_5 + t_r12_c64_6;
  assign t_r12_c64_10 = t_r12_c64_7 + t_r12_c64_8;
  assign t_r12_c64_11 = t_r12_c64_9 + t_r12_c64_10;
  assign t_r12_c64_12 = t_r12_c64_11 + p_13_65;
  assign out_12_64 = t_r12_c64_12 >> 4;

  assign t_r13_c1_0 = p_12_1 << 1;
  assign t_r13_c1_1 = p_13_0 << 1;
  assign t_r13_c1_2 = p_13_1 << 2;
  assign t_r13_c1_3 = p_13_2 << 1;
  assign t_r13_c1_4 = p_14_1 << 1;
  assign t_r13_c1_5 = t_r13_c1_0 + p_12_0;
  assign t_r13_c1_6 = t_r13_c1_1 + p_12_2;
  assign t_r13_c1_7 = t_r13_c1_2 + t_r13_c1_3;
  assign t_r13_c1_8 = t_r13_c1_4 + p_14_0;
  assign t_r13_c1_9 = t_r13_c1_5 + t_r13_c1_6;
  assign t_r13_c1_10 = t_r13_c1_7 + t_r13_c1_8;
  assign t_r13_c1_11 = t_r13_c1_9 + t_r13_c1_10;
  assign t_r13_c1_12 = t_r13_c1_11 + p_14_2;
  assign out_13_1 = t_r13_c1_12 >> 4;

  assign t_r13_c2_0 = p_12_2 << 1;
  assign t_r13_c2_1 = p_13_1 << 1;
  assign t_r13_c2_2 = p_13_2 << 2;
  assign t_r13_c2_3 = p_13_3 << 1;
  assign t_r13_c2_4 = p_14_2 << 1;
  assign t_r13_c2_5 = t_r13_c2_0 + p_12_1;
  assign t_r13_c2_6 = t_r13_c2_1 + p_12_3;
  assign t_r13_c2_7 = t_r13_c2_2 + t_r13_c2_3;
  assign t_r13_c2_8 = t_r13_c2_4 + p_14_1;
  assign t_r13_c2_9 = t_r13_c2_5 + t_r13_c2_6;
  assign t_r13_c2_10 = t_r13_c2_7 + t_r13_c2_8;
  assign t_r13_c2_11 = t_r13_c2_9 + t_r13_c2_10;
  assign t_r13_c2_12 = t_r13_c2_11 + p_14_3;
  assign out_13_2 = t_r13_c2_12 >> 4;

  assign t_r13_c3_0 = p_12_3 << 1;
  assign t_r13_c3_1 = p_13_2 << 1;
  assign t_r13_c3_2 = p_13_3 << 2;
  assign t_r13_c3_3 = p_13_4 << 1;
  assign t_r13_c3_4 = p_14_3 << 1;
  assign t_r13_c3_5 = t_r13_c3_0 + p_12_2;
  assign t_r13_c3_6 = t_r13_c3_1 + p_12_4;
  assign t_r13_c3_7 = t_r13_c3_2 + t_r13_c3_3;
  assign t_r13_c3_8 = t_r13_c3_4 + p_14_2;
  assign t_r13_c3_9 = t_r13_c3_5 + t_r13_c3_6;
  assign t_r13_c3_10 = t_r13_c3_7 + t_r13_c3_8;
  assign t_r13_c3_11 = t_r13_c3_9 + t_r13_c3_10;
  assign t_r13_c3_12 = t_r13_c3_11 + p_14_4;
  assign out_13_3 = t_r13_c3_12 >> 4;

  assign t_r13_c4_0 = p_12_4 << 1;
  assign t_r13_c4_1 = p_13_3 << 1;
  assign t_r13_c4_2 = p_13_4 << 2;
  assign t_r13_c4_3 = p_13_5 << 1;
  assign t_r13_c4_4 = p_14_4 << 1;
  assign t_r13_c4_5 = t_r13_c4_0 + p_12_3;
  assign t_r13_c4_6 = t_r13_c4_1 + p_12_5;
  assign t_r13_c4_7 = t_r13_c4_2 + t_r13_c4_3;
  assign t_r13_c4_8 = t_r13_c4_4 + p_14_3;
  assign t_r13_c4_9 = t_r13_c4_5 + t_r13_c4_6;
  assign t_r13_c4_10 = t_r13_c4_7 + t_r13_c4_8;
  assign t_r13_c4_11 = t_r13_c4_9 + t_r13_c4_10;
  assign t_r13_c4_12 = t_r13_c4_11 + p_14_5;
  assign out_13_4 = t_r13_c4_12 >> 4;

  assign t_r13_c5_0 = p_12_5 << 1;
  assign t_r13_c5_1 = p_13_4 << 1;
  assign t_r13_c5_2 = p_13_5 << 2;
  assign t_r13_c5_3 = p_13_6 << 1;
  assign t_r13_c5_4 = p_14_5 << 1;
  assign t_r13_c5_5 = t_r13_c5_0 + p_12_4;
  assign t_r13_c5_6 = t_r13_c5_1 + p_12_6;
  assign t_r13_c5_7 = t_r13_c5_2 + t_r13_c5_3;
  assign t_r13_c5_8 = t_r13_c5_4 + p_14_4;
  assign t_r13_c5_9 = t_r13_c5_5 + t_r13_c5_6;
  assign t_r13_c5_10 = t_r13_c5_7 + t_r13_c5_8;
  assign t_r13_c5_11 = t_r13_c5_9 + t_r13_c5_10;
  assign t_r13_c5_12 = t_r13_c5_11 + p_14_6;
  assign out_13_5 = t_r13_c5_12 >> 4;

  assign t_r13_c6_0 = p_12_6 << 1;
  assign t_r13_c6_1 = p_13_5 << 1;
  assign t_r13_c6_2 = p_13_6 << 2;
  assign t_r13_c6_3 = p_13_7 << 1;
  assign t_r13_c6_4 = p_14_6 << 1;
  assign t_r13_c6_5 = t_r13_c6_0 + p_12_5;
  assign t_r13_c6_6 = t_r13_c6_1 + p_12_7;
  assign t_r13_c6_7 = t_r13_c6_2 + t_r13_c6_3;
  assign t_r13_c6_8 = t_r13_c6_4 + p_14_5;
  assign t_r13_c6_9 = t_r13_c6_5 + t_r13_c6_6;
  assign t_r13_c6_10 = t_r13_c6_7 + t_r13_c6_8;
  assign t_r13_c6_11 = t_r13_c6_9 + t_r13_c6_10;
  assign t_r13_c6_12 = t_r13_c6_11 + p_14_7;
  assign out_13_6 = t_r13_c6_12 >> 4;

  assign t_r13_c7_0 = p_12_7 << 1;
  assign t_r13_c7_1 = p_13_6 << 1;
  assign t_r13_c7_2 = p_13_7 << 2;
  assign t_r13_c7_3 = p_13_8 << 1;
  assign t_r13_c7_4 = p_14_7 << 1;
  assign t_r13_c7_5 = t_r13_c7_0 + p_12_6;
  assign t_r13_c7_6 = t_r13_c7_1 + p_12_8;
  assign t_r13_c7_7 = t_r13_c7_2 + t_r13_c7_3;
  assign t_r13_c7_8 = t_r13_c7_4 + p_14_6;
  assign t_r13_c7_9 = t_r13_c7_5 + t_r13_c7_6;
  assign t_r13_c7_10 = t_r13_c7_7 + t_r13_c7_8;
  assign t_r13_c7_11 = t_r13_c7_9 + t_r13_c7_10;
  assign t_r13_c7_12 = t_r13_c7_11 + p_14_8;
  assign out_13_7 = t_r13_c7_12 >> 4;

  assign t_r13_c8_0 = p_12_8 << 1;
  assign t_r13_c8_1 = p_13_7 << 1;
  assign t_r13_c8_2 = p_13_8 << 2;
  assign t_r13_c8_3 = p_13_9 << 1;
  assign t_r13_c8_4 = p_14_8 << 1;
  assign t_r13_c8_5 = t_r13_c8_0 + p_12_7;
  assign t_r13_c8_6 = t_r13_c8_1 + p_12_9;
  assign t_r13_c8_7 = t_r13_c8_2 + t_r13_c8_3;
  assign t_r13_c8_8 = t_r13_c8_4 + p_14_7;
  assign t_r13_c8_9 = t_r13_c8_5 + t_r13_c8_6;
  assign t_r13_c8_10 = t_r13_c8_7 + t_r13_c8_8;
  assign t_r13_c8_11 = t_r13_c8_9 + t_r13_c8_10;
  assign t_r13_c8_12 = t_r13_c8_11 + p_14_9;
  assign out_13_8 = t_r13_c8_12 >> 4;

  assign t_r13_c9_0 = p_12_9 << 1;
  assign t_r13_c9_1 = p_13_8 << 1;
  assign t_r13_c9_2 = p_13_9 << 2;
  assign t_r13_c9_3 = p_13_10 << 1;
  assign t_r13_c9_4 = p_14_9 << 1;
  assign t_r13_c9_5 = t_r13_c9_0 + p_12_8;
  assign t_r13_c9_6 = t_r13_c9_1 + p_12_10;
  assign t_r13_c9_7 = t_r13_c9_2 + t_r13_c9_3;
  assign t_r13_c9_8 = t_r13_c9_4 + p_14_8;
  assign t_r13_c9_9 = t_r13_c9_5 + t_r13_c9_6;
  assign t_r13_c9_10 = t_r13_c9_7 + t_r13_c9_8;
  assign t_r13_c9_11 = t_r13_c9_9 + t_r13_c9_10;
  assign t_r13_c9_12 = t_r13_c9_11 + p_14_10;
  assign out_13_9 = t_r13_c9_12 >> 4;

  assign t_r13_c10_0 = p_12_10 << 1;
  assign t_r13_c10_1 = p_13_9 << 1;
  assign t_r13_c10_2 = p_13_10 << 2;
  assign t_r13_c10_3 = p_13_11 << 1;
  assign t_r13_c10_4 = p_14_10 << 1;
  assign t_r13_c10_5 = t_r13_c10_0 + p_12_9;
  assign t_r13_c10_6 = t_r13_c10_1 + p_12_11;
  assign t_r13_c10_7 = t_r13_c10_2 + t_r13_c10_3;
  assign t_r13_c10_8 = t_r13_c10_4 + p_14_9;
  assign t_r13_c10_9 = t_r13_c10_5 + t_r13_c10_6;
  assign t_r13_c10_10 = t_r13_c10_7 + t_r13_c10_8;
  assign t_r13_c10_11 = t_r13_c10_9 + t_r13_c10_10;
  assign t_r13_c10_12 = t_r13_c10_11 + p_14_11;
  assign out_13_10 = t_r13_c10_12 >> 4;

  assign t_r13_c11_0 = p_12_11 << 1;
  assign t_r13_c11_1 = p_13_10 << 1;
  assign t_r13_c11_2 = p_13_11 << 2;
  assign t_r13_c11_3 = p_13_12 << 1;
  assign t_r13_c11_4 = p_14_11 << 1;
  assign t_r13_c11_5 = t_r13_c11_0 + p_12_10;
  assign t_r13_c11_6 = t_r13_c11_1 + p_12_12;
  assign t_r13_c11_7 = t_r13_c11_2 + t_r13_c11_3;
  assign t_r13_c11_8 = t_r13_c11_4 + p_14_10;
  assign t_r13_c11_9 = t_r13_c11_5 + t_r13_c11_6;
  assign t_r13_c11_10 = t_r13_c11_7 + t_r13_c11_8;
  assign t_r13_c11_11 = t_r13_c11_9 + t_r13_c11_10;
  assign t_r13_c11_12 = t_r13_c11_11 + p_14_12;
  assign out_13_11 = t_r13_c11_12 >> 4;

  assign t_r13_c12_0 = p_12_12 << 1;
  assign t_r13_c12_1 = p_13_11 << 1;
  assign t_r13_c12_2 = p_13_12 << 2;
  assign t_r13_c12_3 = p_13_13 << 1;
  assign t_r13_c12_4 = p_14_12 << 1;
  assign t_r13_c12_5 = t_r13_c12_0 + p_12_11;
  assign t_r13_c12_6 = t_r13_c12_1 + p_12_13;
  assign t_r13_c12_7 = t_r13_c12_2 + t_r13_c12_3;
  assign t_r13_c12_8 = t_r13_c12_4 + p_14_11;
  assign t_r13_c12_9 = t_r13_c12_5 + t_r13_c12_6;
  assign t_r13_c12_10 = t_r13_c12_7 + t_r13_c12_8;
  assign t_r13_c12_11 = t_r13_c12_9 + t_r13_c12_10;
  assign t_r13_c12_12 = t_r13_c12_11 + p_14_13;
  assign out_13_12 = t_r13_c12_12 >> 4;

  assign t_r13_c13_0 = p_12_13 << 1;
  assign t_r13_c13_1 = p_13_12 << 1;
  assign t_r13_c13_2 = p_13_13 << 2;
  assign t_r13_c13_3 = p_13_14 << 1;
  assign t_r13_c13_4 = p_14_13 << 1;
  assign t_r13_c13_5 = t_r13_c13_0 + p_12_12;
  assign t_r13_c13_6 = t_r13_c13_1 + p_12_14;
  assign t_r13_c13_7 = t_r13_c13_2 + t_r13_c13_3;
  assign t_r13_c13_8 = t_r13_c13_4 + p_14_12;
  assign t_r13_c13_9 = t_r13_c13_5 + t_r13_c13_6;
  assign t_r13_c13_10 = t_r13_c13_7 + t_r13_c13_8;
  assign t_r13_c13_11 = t_r13_c13_9 + t_r13_c13_10;
  assign t_r13_c13_12 = t_r13_c13_11 + p_14_14;
  assign out_13_13 = t_r13_c13_12 >> 4;

  assign t_r13_c14_0 = p_12_14 << 1;
  assign t_r13_c14_1 = p_13_13 << 1;
  assign t_r13_c14_2 = p_13_14 << 2;
  assign t_r13_c14_3 = p_13_15 << 1;
  assign t_r13_c14_4 = p_14_14 << 1;
  assign t_r13_c14_5 = t_r13_c14_0 + p_12_13;
  assign t_r13_c14_6 = t_r13_c14_1 + p_12_15;
  assign t_r13_c14_7 = t_r13_c14_2 + t_r13_c14_3;
  assign t_r13_c14_8 = t_r13_c14_4 + p_14_13;
  assign t_r13_c14_9 = t_r13_c14_5 + t_r13_c14_6;
  assign t_r13_c14_10 = t_r13_c14_7 + t_r13_c14_8;
  assign t_r13_c14_11 = t_r13_c14_9 + t_r13_c14_10;
  assign t_r13_c14_12 = t_r13_c14_11 + p_14_15;
  assign out_13_14 = t_r13_c14_12 >> 4;

  assign t_r13_c15_0 = p_12_15 << 1;
  assign t_r13_c15_1 = p_13_14 << 1;
  assign t_r13_c15_2 = p_13_15 << 2;
  assign t_r13_c15_3 = p_13_16 << 1;
  assign t_r13_c15_4 = p_14_15 << 1;
  assign t_r13_c15_5 = t_r13_c15_0 + p_12_14;
  assign t_r13_c15_6 = t_r13_c15_1 + p_12_16;
  assign t_r13_c15_7 = t_r13_c15_2 + t_r13_c15_3;
  assign t_r13_c15_8 = t_r13_c15_4 + p_14_14;
  assign t_r13_c15_9 = t_r13_c15_5 + t_r13_c15_6;
  assign t_r13_c15_10 = t_r13_c15_7 + t_r13_c15_8;
  assign t_r13_c15_11 = t_r13_c15_9 + t_r13_c15_10;
  assign t_r13_c15_12 = t_r13_c15_11 + p_14_16;
  assign out_13_15 = t_r13_c15_12 >> 4;

  assign t_r13_c16_0 = p_12_16 << 1;
  assign t_r13_c16_1 = p_13_15 << 1;
  assign t_r13_c16_2 = p_13_16 << 2;
  assign t_r13_c16_3 = p_13_17 << 1;
  assign t_r13_c16_4 = p_14_16 << 1;
  assign t_r13_c16_5 = t_r13_c16_0 + p_12_15;
  assign t_r13_c16_6 = t_r13_c16_1 + p_12_17;
  assign t_r13_c16_7 = t_r13_c16_2 + t_r13_c16_3;
  assign t_r13_c16_8 = t_r13_c16_4 + p_14_15;
  assign t_r13_c16_9 = t_r13_c16_5 + t_r13_c16_6;
  assign t_r13_c16_10 = t_r13_c16_7 + t_r13_c16_8;
  assign t_r13_c16_11 = t_r13_c16_9 + t_r13_c16_10;
  assign t_r13_c16_12 = t_r13_c16_11 + p_14_17;
  assign out_13_16 = t_r13_c16_12 >> 4;

  assign t_r13_c17_0 = p_12_17 << 1;
  assign t_r13_c17_1 = p_13_16 << 1;
  assign t_r13_c17_2 = p_13_17 << 2;
  assign t_r13_c17_3 = p_13_18 << 1;
  assign t_r13_c17_4 = p_14_17 << 1;
  assign t_r13_c17_5 = t_r13_c17_0 + p_12_16;
  assign t_r13_c17_6 = t_r13_c17_1 + p_12_18;
  assign t_r13_c17_7 = t_r13_c17_2 + t_r13_c17_3;
  assign t_r13_c17_8 = t_r13_c17_4 + p_14_16;
  assign t_r13_c17_9 = t_r13_c17_5 + t_r13_c17_6;
  assign t_r13_c17_10 = t_r13_c17_7 + t_r13_c17_8;
  assign t_r13_c17_11 = t_r13_c17_9 + t_r13_c17_10;
  assign t_r13_c17_12 = t_r13_c17_11 + p_14_18;
  assign out_13_17 = t_r13_c17_12 >> 4;

  assign t_r13_c18_0 = p_12_18 << 1;
  assign t_r13_c18_1 = p_13_17 << 1;
  assign t_r13_c18_2 = p_13_18 << 2;
  assign t_r13_c18_3 = p_13_19 << 1;
  assign t_r13_c18_4 = p_14_18 << 1;
  assign t_r13_c18_5 = t_r13_c18_0 + p_12_17;
  assign t_r13_c18_6 = t_r13_c18_1 + p_12_19;
  assign t_r13_c18_7 = t_r13_c18_2 + t_r13_c18_3;
  assign t_r13_c18_8 = t_r13_c18_4 + p_14_17;
  assign t_r13_c18_9 = t_r13_c18_5 + t_r13_c18_6;
  assign t_r13_c18_10 = t_r13_c18_7 + t_r13_c18_8;
  assign t_r13_c18_11 = t_r13_c18_9 + t_r13_c18_10;
  assign t_r13_c18_12 = t_r13_c18_11 + p_14_19;
  assign out_13_18 = t_r13_c18_12 >> 4;

  assign t_r13_c19_0 = p_12_19 << 1;
  assign t_r13_c19_1 = p_13_18 << 1;
  assign t_r13_c19_2 = p_13_19 << 2;
  assign t_r13_c19_3 = p_13_20 << 1;
  assign t_r13_c19_4 = p_14_19 << 1;
  assign t_r13_c19_5 = t_r13_c19_0 + p_12_18;
  assign t_r13_c19_6 = t_r13_c19_1 + p_12_20;
  assign t_r13_c19_7 = t_r13_c19_2 + t_r13_c19_3;
  assign t_r13_c19_8 = t_r13_c19_4 + p_14_18;
  assign t_r13_c19_9 = t_r13_c19_5 + t_r13_c19_6;
  assign t_r13_c19_10 = t_r13_c19_7 + t_r13_c19_8;
  assign t_r13_c19_11 = t_r13_c19_9 + t_r13_c19_10;
  assign t_r13_c19_12 = t_r13_c19_11 + p_14_20;
  assign out_13_19 = t_r13_c19_12 >> 4;

  assign t_r13_c20_0 = p_12_20 << 1;
  assign t_r13_c20_1 = p_13_19 << 1;
  assign t_r13_c20_2 = p_13_20 << 2;
  assign t_r13_c20_3 = p_13_21 << 1;
  assign t_r13_c20_4 = p_14_20 << 1;
  assign t_r13_c20_5 = t_r13_c20_0 + p_12_19;
  assign t_r13_c20_6 = t_r13_c20_1 + p_12_21;
  assign t_r13_c20_7 = t_r13_c20_2 + t_r13_c20_3;
  assign t_r13_c20_8 = t_r13_c20_4 + p_14_19;
  assign t_r13_c20_9 = t_r13_c20_5 + t_r13_c20_6;
  assign t_r13_c20_10 = t_r13_c20_7 + t_r13_c20_8;
  assign t_r13_c20_11 = t_r13_c20_9 + t_r13_c20_10;
  assign t_r13_c20_12 = t_r13_c20_11 + p_14_21;
  assign out_13_20 = t_r13_c20_12 >> 4;

  assign t_r13_c21_0 = p_12_21 << 1;
  assign t_r13_c21_1 = p_13_20 << 1;
  assign t_r13_c21_2 = p_13_21 << 2;
  assign t_r13_c21_3 = p_13_22 << 1;
  assign t_r13_c21_4 = p_14_21 << 1;
  assign t_r13_c21_5 = t_r13_c21_0 + p_12_20;
  assign t_r13_c21_6 = t_r13_c21_1 + p_12_22;
  assign t_r13_c21_7 = t_r13_c21_2 + t_r13_c21_3;
  assign t_r13_c21_8 = t_r13_c21_4 + p_14_20;
  assign t_r13_c21_9 = t_r13_c21_5 + t_r13_c21_6;
  assign t_r13_c21_10 = t_r13_c21_7 + t_r13_c21_8;
  assign t_r13_c21_11 = t_r13_c21_9 + t_r13_c21_10;
  assign t_r13_c21_12 = t_r13_c21_11 + p_14_22;
  assign out_13_21 = t_r13_c21_12 >> 4;

  assign t_r13_c22_0 = p_12_22 << 1;
  assign t_r13_c22_1 = p_13_21 << 1;
  assign t_r13_c22_2 = p_13_22 << 2;
  assign t_r13_c22_3 = p_13_23 << 1;
  assign t_r13_c22_4 = p_14_22 << 1;
  assign t_r13_c22_5 = t_r13_c22_0 + p_12_21;
  assign t_r13_c22_6 = t_r13_c22_1 + p_12_23;
  assign t_r13_c22_7 = t_r13_c22_2 + t_r13_c22_3;
  assign t_r13_c22_8 = t_r13_c22_4 + p_14_21;
  assign t_r13_c22_9 = t_r13_c22_5 + t_r13_c22_6;
  assign t_r13_c22_10 = t_r13_c22_7 + t_r13_c22_8;
  assign t_r13_c22_11 = t_r13_c22_9 + t_r13_c22_10;
  assign t_r13_c22_12 = t_r13_c22_11 + p_14_23;
  assign out_13_22 = t_r13_c22_12 >> 4;

  assign t_r13_c23_0 = p_12_23 << 1;
  assign t_r13_c23_1 = p_13_22 << 1;
  assign t_r13_c23_2 = p_13_23 << 2;
  assign t_r13_c23_3 = p_13_24 << 1;
  assign t_r13_c23_4 = p_14_23 << 1;
  assign t_r13_c23_5 = t_r13_c23_0 + p_12_22;
  assign t_r13_c23_6 = t_r13_c23_1 + p_12_24;
  assign t_r13_c23_7 = t_r13_c23_2 + t_r13_c23_3;
  assign t_r13_c23_8 = t_r13_c23_4 + p_14_22;
  assign t_r13_c23_9 = t_r13_c23_5 + t_r13_c23_6;
  assign t_r13_c23_10 = t_r13_c23_7 + t_r13_c23_8;
  assign t_r13_c23_11 = t_r13_c23_9 + t_r13_c23_10;
  assign t_r13_c23_12 = t_r13_c23_11 + p_14_24;
  assign out_13_23 = t_r13_c23_12 >> 4;

  assign t_r13_c24_0 = p_12_24 << 1;
  assign t_r13_c24_1 = p_13_23 << 1;
  assign t_r13_c24_2 = p_13_24 << 2;
  assign t_r13_c24_3 = p_13_25 << 1;
  assign t_r13_c24_4 = p_14_24 << 1;
  assign t_r13_c24_5 = t_r13_c24_0 + p_12_23;
  assign t_r13_c24_6 = t_r13_c24_1 + p_12_25;
  assign t_r13_c24_7 = t_r13_c24_2 + t_r13_c24_3;
  assign t_r13_c24_8 = t_r13_c24_4 + p_14_23;
  assign t_r13_c24_9 = t_r13_c24_5 + t_r13_c24_6;
  assign t_r13_c24_10 = t_r13_c24_7 + t_r13_c24_8;
  assign t_r13_c24_11 = t_r13_c24_9 + t_r13_c24_10;
  assign t_r13_c24_12 = t_r13_c24_11 + p_14_25;
  assign out_13_24 = t_r13_c24_12 >> 4;

  assign t_r13_c25_0 = p_12_25 << 1;
  assign t_r13_c25_1 = p_13_24 << 1;
  assign t_r13_c25_2 = p_13_25 << 2;
  assign t_r13_c25_3 = p_13_26 << 1;
  assign t_r13_c25_4 = p_14_25 << 1;
  assign t_r13_c25_5 = t_r13_c25_0 + p_12_24;
  assign t_r13_c25_6 = t_r13_c25_1 + p_12_26;
  assign t_r13_c25_7 = t_r13_c25_2 + t_r13_c25_3;
  assign t_r13_c25_8 = t_r13_c25_4 + p_14_24;
  assign t_r13_c25_9 = t_r13_c25_5 + t_r13_c25_6;
  assign t_r13_c25_10 = t_r13_c25_7 + t_r13_c25_8;
  assign t_r13_c25_11 = t_r13_c25_9 + t_r13_c25_10;
  assign t_r13_c25_12 = t_r13_c25_11 + p_14_26;
  assign out_13_25 = t_r13_c25_12 >> 4;

  assign t_r13_c26_0 = p_12_26 << 1;
  assign t_r13_c26_1 = p_13_25 << 1;
  assign t_r13_c26_2 = p_13_26 << 2;
  assign t_r13_c26_3 = p_13_27 << 1;
  assign t_r13_c26_4 = p_14_26 << 1;
  assign t_r13_c26_5 = t_r13_c26_0 + p_12_25;
  assign t_r13_c26_6 = t_r13_c26_1 + p_12_27;
  assign t_r13_c26_7 = t_r13_c26_2 + t_r13_c26_3;
  assign t_r13_c26_8 = t_r13_c26_4 + p_14_25;
  assign t_r13_c26_9 = t_r13_c26_5 + t_r13_c26_6;
  assign t_r13_c26_10 = t_r13_c26_7 + t_r13_c26_8;
  assign t_r13_c26_11 = t_r13_c26_9 + t_r13_c26_10;
  assign t_r13_c26_12 = t_r13_c26_11 + p_14_27;
  assign out_13_26 = t_r13_c26_12 >> 4;

  assign t_r13_c27_0 = p_12_27 << 1;
  assign t_r13_c27_1 = p_13_26 << 1;
  assign t_r13_c27_2 = p_13_27 << 2;
  assign t_r13_c27_3 = p_13_28 << 1;
  assign t_r13_c27_4 = p_14_27 << 1;
  assign t_r13_c27_5 = t_r13_c27_0 + p_12_26;
  assign t_r13_c27_6 = t_r13_c27_1 + p_12_28;
  assign t_r13_c27_7 = t_r13_c27_2 + t_r13_c27_3;
  assign t_r13_c27_8 = t_r13_c27_4 + p_14_26;
  assign t_r13_c27_9 = t_r13_c27_5 + t_r13_c27_6;
  assign t_r13_c27_10 = t_r13_c27_7 + t_r13_c27_8;
  assign t_r13_c27_11 = t_r13_c27_9 + t_r13_c27_10;
  assign t_r13_c27_12 = t_r13_c27_11 + p_14_28;
  assign out_13_27 = t_r13_c27_12 >> 4;

  assign t_r13_c28_0 = p_12_28 << 1;
  assign t_r13_c28_1 = p_13_27 << 1;
  assign t_r13_c28_2 = p_13_28 << 2;
  assign t_r13_c28_3 = p_13_29 << 1;
  assign t_r13_c28_4 = p_14_28 << 1;
  assign t_r13_c28_5 = t_r13_c28_0 + p_12_27;
  assign t_r13_c28_6 = t_r13_c28_1 + p_12_29;
  assign t_r13_c28_7 = t_r13_c28_2 + t_r13_c28_3;
  assign t_r13_c28_8 = t_r13_c28_4 + p_14_27;
  assign t_r13_c28_9 = t_r13_c28_5 + t_r13_c28_6;
  assign t_r13_c28_10 = t_r13_c28_7 + t_r13_c28_8;
  assign t_r13_c28_11 = t_r13_c28_9 + t_r13_c28_10;
  assign t_r13_c28_12 = t_r13_c28_11 + p_14_29;
  assign out_13_28 = t_r13_c28_12 >> 4;

  assign t_r13_c29_0 = p_12_29 << 1;
  assign t_r13_c29_1 = p_13_28 << 1;
  assign t_r13_c29_2 = p_13_29 << 2;
  assign t_r13_c29_3 = p_13_30 << 1;
  assign t_r13_c29_4 = p_14_29 << 1;
  assign t_r13_c29_5 = t_r13_c29_0 + p_12_28;
  assign t_r13_c29_6 = t_r13_c29_1 + p_12_30;
  assign t_r13_c29_7 = t_r13_c29_2 + t_r13_c29_3;
  assign t_r13_c29_8 = t_r13_c29_4 + p_14_28;
  assign t_r13_c29_9 = t_r13_c29_5 + t_r13_c29_6;
  assign t_r13_c29_10 = t_r13_c29_7 + t_r13_c29_8;
  assign t_r13_c29_11 = t_r13_c29_9 + t_r13_c29_10;
  assign t_r13_c29_12 = t_r13_c29_11 + p_14_30;
  assign out_13_29 = t_r13_c29_12 >> 4;

  assign t_r13_c30_0 = p_12_30 << 1;
  assign t_r13_c30_1 = p_13_29 << 1;
  assign t_r13_c30_2 = p_13_30 << 2;
  assign t_r13_c30_3 = p_13_31 << 1;
  assign t_r13_c30_4 = p_14_30 << 1;
  assign t_r13_c30_5 = t_r13_c30_0 + p_12_29;
  assign t_r13_c30_6 = t_r13_c30_1 + p_12_31;
  assign t_r13_c30_7 = t_r13_c30_2 + t_r13_c30_3;
  assign t_r13_c30_8 = t_r13_c30_4 + p_14_29;
  assign t_r13_c30_9 = t_r13_c30_5 + t_r13_c30_6;
  assign t_r13_c30_10 = t_r13_c30_7 + t_r13_c30_8;
  assign t_r13_c30_11 = t_r13_c30_9 + t_r13_c30_10;
  assign t_r13_c30_12 = t_r13_c30_11 + p_14_31;
  assign out_13_30 = t_r13_c30_12 >> 4;

  assign t_r13_c31_0 = p_12_31 << 1;
  assign t_r13_c31_1 = p_13_30 << 1;
  assign t_r13_c31_2 = p_13_31 << 2;
  assign t_r13_c31_3 = p_13_32 << 1;
  assign t_r13_c31_4 = p_14_31 << 1;
  assign t_r13_c31_5 = t_r13_c31_0 + p_12_30;
  assign t_r13_c31_6 = t_r13_c31_1 + p_12_32;
  assign t_r13_c31_7 = t_r13_c31_2 + t_r13_c31_3;
  assign t_r13_c31_8 = t_r13_c31_4 + p_14_30;
  assign t_r13_c31_9 = t_r13_c31_5 + t_r13_c31_6;
  assign t_r13_c31_10 = t_r13_c31_7 + t_r13_c31_8;
  assign t_r13_c31_11 = t_r13_c31_9 + t_r13_c31_10;
  assign t_r13_c31_12 = t_r13_c31_11 + p_14_32;
  assign out_13_31 = t_r13_c31_12 >> 4;

  assign t_r13_c32_0 = p_12_32 << 1;
  assign t_r13_c32_1 = p_13_31 << 1;
  assign t_r13_c32_2 = p_13_32 << 2;
  assign t_r13_c32_3 = p_13_33 << 1;
  assign t_r13_c32_4 = p_14_32 << 1;
  assign t_r13_c32_5 = t_r13_c32_0 + p_12_31;
  assign t_r13_c32_6 = t_r13_c32_1 + p_12_33;
  assign t_r13_c32_7 = t_r13_c32_2 + t_r13_c32_3;
  assign t_r13_c32_8 = t_r13_c32_4 + p_14_31;
  assign t_r13_c32_9 = t_r13_c32_5 + t_r13_c32_6;
  assign t_r13_c32_10 = t_r13_c32_7 + t_r13_c32_8;
  assign t_r13_c32_11 = t_r13_c32_9 + t_r13_c32_10;
  assign t_r13_c32_12 = t_r13_c32_11 + p_14_33;
  assign out_13_32 = t_r13_c32_12 >> 4;

  assign t_r13_c33_0 = p_12_33 << 1;
  assign t_r13_c33_1 = p_13_32 << 1;
  assign t_r13_c33_2 = p_13_33 << 2;
  assign t_r13_c33_3 = p_13_34 << 1;
  assign t_r13_c33_4 = p_14_33 << 1;
  assign t_r13_c33_5 = t_r13_c33_0 + p_12_32;
  assign t_r13_c33_6 = t_r13_c33_1 + p_12_34;
  assign t_r13_c33_7 = t_r13_c33_2 + t_r13_c33_3;
  assign t_r13_c33_8 = t_r13_c33_4 + p_14_32;
  assign t_r13_c33_9 = t_r13_c33_5 + t_r13_c33_6;
  assign t_r13_c33_10 = t_r13_c33_7 + t_r13_c33_8;
  assign t_r13_c33_11 = t_r13_c33_9 + t_r13_c33_10;
  assign t_r13_c33_12 = t_r13_c33_11 + p_14_34;
  assign out_13_33 = t_r13_c33_12 >> 4;

  assign t_r13_c34_0 = p_12_34 << 1;
  assign t_r13_c34_1 = p_13_33 << 1;
  assign t_r13_c34_2 = p_13_34 << 2;
  assign t_r13_c34_3 = p_13_35 << 1;
  assign t_r13_c34_4 = p_14_34 << 1;
  assign t_r13_c34_5 = t_r13_c34_0 + p_12_33;
  assign t_r13_c34_6 = t_r13_c34_1 + p_12_35;
  assign t_r13_c34_7 = t_r13_c34_2 + t_r13_c34_3;
  assign t_r13_c34_8 = t_r13_c34_4 + p_14_33;
  assign t_r13_c34_9 = t_r13_c34_5 + t_r13_c34_6;
  assign t_r13_c34_10 = t_r13_c34_7 + t_r13_c34_8;
  assign t_r13_c34_11 = t_r13_c34_9 + t_r13_c34_10;
  assign t_r13_c34_12 = t_r13_c34_11 + p_14_35;
  assign out_13_34 = t_r13_c34_12 >> 4;

  assign t_r13_c35_0 = p_12_35 << 1;
  assign t_r13_c35_1 = p_13_34 << 1;
  assign t_r13_c35_2 = p_13_35 << 2;
  assign t_r13_c35_3 = p_13_36 << 1;
  assign t_r13_c35_4 = p_14_35 << 1;
  assign t_r13_c35_5 = t_r13_c35_0 + p_12_34;
  assign t_r13_c35_6 = t_r13_c35_1 + p_12_36;
  assign t_r13_c35_7 = t_r13_c35_2 + t_r13_c35_3;
  assign t_r13_c35_8 = t_r13_c35_4 + p_14_34;
  assign t_r13_c35_9 = t_r13_c35_5 + t_r13_c35_6;
  assign t_r13_c35_10 = t_r13_c35_7 + t_r13_c35_8;
  assign t_r13_c35_11 = t_r13_c35_9 + t_r13_c35_10;
  assign t_r13_c35_12 = t_r13_c35_11 + p_14_36;
  assign out_13_35 = t_r13_c35_12 >> 4;

  assign t_r13_c36_0 = p_12_36 << 1;
  assign t_r13_c36_1 = p_13_35 << 1;
  assign t_r13_c36_2 = p_13_36 << 2;
  assign t_r13_c36_3 = p_13_37 << 1;
  assign t_r13_c36_4 = p_14_36 << 1;
  assign t_r13_c36_5 = t_r13_c36_0 + p_12_35;
  assign t_r13_c36_6 = t_r13_c36_1 + p_12_37;
  assign t_r13_c36_7 = t_r13_c36_2 + t_r13_c36_3;
  assign t_r13_c36_8 = t_r13_c36_4 + p_14_35;
  assign t_r13_c36_9 = t_r13_c36_5 + t_r13_c36_6;
  assign t_r13_c36_10 = t_r13_c36_7 + t_r13_c36_8;
  assign t_r13_c36_11 = t_r13_c36_9 + t_r13_c36_10;
  assign t_r13_c36_12 = t_r13_c36_11 + p_14_37;
  assign out_13_36 = t_r13_c36_12 >> 4;

  assign t_r13_c37_0 = p_12_37 << 1;
  assign t_r13_c37_1 = p_13_36 << 1;
  assign t_r13_c37_2 = p_13_37 << 2;
  assign t_r13_c37_3 = p_13_38 << 1;
  assign t_r13_c37_4 = p_14_37 << 1;
  assign t_r13_c37_5 = t_r13_c37_0 + p_12_36;
  assign t_r13_c37_6 = t_r13_c37_1 + p_12_38;
  assign t_r13_c37_7 = t_r13_c37_2 + t_r13_c37_3;
  assign t_r13_c37_8 = t_r13_c37_4 + p_14_36;
  assign t_r13_c37_9 = t_r13_c37_5 + t_r13_c37_6;
  assign t_r13_c37_10 = t_r13_c37_7 + t_r13_c37_8;
  assign t_r13_c37_11 = t_r13_c37_9 + t_r13_c37_10;
  assign t_r13_c37_12 = t_r13_c37_11 + p_14_38;
  assign out_13_37 = t_r13_c37_12 >> 4;

  assign t_r13_c38_0 = p_12_38 << 1;
  assign t_r13_c38_1 = p_13_37 << 1;
  assign t_r13_c38_2 = p_13_38 << 2;
  assign t_r13_c38_3 = p_13_39 << 1;
  assign t_r13_c38_4 = p_14_38 << 1;
  assign t_r13_c38_5 = t_r13_c38_0 + p_12_37;
  assign t_r13_c38_6 = t_r13_c38_1 + p_12_39;
  assign t_r13_c38_7 = t_r13_c38_2 + t_r13_c38_3;
  assign t_r13_c38_8 = t_r13_c38_4 + p_14_37;
  assign t_r13_c38_9 = t_r13_c38_5 + t_r13_c38_6;
  assign t_r13_c38_10 = t_r13_c38_7 + t_r13_c38_8;
  assign t_r13_c38_11 = t_r13_c38_9 + t_r13_c38_10;
  assign t_r13_c38_12 = t_r13_c38_11 + p_14_39;
  assign out_13_38 = t_r13_c38_12 >> 4;

  assign t_r13_c39_0 = p_12_39 << 1;
  assign t_r13_c39_1 = p_13_38 << 1;
  assign t_r13_c39_2 = p_13_39 << 2;
  assign t_r13_c39_3 = p_13_40 << 1;
  assign t_r13_c39_4 = p_14_39 << 1;
  assign t_r13_c39_5 = t_r13_c39_0 + p_12_38;
  assign t_r13_c39_6 = t_r13_c39_1 + p_12_40;
  assign t_r13_c39_7 = t_r13_c39_2 + t_r13_c39_3;
  assign t_r13_c39_8 = t_r13_c39_4 + p_14_38;
  assign t_r13_c39_9 = t_r13_c39_5 + t_r13_c39_6;
  assign t_r13_c39_10 = t_r13_c39_7 + t_r13_c39_8;
  assign t_r13_c39_11 = t_r13_c39_9 + t_r13_c39_10;
  assign t_r13_c39_12 = t_r13_c39_11 + p_14_40;
  assign out_13_39 = t_r13_c39_12 >> 4;

  assign t_r13_c40_0 = p_12_40 << 1;
  assign t_r13_c40_1 = p_13_39 << 1;
  assign t_r13_c40_2 = p_13_40 << 2;
  assign t_r13_c40_3 = p_13_41 << 1;
  assign t_r13_c40_4 = p_14_40 << 1;
  assign t_r13_c40_5 = t_r13_c40_0 + p_12_39;
  assign t_r13_c40_6 = t_r13_c40_1 + p_12_41;
  assign t_r13_c40_7 = t_r13_c40_2 + t_r13_c40_3;
  assign t_r13_c40_8 = t_r13_c40_4 + p_14_39;
  assign t_r13_c40_9 = t_r13_c40_5 + t_r13_c40_6;
  assign t_r13_c40_10 = t_r13_c40_7 + t_r13_c40_8;
  assign t_r13_c40_11 = t_r13_c40_9 + t_r13_c40_10;
  assign t_r13_c40_12 = t_r13_c40_11 + p_14_41;
  assign out_13_40 = t_r13_c40_12 >> 4;

  assign t_r13_c41_0 = p_12_41 << 1;
  assign t_r13_c41_1 = p_13_40 << 1;
  assign t_r13_c41_2 = p_13_41 << 2;
  assign t_r13_c41_3 = p_13_42 << 1;
  assign t_r13_c41_4 = p_14_41 << 1;
  assign t_r13_c41_5 = t_r13_c41_0 + p_12_40;
  assign t_r13_c41_6 = t_r13_c41_1 + p_12_42;
  assign t_r13_c41_7 = t_r13_c41_2 + t_r13_c41_3;
  assign t_r13_c41_8 = t_r13_c41_4 + p_14_40;
  assign t_r13_c41_9 = t_r13_c41_5 + t_r13_c41_6;
  assign t_r13_c41_10 = t_r13_c41_7 + t_r13_c41_8;
  assign t_r13_c41_11 = t_r13_c41_9 + t_r13_c41_10;
  assign t_r13_c41_12 = t_r13_c41_11 + p_14_42;
  assign out_13_41 = t_r13_c41_12 >> 4;

  assign t_r13_c42_0 = p_12_42 << 1;
  assign t_r13_c42_1 = p_13_41 << 1;
  assign t_r13_c42_2 = p_13_42 << 2;
  assign t_r13_c42_3 = p_13_43 << 1;
  assign t_r13_c42_4 = p_14_42 << 1;
  assign t_r13_c42_5 = t_r13_c42_0 + p_12_41;
  assign t_r13_c42_6 = t_r13_c42_1 + p_12_43;
  assign t_r13_c42_7 = t_r13_c42_2 + t_r13_c42_3;
  assign t_r13_c42_8 = t_r13_c42_4 + p_14_41;
  assign t_r13_c42_9 = t_r13_c42_5 + t_r13_c42_6;
  assign t_r13_c42_10 = t_r13_c42_7 + t_r13_c42_8;
  assign t_r13_c42_11 = t_r13_c42_9 + t_r13_c42_10;
  assign t_r13_c42_12 = t_r13_c42_11 + p_14_43;
  assign out_13_42 = t_r13_c42_12 >> 4;

  assign t_r13_c43_0 = p_12_43 << 1;
  assign t_r13_c43_1 = p_13_42 << 1;
  assign t_r13_c43_2 = p_13_43 << 2;
  assign t_r13_c43_3 = p_13_44 << 1;
  assign t_r13_c43_4 = p_14_43 << 1;
  assign t_r13_c43_5 = t_r13_c43_0 + p_12_42;
  assign t_r13_c43_6 = t_r13_c43_1 + p_12_44;
  assign t_r13_c43_7 = t_r13_c43_2 + t_r13_c43_3;
  assign t_r13_c43_8 = t_r13_c43_4 + p_14_42;
  assign t_r13_c43_9 = t_r13_c43_5 + t_r13_c43_6;
  assign t_r13_c43_10 = t_r13_c43_7 + t_r13_c43_8;
  assign t_r13_c43_11 = t_r13_c43_9 + t_r13_c43_10;
  assign t_r13_c43_12 = t_r13_c43_11 + p_14_44;
  assign out_13_43 = t_r13_c43_12 >> 4;

  assign t_r13_c44_0 = p_12_44 << 1;
  assign t_r13_c44_1 = p_13_43 << 1;
  assign t_r13_c44_2 = p_13_44 << 2;
  assign t_r13_c44_3 = p_13_45 << 1;
  assign t_r13_c44_4 = p_14_44 << 1;
  assign t_r13_c44_5 = t_r13_c44_0 + p_12_43;
  assign t_r13_c44_6 = t_r13_c44_1 + p_12_45;
  assign t_r13_c44_7 = t_r13_c44_2 + t_r13_c44_3;
  assign t_r13_c44_8 = t_r13_c44_4 + p_14_43;
  assign t_r13_c44_9 = t_r13_c44_5 + t_r13_c44_6;
  assign t_r13_c44_10 = t_r13_c44_7 + t_r13_c44_8;
  assign t_r13_c44_11 = t_r13_c44_9 + t_r13_c44_10;
  assign t_r13_c44_12 = t_r13_c44_11 + p_14_45;
  assign out_13_44 = t_r13_c44_12 >> 4;

  assign t_r13_c45_0 = p_12_45 << 1;
  assign t_r13_c45_1 = p_13_44 << 1;
  assign t_r13_c45_2 = p_13_45 << 2;
  assign t_r13_c45_3 = p_13_46 << 1;
  assign t_r13_c45_4 = p_14_45 << 1;
  assign t_r13_c45_5 = t_r13_c45_0 + p_12_44;
  assign t_r13_c45_6 = t_r13_c45_1 + p_12_46;
  assign t_r13_c45_7 = t_r13_c45_2 + t_r13_c45_3;
  assign t_r13_c45_8 = t_r13_c45_4 + p_14_44;
  assign t_r13_c45_9 = t_r13_c45_5 + t_r13_c45_6;
  assign t_r13_c45_10 = t_r13_c45_7 + t_r13_c45_8;
  assign t_r13_c45_11 = t_r13_c45_9 + t_r13_c45_10;
  assign t_r13_c45_12 = t_r13_c45_11 + p_14_46;
  assign out_13_45 = t_r13_c45_12 >> 4;

  assign t_r13_c46_0 = p_12_46 << 1;
  assign t_r13_c46_1 = p_13_45 << 1;
  assign t_r13_c46_2 = p_13_46 << 2;
  assign t_r13_c46_3 = p_13_47 << 1;
  assign t_r13_c46_4 = p_14_46 << 1;
  assign t_r13_c46_5 = t_r13_c46_0 + p_12_45;
  assign t_r13_c46_6 = t_r13_c46_1 + p_12_47;
  assign t_r13_c46_7 = t_r13_c46_2 + t_r13_c46_3;
  assign t_r13_c46_8 = t_r13_c46_4 + p_14_45;
  assign t_r13_c46_9 = t_r13_c46_5 + t_r13_c46_6;
  assign t_r13_c46_10 = t_r13_c46_7 + t_r13_c46_8;
  assign t_r13_c46_11 = t_r13_c46_9 + t_r13_c46_10;
  assign t_r13_c46_12 = t_r13_c46_11 + p_14_47;
  assign out_13_46 = t_r13_c46_12 >> 4;

  assign t_r13_c47_0 = p_12_47 << 1;
  assign t_r13_c47_1 = p_13_46 << 1;
  assign t_r13_c47_2 = p_13_47 << 2;
  assign t_r13_c47_3 = p_13_48 << 1;
  assign t_r13_c47_4 = p_14_47 << 1;
  assign t_r13_c47_5 = t_r13_c47_0 + p_12_46;
  assign t_r13_c47_6 = t_r13_c47_1 + p_12_48;
  assign t_r13_c47_7 = t_r13_c47_2 + t_r13_c47_3;
  assign t_r13_c47_8 = t_r13_c47_4 + p_14_46;
  assign t_r13_c47_9 = t_r13_c47_5 + t_r13_c47_6;
  assign t_r13_c47_10 = t_r13_c47_7 + t_r13_c47_8;
  assign t_r13_c47_11 = t_r13_c47_9 + t_r13_c47_10;
  assign t_r13_c47_12 = t_r13_c47_11 + p_14_48;
  assign out_13_47 = t_r13_c47_12 >> 4;

  assign t_r13_c48_0 = p_12_48 << 1;
  assign t_r13_c48_1 = p_13_47 << 1;
  assign t_r13_c48_2 = p_13_48 << 2;
  assign t_r13_c48_3 = p_13_49 << 1;
  assign t_r13_c48_4 = p_14_48 << 1;
  assign t_r13_c48_5 = t_r13_c48_0 + p_12_47;
  assign t_r13_c48_6 = t_r13_c48_1 + p_12_49;
  assign t_r13_c48_7 = t_r13_c48_2 + t_r13_c48_3;
  assign t_r13_c48_8 = t_r13_c48_4 + p_14_47;
  assign t_r13_c48_9 = t_r13_c48_5 + t_r13_c48_6;
  assign t_r13_c48_10 = t_r13_c48_7 + t_r13_c48_8;
  assign t_r13_c48_11 = t_r13_c48_9 + t_r13_c48_10;
  assign t_r13_c48_12 = t_r13_c48_11 + p_14_49;
  assign out_13_48 = t_r13_c48_12 >> 4;

  assign t_r13_c49_0 = p_12_49 << 1;
  assign t_r13_c49_1 = p_13_48 << 1;
  assign t_r13_c49_2 = p_13_49 << 2;
  assign t_r13_c49_3 = p_13_50 << 1;
  assign t_r13_c49_4 = p_14_49 << 1;
  assign t_r13_c49_5 = t_r13_c49_0 + p_12_48;
  assign t_r13_c49_6 = t_r13_c49_1 + p_12_50;
  assign t_r13_c49_7 = t_r13_c49_2 + t_r13_c49_3;
  assign t_r13_c49_8 = t_r13_c49_4 + p_14_48;
  assign t_r13_c49_9 = t_r13_c49_5 + t_r13_c49_6;
  assign t_r13_c49_10 = t_r13_c49_7 + t_r13_c49_8;
  assign t_r13_c49_11 = t_r13_c49_9 + t_r13_c49_10;
  assign t_r13_c49_12 = t_r13_c49_11 + p_14_50;
  assign out_13_49 = t_r13_c49_12 >> 4;

  assign t_r13_c50_0 = p_12_50 << 1;
  assign t_r13_c50_1 = p_13_49 << 1;
  assign t_r13_c50_2 = p_13_50 << 2;
  assign t_r13_c50_3 = p_13_51 << 1;
  assign t_r13_c50_4 = p_14_50 << 1;
  assign t_r13_c50_5 = t_r13_c50_0 + p_12_49;
  assign t_r13_c50_6 = t_r13_c50_1 + p_12_51;
  assign t_r13_c50_7 = t_r13_c50_2 + t_r13_c50_3;
  assign t_r13_c50_8 = t_r13_c50_4 + p_14_49;
  assign t_r13_c50_9 = t_r13_c50_5 + t_r13_c50_6;
  assign t_r13_c50_10 = t_r13_c50_7 + t_r13_c50_8;
  assign t_r13_c50_11 = t_r13_c50_9 + t_r13_c50_10;
  assign t_r13_c50_12 = t_r13_c50_11 + p_14_51;
  assign out_13_50 = t_r13_c50_12 >> 4;

  assign t_r13_c51_0 = p_12_51 << 1;
  assign t_r13_c51_1 = p_13_50 << 1;
  assign t_r13_c51_2 = p_13_51 << 2;
  assign t_r13_c51_3 = p_13_52 << 1;
  assign t_r13_c51_4 = p_14_51 << 1;
  assign t_r13_c51_5 = t_r13_c51_0 + p_12_50;
  assign t_r13_c51_6 = t_r13_c51_1 + p_12_52;
  assign t_r13_c51_7 = t_r13_c51_2 + t_r13_c51_3;
  assign t_r13_c51_8 = t_r13_c51_4 + p_14_50;
  assign t_r13_c51_9 = t_r13_c51_5 + t_r13_c51_6;
  assign t_r13_c51_10 = t_r13_c51_7 + t_r13_c51_8;
  assign t_r13_c51_11 = t_r13_c51_9 + t_r13_c51_10;
  assign t_r13_c51_12 = t_r13_c51_11 + p_14_52;
  assign out_13_51 = t_r13_c51_12 >> 4;

  assign t_r13_c52_0 = p_12_52 << 1;
  assign t_r13_c52_1 = p_13_51 << 1;
  assign t_r13_c52_2 = p_13_52 << 2;
  assign t_r13_c52_3 = p_13_53 << 1;
  assign t_r13_c52_4 = p_14_52 << 1;
  assign t_r13_c52_5 = t_r13_c52_0 + p_12_51;
  assign t_r13_c52_6 = t_r13_c52_1 + p_12_53;
  assign t_r13_c52_7 = t_r13_c52_2 + t_r13_c52_3;
  assign t_r13_c52_8 = t_r13_c52_4 + p_14_51;
  assign t_r13_c52_9 = t_r13_c52_5 + t_r13_c52_6;
  assign t_r13_c52_10 = t_r13_c52_7 + t_r13_c52_8;
  assign t_r13_c52_11 = t_r13_c52_9 + t_r13_c52_10;
  assign t_r13_c52_12 = t_r13_c52_11 + p_14_53;
  assign out_13_52 = t_r13_c52_12 >> 4;

  assign t_r13_c53_0 = p_12_53 << 1;
  assign t_r13_c53_1 = p_13_52 << 1;
  assign t_r13_c53_2 = p_13_53 << 2;
  assign t_r13_c53_3 = p_13_54 << 1;
  assign t_r13_c53_4 = p_14_53 << 1;
  assign t_r13_c53_5 = t_r13_c53_0 + p_12_52;
  assign t_r13_c53_6 = t_r13_c53_1 + p_12_54;
  assign t_r13_c53_7 = t_r13_c53_2 + t_r13_c53_3;
  assign t_r13_c53_8 = t_r13_c53_4 + p_14_52;
  assign t_r13_c53_9 = t_r13_c53_5 + t_r13_c53_6;
  assign t_r13_c53_10 = t_r13_c53_7 + t_r13_c53_8;
  assign t_r13_c53_11 = t_r13_c53_9 + t_r13_c53_10;
  assign t_r13_c53_12 = t_r13_c53_11 + p_14_54;
  assign out_13_53 = t_r13_c53_12 >> 4;

  assign t_r13_c54_0 = p_12_54 << 1;
  assign t_r13_c54_1 = p_13_53 << 1;
  assign t_r13_c54_2 = p_13_54 << 2;
  assign t_r13_c54_3 = p_13_55 << 1;
  assign t_r13_c54_4 = p_14_54 << 1;
  assign t_r13_c54_5 = t_r13_c54_0 + p_12_53;
  assign t_r13_c54_6 = t_r13_c54_1 + p_12_55;
  assign t_r13_c54_7 = t_r13_c54_2 + t_r13_c54_3;
  assign t_r13_c54_8 = t_r13_c54_4 + p_14_53;
  assign t_r13_c54_9 = t_r13_c54_5 + t_r13_c54_6;
  assign t_r13_c54_10 = t_r13_c54_7 + t_r13_c54_8;
  assign t_r13_c54_11 = t_r13_c54_9 + t_r13_c54_10;
  assign t_r13_c54_12 = t_r13_c54_11 + p_14_55;
  assign out_13_54 = t_r13_c54_12 >> 4;

  assign t_r13_c55_0 = p_12_55 << 1;
  assign t_r13_c55_1 = p_13_54 << 1;
  assign t_r13_c55_2 = p_13_55 << 2;
  assign t_r13_c55_3 = p_13_56 << 1;
  assign t_r13_c55_4 = p_14_55 << 1;
  assign t_r13_c55_5 = t_r13_c55_0 + p_12_54;
  assign t_r13_c55_6 = t_r13_c55_1 + p_12_56;
  assign t_r13_c55_7 = t_r13_c55_2 + t_r13_c55_3;
  assign t_r13_c55_8 = t_r13_c55_4 + p_14_54;
  assign t_r13_c55_9 = t_r13_c55_5 + t_r13_c55_6;
  assign t_r13_c55_10 = t_r13_c55_7 + t_r13_c55_8;
  assign t_r13_c55_11 = t_r13_c55_9 + t_r13_c55_10;
  assign t_r13_c55_12 = t_r13_c55_11 + p_14_56;
  assign out_13_55 = t_r13_c55_12 >> 4;

  assign t_r13_c56_0 = p_12_56 << 1;
  assign t_r13_c56_1 = p_13_55 << 1;
  assign t_r13_c56_2 = p_13_56 << 2;
  assign t_r13_c56_3 = p_13_57 << 1;
  assign t_r13_c56_4 = p_14_56 << 1;
  assign t_r13_c56_5 = t_r13_c56_0 + p_12_55;
  assign t_r13_c56_6 = t_r13_c56_1 + p_12_57;
  assign t_r13_c56_7 = t_r13_c56_2 + t_r13_c56_3;
  assign t_r13_c56_8 = t_r13_c56_4 + p_14_55;
  assign t_r13_c56_9 = t_r13_c56_5 + t_r13_c56_6;
  assign t_r13_c56_10 = t_r13_c56_7 + t_r13_c56_8;
  assign t_r13_c56_11 = t_r13_c56_9 + t_r13_c56_10;
  assign t_r13_c56_12 = t_r13_c56_11 + p_14_57;
  assign out_13_56 = t_r13_c56_12 >> 4;

  assign t_r13_c57_0 = p_12_57 << 1;
  assign t_r13_c57_1 = p_13_56 << 1;
  assign t_r13_c57_2 = p_13_57 << 2;
  assign t_r13_c57_3 = p_13_58 << 1;
  assign t_r13_c57_4 = p_14_57 << 1;
  assign t_r13_c57_5 = t_r13_c57_0 + p_12_56;
  assign t_r13_c57_6 = t_r13_c57_1 + p_12_58;
  assign t_r13_c57_7 = t_r13_c57_2 + t_r13_c57_3;
  assign t_r13_c57_8 = t_r13_c57_4 + p_14_56;
  assign t_r13_c57_9 = t_r13_c57_5 + t_r13_c57_6;
  assign t_r13_c57_10 = t_r13_c57_7 + t_r13_c57_8;
  assign t_r13_c57_11 = t_r13_c57_9 + t_r13_c57_10;
  assign t_r13_c57_12 = t_r13_c57_11 + p_14_58;
  assign out_13_57 = t_r13_c57_12 >> 4;

  assign t_r13_c58_0 = p_12_58 << 1;
  assign t_r13_c58_1 = p_13_57 << 1;
  assign t_r13_c58_2 = p_13_58 << 2;
  assign t_r13_c58_3 = p_13_59 << 1;
  assign t_r13_c58_4 = p_14_58 << 1;
  assign t_r13_c58_5 = t_r13_c58_0 + p_12_57;
  assign t_r13_c58_6 = t_r13_c58_1 + p_12_59;
  assign t_r13_c58_7 = t_r13_c58_2 + t_r13_c58_3;
  assign t_r13_c58_8 = t_r13_c58_4 + p_14_57;
  assign t_r13_c58_9 = t_r13_c58_5 + t_r13_c58_6;
  assign t_r13_c58_10 = t_r13_c58_7 + t_r13_c58_8;
  assign t_r13_c58_11 = t_r13_c58_9 + t_r13_c58_10;
  assign t_r13_c58_12 = t_r13_c58_11 + p_14_59;
  assign out_13_58 = t_r13_c58_12 >> 4;

  assign t_r13_c59_0 = p_12_59 << 1;
  assign t_r13_c59_1 = p_13_58 << 1;
  assign t_r13_c59_2 = p_13_59 << 2;
  assign t_r13_c59_3 = p_13_60 << 1;
  assign t_r13_c59_4 = p_14_59 << 1;
  assign t_r13_c59_5 = t_r13_c59_0 + p_12_58;
  assign t_r13_c59_6 = t_r13_c59_1 + p_12_60;
  assign t_r13_c59_7 = t_r13_c59_2 + t_r13_c59_3;
  assign t_r13_c59_8 = t_r13_c59_4 + p_14_58;
  assign t_r13_c59_9 = t_r13_c59_5 + t_r13_c59_6;
  assign t_r13_c59_10 = t_r13_c59_7 + t_r13_c59_8;
  assign t_r13_c59_11 = t_r13_c59_9 + t_r13_c59_10;
  assign t_r13_c59_12 = t_r13_c59_11 + p_14_60;
  assign out_13_59 = t_r13_c59_12 >> 4;

  assign t_r13_c60_0 = p_12_60 << 1;
  assign t_r13_c60_1 = p_13_59 << 1;
  assign t_r13_c60_2 = p_13_60 << 2;
  assign t_r13_c60_3 = p_13_61 << 1;
  assign t_r13_c60_4 = p_14_60 << 1;
  assign t_r13_c60_5 = t_r13_c60_0 + p_12_59;
  assign t_r13_c60_6 = t_r13_c60_1 + p_12_61;
  assign t_r13_c60_7 = t_r13_c60_2 + t_r13_c60_3;
  assign t_r13_c60_8 = t_r13_c60_4 + p_14_59;
  assign t_r13_c60_9 = t_r13_c60_5 + t_r13_c60_6;
  assign t_r13_c60_10 = t_r13_c60_7 + t_r13_c60_8;
  assign t_r13_c60_11 = t_r13_c60_9 + t_r13_c60_10;
  assign t_r13_c60_12 = t_r13_c60_11 + p_14_61;
  assign out_13_60 = t_r13_c60_12 >> 4;

  assign t_r13_c61_0 = p_12_61 << 1;
  assign t_r13_c61_1 = p_13_60 << 1;
  assign t_r13_c61_2 = p_13_61 << 2;
  assign t_r13_c61_3 = p_13_62 << 1;
  assign t_r13_c61_4 = p_14_61 << 1;
  assign t_r13_c61_5 = t_r13_c61_0 + p_12_60;
  assign t_r13_c61_6 = t_r13_c61_1 + p_12_62;
  assign t_r13_c61_7 = t_r13_c61_2 + t_r13_c61_3;
  assign t_r13_c61_8 = t_r13_c61_4 + p_14_60;
  assign t_r13_c61_9 = t_r13_c61_5 + t_r13_c61_6;
  assign t_r13_c61_10 = t_r13_c61_7 + t_r13_c61_8;
  assign t_r13_c61_11 = t_r13_c61_9 + t_r13_c61_10;
  assign t_r13_c61_12 = t_r13_c61_11 + p_14_62;
  assign out_13_61 = t_r13_c61_12 >> 4;

  assign t_r13_c62_0 = p_12_62 << 1;
  assign t_r13_c62_1 = p_13_61 << 1;
  assign t_r13_c62_2 = p_13_62 << 2;
  assign t_r13_c62_3 = p_13_63 << 1;
  assign t_r13_c62_4 = p_14_62 << 1;
  assign t_r13_c62_5 = t_r13_c62_0 + p_12_61;
  assign t_r13_c62_6 = t_r13_c62_1 + p_12_63;
  assign t_r13_c62_7 = t_r13_c62_2 + t_r13_c62_3;
  assign t_r13_c62_8 = t_r13_c62_4 + p_14_61;
  assign t_r13_c62_9 = t_r13_c62_5 + t_r13_c62_6;
  assign t_r13_c62_10 = t_r13_c62_7 + t_r13_c62_8;
  assign t_r13_c62_11 = t_r13_c62_9 + t_r13_c62_10;
  assign t_r13_c62_12 = t_r13_c62_11 + p_14_63;
  assign out_13_62 = t_r13_c62_12 >> 4;

  assign t_r13_c63_0 = p_12_63 << 1;
  assign t_r13_c63_1 = p_13_62 << 1;
  assign t_r13_c63_2 = p_13_63 << 2;
  assign t_r13_c63_3 = p_13_64 << 1;
  assign t_r13_c63_4 = p_14_63 << 1;
  assign t_r13_c63_5 = t_r13_c63_0 + p_12_62;
  assign t_r13_c63_6 = t_r13_c63_1 + p_12_64;
  assign t_r13_c63_7 = t_r13_c63_2 + t_r13_c63_3;
  assign t_r13_c63_8 = t_r13_c63_4 + p_14_62;
  assign t_r13_c63_9 = t_r13_c63_5 + t_r13_c63_6;
  assign t_r13_c63_10 = t_r13_c63_7 + t_r13_c63_8;
  assign t_r13_c63_11 = t_r13_c63_9 + t_r13_c63_10;
  assign t_r13_c63_12 = t_r13_c63_11 + p_14_64;
  assign out_13_63 = t_r13_c63_12 >> 4;

  assign t_r13_c64_0 = p_12_64 << 1;
  assign t_r13_c64_1 = p_13_63 << 1;
  assign t_r13_c64_2 = p_13_64 << 2;
  assign t_r13_c64_3 = p_13_65 << 1;
  assign t_r13_c64_4 = p_14_64 << 1;
  assign t_r13_c64_5 = t_r13_c64_0 + p_12_63;
  assign t_r13_c64_6 = t_r13_c64_1 + p_12_65;
  assign t_r13_c64_7 = t_r13_c64_2 + t_r13_c64_3;
  assign t_r13_c64_8 = t_r13_c64_4 + p_14_63;
  assign t_r13_c64_9 = t_r13_c64_5 + t_r13_c64_6;
  assign t_r13_c64_10 = t_r13_c64_7 + t_r13_c64_8;
  assign t_r13_c64_11 = t_r13_c64_9 + t_r13_c64_10;
  assign t_r13_c64_12 = t_r13_c64_11 + p_14_65;
  assign out_13_64 = t_r13_c64_12 >> 4;

  assign t_r14_c1_0 = p_13_1 << 1;
  assign t_r14_c1_1 = p_14_0 << 1;
  assign t_r14_c1_2 = p_14_1 << 2;
  assign t_r14_c1_3 = p_14_2 << 1;
  assign t_r14_c1_4 = p_15_1 << 1;
  assign t_r14_c1_5 = t_r14_c1_0 + p_13_0;
  assign t_r14_c1_6 = t_r14_c1_1 + p_13_2;
  assign t_r14_c1_7 = t_r14_c1_2 + t_r14_c1_3;
  assign t_r14_c1_8 = t_r14_c1_4 + p_15_0;
  assign t_r14_c1_9 = t_r14_c1_5 + t_r14_c1_6;
  assign t_r14_c1_10 = t_r14_c1_7 + t_r14_c1_8;
  assign t_r14_c1_11 = t_r14_c1_9 + t_r14_c1_10;
  assign t_r14_c1_12 = t_r14_c1_11 + p_15_2;
  assign out_14_1 = t_r14_c1_12 >> 4;

  assign t_r14_c2_0 = p_13_2 << 1;
  assign t_r14_c2_1 = p_14_1 << 1;
  assign t_r14_c2_2 = p_14_2 << 2;
  assign t_r14_c2_3 = p_14_3 << 1;
  assign t_r14_c2_4 = p_15_2 << 1;
  assign t_r14_c2_5 = t_r14_c2_0 + p_13_1;
  assign t_r14_c2_6 = t_r14_c2_1 + p_13_3;
  assign t_r14_c2_7 = t_r14_c2_2 + t_r14_c2_3;
  assign t_r14_c2_8 = t_r14_c2_4 + p_15_1;
  assign t_r14_c2_9 = t_r14_c2_5 + t_r14_c2_6;
  assign t_r14_c2_10 = t_r14_c2_7 + t_r14_c2_8;
  assign t_r14_c2_11 = t_r14_c2_9 + t_r14_c2_10;
  assign t_r14_c2_12 = t_r14_c2_11 + p_15_3;
  assign out_14_2 = t_r14_c2_12 >> 4;

  assign t_r14_c3_0 = p_13_3 << 1;
  assign t_r14_c3_1 = p_14_2 << 1;
  assign t_r14_c3_2 = p_14_3 << 2;
  assign t_r14_c3_3 = p_14_4 << 1;
  assign t_r14_c3_4 = p_15_3 << 1;
  assign t_r14_c3_5 = t_r14_c3_0 + p_13_2;
  assign t_r14_c3_6 = t_r14_c3_1 + p_13_4;
  assign t_r14_c3_7 = t_r14_c3_2 + t_r14_c3_3;
  assign t_r14_c3_8 = t_r14_c3_4 + p_15_2;
  assign t_r14_c3_9 = t_r14_c3_5 + t_r14_c3_6;
  assign t_r14_c3_10 = t_r14_c3_7 + t_r14_c3_8;
  assign t_r14_c3_11 = t_r14_c3_9 + t_r14_c3_10;
  assign t_r14_c3_12 = t_r14_c3_11 + p_15_4;
  assign out_14_3 = t_r14_c3_12 >> 4;

  assign t_r14_c4_0 = p_13_4 << 1;
  assign t_r14_c4_1 = p_14_3 << 1;
  assign t_r14_c4_2 = p_14_4 << 2;
  assign t_r14_c4_3 = p_14_5 << 1;
  assign t_r14_c4_4 = p_15_4 << 1;
  assign t_r14_c4_5 = t_r14_c4_0 + p_13_3;
  assign t_r14_c4_6 = t_r14_c4_1 + p_13_5;
  assign t_r14_c4_7 = t_r14_c4_2 + t_r14_c4_3;
  assign t_r14_c4_8 = t_r14_c4_4 + p_15_3;
  assign t_r14_c4_9 = t_r14_c4_5 + t_r14_c4_6;
  assign t_r14_c4_10 = t_r14_c4_7 + t_r14_c4_8;
  assign t_r14_c4_11 = t_r14_c4_9 + t_r14_c4_10;
  assign t_r14_c4_12 = t_r14_c4_11 + p_15_5;
  assign out_14_4 = t_r14_c4_12 >> 4;

  assign t_r14_c5_0 = p_13_5 << 1;
  assign t_r14_c5_1 = p_14_4 << 1;
  assign t_r14_c5_2 = p_14_5 << 2;
  assign t_r14_c5_3 = p_14_6 << 1;
  assign t_r14_c5_4 = p_15_5 << 1;
  assign t_r14_c5_5 = t_r14_c5_0 + p_13_4;
  assign t_r14_c5_6 = t_r14_c5_1 + p_13_6;
  assign t_r14_c5_7 = t_r14_c5_2 + t_r14_c5_3;
  assign t_r14_c5_8 = t_r14_c5_4 + p_15_4;
  assign t_r14_c5_9 = t_r14_c5_5 + t_r14_c5_6;
  assign t_r14_c5_10 = t_r14_c5_7 + t_r14_c5_8;
  assign t_r14_c5_11 = t_r14_c5_9 + t_r14_c5_10;
  assign t_r14_c5_12 = t_r14_c5_11 + p_15_6;
  assign out_14_5 = t_r14_c5_12 >> 4;

  assign t_r14_c6_0 = p_13_6 << 1;
  assign t_r14_c6_1 = p_14_5 << 1;
  assign t_r14_c6_2 = p_14_6 << 2;
  assign t_r14_c6_3 = p_14_7 << 1;
  assign t_r14_c6_4 = p_15_6 << 1;
  assign t_r14_c6_5 = t_r14_c6_0 + p_13_5;
  assign t_r14_c6_6 = t_r14_c6_1 + p_13_7;
  assign t_r14_c6_7 = t_r14_c6_2 + t_r14_c6_3;
  assign t_r14_c6_8 = t_r14_c6_4 + p_15_5;
  assign t_r14_c6_9 = t_r14_c6_5 + t_r14_c6_6;
  assign t_r14_c6_10 = t_r14_c6_7 + t_r14_c6_8;
  assign t_r14_c6_11 = t_r14_c6_9 + t_r14_c6_10;
  assign t_r14_c6_12 = t_r14_c6_11 + p_15_7;
  assign out_14_6 = t_r14_c6_12 >> 4;

  assign t_r14_c7_0 = p_13_7 << 1;
  assign t_r14_c7_1 = p_14_6 << 1;
  assign t_r14_c7_2 = p_14_7 << 2;
  assign t_r14_c7_3 = p_14_8 << 1;
  assign t_r14_c7_4 = p_15_7 << 1;
  assign t_r14_c7_5 = t_r14_c7_0 + p_13_6;
  assign t_r14_c7_6 = t_r14_c7_1 + p_13_8;
  assign t_r14_c7_7 = t_r14_c7_2 + t_r14_c7_3;
  assign t_r14_c7_8 = t_r14_c7_4 + p_15_6;
  assign t_r14_c7_9 = t_r14_c7_5 + t_r14_c7_6;
  assign t_r14_c7_10 = t_r14_c7_7 + t_r14_c7_8;
  assign t_r14_c7_11 = t_r14_c7_9 + t_r14_c7_10;
  assign t_r14_c7_12 = t_r14_c7_11 + p_15_8;
  assign out_14_7 = t_r14_c7_12 >> 4;

  assign t_r14_c8_0 = p_13_8 << 1;
  assign t_r14_c8_1 = p_14_7 << 1;
  assign t_r14_c8_2 = p_14_8 << 2;
  assign t_r14_c8_3 = p_14_9 << 1;
  assign t_r14_c8_4 = p_15_8 << 1;
  assign t_r14_c8_5 = t_r14_c8_0 + p_13_7;
  assign t_r14_c8_6 = t_r14_c8_1 + p_13_9;
  assign t_r14_c8_7 = t_r14_c8_2 + t_r14_c8_3;
  assign t_r14_c8_8 = t_r14_c8_4 + p_15_7;
  assign t_r14_c8_9 = t_r14_c8_5 + t_r14_c8_6;
  assign t_r14_c8_10 = t_r14_c8_7 + t_r14_c8_8;
  assign t_r14_c8_11 = t_r14_c8_9 + t_r14_c8_10;
  assign t_r14_c8_12 = t_r14_c8_11 + p_15_9;
  assign out_14_8 = t_r14_c8_12 >> 4;

  assign t_r14_c9_0 = p_13_9 << 1;
  assign t_r14_c9_1 = p_14_8 << 1;
  assign t_r14_c9_2 = p_14_9 << 2;
  assign t_r14_c9_3 = p_14_10 << 1;
  assign t_r14_c9_4 = p_15_9 << 1;
  assign t_r14_c9_5 = t_r14_c9_0 + p_13_8;
  assign t_r14_c9_6 = t_r14_c9_1 + p_13_10;
  assign t_r14_c9_7 = t_r14_c9_2 + t_r14_c9_3;
  assign t_r14_c9_8 = t_r14_c9_4 + p_15_8;
  assign t_r14_c9_9 = t_r14_c9_5 + t_r14_c9_6;
  assign t_r14_c9_10 = t_r14_c9_7 + t_r14_c9_8;
  assign t_r14_c9_11 = t_r14_c9_9 + t_r14_c9_10;
  assign t_r14_c9_12 = t_r14_c9_11 + p_15_10;
  assign out_14_9 = t_r14_c9_12 >> 4;

  assign t_r14_c10_0 = p_13_10 << 1;
  assign t_r14_c10_1 = p_14_9 << 1;
  assign t_r14_c10_2 = p_14_10 << 2;
  assign t_r14_c10_3 = p_14_11 << 1;
  assign t_r14_c10_4 = p_15_10 << 1;
  assign t_r14_c10_5 = t_r14_c10_0 + p_13_9;
  assign t_r14_c10_6 = t_r14_c10_1 + p_13_11;
  assign t_r14_c10_7 = t_r14_c10_2 + t_r14_c10_3;
  assign t_r14_c10_8 = t_r14_c10_4 + p_15_9;
  assign t_r14_c10_9 = t_r14_c10_5 + t_r14_c10_6;
  assign t_r14_c10_10 = t_r14_c10_7 + t_r14_c10_8;
  assign t_r14_c10_11 = t_r14_c10_9 + t_r14_c10_10;
  assign t_r14_c10_12 = t_r14_c10_11 + p_15_11;
  assign out_14_10 = t_r14_c10_12 >> 4;

  assign t_r14_c11_0 = p_13_11 << 1;
  assign t_r14_c11_1 = p_14_10 << 1;
  assign t_r14_c11_2 = p_14_11 << 2;
  assign t_r14_c11_3 = p_14_12 << 1;
  assign t_r14_c11_4 = p_15_11 << 1;
  assign t_r14_c11_5 = t_r14_c11_0 + p_13_10;
  assign t_r14_c11_6 = t_r14_c11_1 + p_13_12;
  assign t_r14_c11_7 = t_r14_c11_2 + t_r14_c11_3;
  assign t_r14_c11_8 = t_r14_c11_4 + p_15_10;
  assign t_r14_c11_9 = t_r14_c11_5 + t_r14_c11_6;
  assign t_r14_c11_10 = t_r14_c11_7 + t_r14_c11_8;
  assign t_r14_c11_11 = t_r14_c11_9 + t_r14_c11_10;
  assign t_r14_c11_12 = t_r14_c11_11 + p_15_12;
  assign out_14_11 = t_r14_c11_12 >> 4;

  assign t_r14_c12_0 = p_13_12 << 1;
  assign t_r14_c12_1 = p_14_11 << 1;
  assign t_r14_c12_2 = p_14_12 << 2;
  assign t_r14_c12_3 = p_14_13 << 1;
  assign t_r14_c12_4 = p_15_12 << 1;
  assign t_r14_c12_5 = t_r14_c12_0 + p_13_11;
  assign t_r14_c12_6 = t_r14_c12_1 + p_13_13;
  assign t_r14_c12_7 = t_r14_c12_2 + t_r14_c12_3;
  assign t_r14_c12_8 = t_r14_c12_4 + p_15_11;
  assign t_r14_c12_9 = t_r14_c12_5 + t_r14_c12_6;
  assign t_r14_c12_10 = t_r14_c12_7 + t_r14_c12_8;
  assign t_r14_c12_11 = t_r14_c12_9 + t_r14_c12_10;
  assign t_r14_c12_12 = t_r14_c12_11 + p_15_13;
  assign out_14_12 = t_r14_c12_12 >> 4;

  assign t_r14_c13_0 = p_13_13 << 1;
  assign t_r14_c13_1 = p_14_12 << 1;
  assign t_r14_c13_2 = p_14_13 << 2;
  assign t_r14_c13_3 = p_14_14 << 1;
  assign t_r14_c13_4 = p_15_13 << 1;
  assign t_r14_c13_5 = t_r14_c13_0 + p_13_12;
  assign t_r14_c13_6 = t_r14_c13_1 + p_13_14;
  assign t_r14_c13_7 = t_r14_c13_2 + t_r14_c13_3;
  assign t_r14_c13_8 = t_r14_c13_4 + p_15_12;
  assign t_r14_c13_9 = t_r14_c13_5 + t_r14_c13_6;
  assign t_r14_c13_10 = t_r14_c13_7 + t_r14_c13_8;
  assign t_r14_c13_11 = t_r14_c13_9 + t_r14_c13_10;
  assign t_r14_c13_12 = t_r14_c13_11 + p_15_14;
  assign out_14_13 = t_r14_c13_12 >> 4;

  assign t_r14_c14_0 = p_13_14 << 1;
  assign t_r14_c14_1 = p_14_13 << 1;
  assign t_r14_c14_2 = p_14_14 << 2;
  assign t_r14_c14_3 = p_14_15 << 1;
  assign t_r14_c14_4 = p_15_14 << 1;
  assign t_r14_c14_5 = t_r14_c14_0 + p_13_13;
  assign t_r14_c14_6 = t_r14_c14_1 + p_13_15;
  assign t_r14_c14_7 = t_r14_c14_2 + t_r14_c14_3;
  assign t_r14_c14_8 = t_r14_c14_4 + p_15_13;
  assign t_r14_c14_9 = t_r14_c14_5 + t_r14_c14_6;
  assign t_r14_c14_10 = t_r14_c14_7 + t_r14_c14_8;
  assign t_r14_c14_11 = t_r14_c14_9 + t_r14_c14_10;
  assign t_r14_c14_12 = t_r14_c14_11 + p_15_15;
  assign out_14_14 = t_r14_c14_12 >> 4;

  assign t_r14_c15_0 = p_13_15 << 1;
  assign t_r14_c15_1 = p_14_14 << 1;
  assign t_r14_c15_2 = p_14_15 << 2;
  assign t_r14_c15_3 = p_14_16 << 1;
  assign t_r14_c15_4 = p_15_15 << 1;
  assign t_r14_c15_5 = t_r14_c15_0 + p_13_14;
  assign t_r14_c15_6 = t_r14_c15_1 + p_13_16;
  assign t_r14_c15_7 = t_r14_c15_2 + t_r14_c15_3;
  assign t_r14_c15_8 = t_r14_c15_4 + p_15_14;
  assign t_r14_c15_9 = t_r14_c15_5 + t_r14_c15_6;
  assign t_r14_c15_10 = t_r14_c15_7 + t_r14_c15_8;
  assign t_r14_c15_11 = t_r14_c15_9 + t_r14_c15_10;
  assign t_r14_c15_12 = t_r14_c15_11 + p_15_16;
  assign out_14_15 = t_r14_c15_12 >> 4;

  assign t_r14_c16_0 = p_13_16 << 1;
  assign t_r14_c16_1 = p_14_15 << 1;
  assign t_r14_c16_2 = p_14_16 << 2;
  assign t_r14_c16_3 = p_14_17 << 1;
  assign t_r14_c16_4 = p_15_16 << 1;
  assign t_r14_c16_5 = t_r14_c16_0 + p_13_15;
  assign t_r14_c16_6 = t_r14_c16_1 + p_13_17;
  assign t_r14_c16_7 = t_r14_c16_2 + t_r14_c16_3;
  assign t_r14_c16_8 = t_r14_c16_4 + p_15_15;
  assign t_r14_c16_9 = t_r14_c16_5 + t_r14_c16_6;
  assign t_r14_c16_10 = t_r14_c16_7 + t_r14_c16_8;
  assign t_r14_c16_11 = t_r14_c16_9 + t_r14_c16_10;
  assign t_r14_c16_12 = t_r14_c16_11 + p_15_17;
  assign out_14_16 = t_r14_c16_12 >> 4;

  assign t_r14_c17_0 = p_13_17 << 1;
  assign t_r14_c17_1 = p_14_16 << 1;
  assign t_r14_c17_2 = p_14_17 << 2;
  assign t_r14_c17_3 = p_14_18 << 1;
  assign t_r14_c17_4 = p_15_17 << 1;
  assign t_r14_c17_5 = t_r14_c17_0 + p_13_16;
  assign t_r14_c17_6 = t_r14_c17_1 + p_13_18;
  assign t_r14_c17_7 = t_r14_c17_2 + t_r14_c17_3;
  assign t_r14_c17_8 = t_r14_c17_4 + p_15_16;
  assign t_r14_c17_9 = t_r14_c17_5 + t_r14_c17_6;
  assign t_r14_c17_10 = t_r14_c17_7 + t_r14_c17_8;
  assign t_r14_c17_11 = t_r14_c17_9 + t_r14_c17_10;
  assign t_r14_c17_12 = t_r14_c17_11 + p_15_18;
  assign out_14_17 = t_r14_c17_12 >> 4;

  assign t_r14_c18_0 = p_13_18 << 1;
  assign t_r14_c18_1 = p_14_17 << 1;
  assign t_r14_c18_2 = p_14_18 << 2;
  assign t_r14_c18_3 = p_14_19 << 1;
  assign t_r14_c18_4 = p_15_18 << 1;
  assign t_r14_c18_5 = t_r14_c18_0 + p_13_17;
  assign t_r14_c18_6 = t_r14_c18_1 + p_13_19;
  assign t_r14_c18_7 = t_r14_c18_2 + t_r14_c18_3;
  assign t_r14_c18_8 = t_r14_c18_4 + p_15_17;
  assign t_r14_c18_9 = t_r14_c18_5 + t_r14_c18_6;
  assign t_r14_c18_10 = t_r14_c18_7 + t_r14_c18_8;
  assign t_r14_c18_11 = t_r14_c18_9 + t_r14_c18_10;
  assign t_r14_c18_12 = t_r14_c18_11 + p_15_19;
  assign out_14_18 = t_r14_c18_12 >> 4;

  assign t_r14_c19_0 = p_13_19 << 1;
  assign t_r14_c19_1 = p_14_18 << 1;
  assign t_r14_c19_2 = p_14_19 << 2;
  assign t_r14_c19_3 = p_14_20 << 1;
  assign t_r14_c19_4 = p_15_19 << 1;
  assign t_r14_c19_5 = t_r14_c19_0 + p_13_18;
  assign t_r14_c19_6 = t_r14_c19_1 + p_13_20;
  assign t_r14_c19_7 = t_r14_c19_2 + t_r14_c19_3;
  assign t_r14_c19_8 = t_r14_c19_4 + p_15_18;
  assign t_r14_c19_9 = t_r14_c19_5 + t_r14_c19_6;
  assign t_r14_c19_10 = t_r14_c19_7 + t_r14_c19_8;
  assign t_r14_c19_11 = t_r14_c19_9 + t_r14_c19_10;
  assign t_r14_c19_12 = t_r14_c19_11 + p_15_20;
  assign out_14_19 = t_r14_c19_12 >> 4;

  assign t_r14_c20_0 = p_13_20 << 1;
  assign t_r14_c20_1 = p_14_19 << 1;
  assign t_r14_c20_2 = p_14_20 << 2;
  assign t_r14_c20_3 = p_14_21 << 1;
  assign t_r14_c20_4 = p_15_20 << 1;
  assign t_r14_c20_5 = t_r14_c20_0 + p_13_19;
  assign t_r14_c20_6 = t_r14_c20_1 + p_13_21;
  assign t_r14_c20_7 = t_r14_c20_2 + t_r14_c20_3;
  assign t_r14_c20_8 = t_r14_c20_4 + p_15_19;
  assign t_r14_c20_9 = t_r14_c20_5 + t_r14_c20_6;
  assign t_r14_c20_10 = t_r14_c20_7 + t_r14_c20_8;
  assign t_r14_c20_11 = t_r14_c20_9 + t_r14_c20_10;
  assign t_r14_c20_12 = t_r14_c20_11 + p_15_21;
  assign out_14_20 = t_r14_c20_12 >> 4;

  assign t_r14_c21_0 = p_13_21 << 1;
  assign t_r14_c21_1 = p_14_20 << 1;
  assign t_r14_c21_2 = p_14_21 << 2;
  assign t_r14_c21_3 = p_14_22 << 1;
  assign t_r14_c21_4 = p_15_21 << 1;
  assign t_r14_c21_5 = t_r14_c21_0 + p_13_20;
  assign t_r14_c21_6 = t_r14_c21_1 + p_13_22;
  assign t_r14_c21_7 = t_r14_c21_2 + t_r14_c21_3;
  assign t_r14_c21_8 = t_r14_c21_4 + p_15_20;
  assign t_r14_c21_9 = t_r14_c21_5 + t_r14_c21_6;
  assign t_r14_c21_10 = t_r14_c21_7 + t_r14_c21_8;
  assign t_r14_c21_11 = t_r14_c21_9 + t_r14_c21_10;
  assign t_r14_c21_12 = t_r14_c21_11 + p_15_22;
  assign out_14_21 = t_r14_c21_12 >> 4;

  assign t_r14_c22_0 = p_13_22 << 1;
  assign t_r14_c22_1 = p_14_21 << 1;
  assign t_r14_c22_2 = p_14_22 << 2;
  assign t_r14_c22_3 = p_14_23 << 1;
  assign t_r14_c22_4 = p_15_22 << 1;
  assign t_r14_c22_5 = t_r14_c22_0 + p_13_21;
  assign t_r14_c22_6 = t_r14_c22_1 + p_13_23;
  assign t_r14_c22_7 = t_r14_c22_2 + t_r14_c22_3;
  assign t_r14_c22_8 = t_r14_c22_4 + p_15_21;
  assign t_r14_c22_9 = t_r14_c22_5 + t_r14_c22_6;
  assign t_r14_c22_10 = t_r14_c22_7 + t_r14_c22_8;
  assign t_r14_c22_11 = t_r14_c22_9 + t_r14_c22_10;
  assign t_r14_c22_12 = t_r14_c22_11 + p_15_23;
  assign out_14_22 = t_r14_c22_12 >> 4;

  assign t_r14_c23_0 = p_13_23 << 1;
  assign t_r14_c23_1 = p_14_22 << 1;
  assign t_r14_c23_2 = p_14_23 << 2;
  assign t_r14_c23_3 = p_14_24 << 1;
  assign t_r14_c23_4 = p_15_23 << 1;
  assign t_r14_c23_5 = t_r14_c23_0 + p_13_22;
  assign t_r14_c23_6 = t_r14_c23_1 + p_13_24;
  assign t_r14_c23_7 = t_r14_c23_2 + t_r14_c23_3;
  assign t_r14_c23_8 = t_r14_c23_4 + p_15_22;
  assign t_r14_c23_9 = t_r14_c23_5 + t_r14_c23_6;
  assign t_r14_c23_10 = t_r14_c23_7 + t_r14_c23_8;
  assign t_r14_c23_11 = t_r14_c23_9 + t_r14_c23_10;
  assign t_r14_c23_12 = t_r14_c23_11 + p_15_24;
  assign out_14_23 = t_r14_c23_12 >> 4;

  assign t_r14_c24_0 = p_13_24 << 1;
  assign t_r14_c24_1 = p_14_23 << 1;
  assign t_r14_c24_2 = p_14_24 << 2;
  assign t_r14_c24_3 = p_14_25 << 1;
  assign t_r14_c24_4 = p_15_24 << 1;
  assign t_r14_c24_5 = t_r14_c24_0 + p_13_23;
  assign t_r14_c24_6 = t_r14_c24_1 + p_13_25;
  assign t_r14_c24_7 = t_r14_c24_2 + t_r14_c24_3;
  assign t_r14_c24_8 = t_r14_c24_4 + p_15_23;
  assign t_r14_c24_9 = t_r14_c24_5 + t_r14_c24_6;
  assign t_r14_c24_10 = t_r14_c24_7 + t_r14_c24_8;
  assign t_r14_c24_11 = t_r14_c24_9 + t_r14_c24_10;
  assign t_r14_c24_12 = t_r14_c24_11 + p_15_25;
  assign out_14_24 = t_r14_c24_12 >> 4;

  assign t_r14_c25_0 = p_13_25 << 1;
  assign t_r14_c25_1 = p_14_24 << 1;
  assign t_r14_c25_2 = p_14_25 << 2;
  assign t_r14_c25_3 = p_14_26 << 1;
  assign t_r14_c25_4 = p_15_25 << 1;
  assign t_r14_c25_5 = t_r14_c25_0 + p_13_24;
  assign t_r14_c25_6 = t_r14_c25_1 + p_13_26;
  assign t_r14_c25_7 = t_r14_c25_2 + t_r14_c25_3;
  assign t_r14_c25_8 = t_r14_c25_4 + p_15_24;
  assign t_r14_c25_9 = t_r14_c25_5 + t_r14_c25_6;
  assign t_r14_c25_10 = t_r14_c25_7 + t_r14_c25_8;
  assign t_r14_c25_11 = t_r14_c25_9 + t_r14_c25_10;
  assign t_r14_c25_12 = t_r14_c25_11 + p_15_26;
  assign out_14_25 = t_r14_c25_12 >> 4;

  assign t_r14_c26_0 = p_13_26 << 1;
  assign t_r14_c26_1 = p_14_25 << 1;
  assign t_r14_c26_2 = p_14_26 << 2;
  assign t_r14_c26_3 = p_14_27 << 1;
  assign t_r14_c26_4 = p_15_26 << 1;
  assign t_r14_c26_5 = t_r14_c26_0 + p_13_25;
  assign t_r14_c26_6 = t_r14_c26_1 + p_13_27;
  assign t_r14_c26_7 = t_r14_c26_2 + t_r14_c26_3;
  assign t_r14_c26_8 = t_r14_c26_4 + p_15_25;
  assign t_r14_c26_9 = t_r14_c26_5 + t_r14_c26_6;
  assign t_r14_c26_10 = t_r14_c26_7 + t_r14_c26_8;
  assign t_r14_c26_11 = t_r14_c26_9 + t_r14_c26_10;
  assign t_r14_c26_12 = t_r14_c26_11 + p_15_27;
  assign out_14_26 = t_r14_c26_12 >> 4;

  assign t_r14_c27_0 = p_13_27 << 1;
  assign t_r14_c27_1 = p_14_26 << 1;
  assign t_r14_c27_2 = p_14_27 << 2;
  assign t_r14_c27_3 = p_14_28 << 1;
  assign t_r14_c27_4 = p_15_27 << 1;
  assign t_r14_c27_5 = t_r14_c27_0 + p_13_26;
  assign t_r14_c27_6 = t_r14_c27_1 + p_13_28;
  assign t_r14_c27_7 = t_r14_c27_2 + t_r14_c27_3;
  assign t_r14_c27_8 = t_r14_c27_4 + p_15_26;
  assign t_r14_c27_9 = t_r14_c27_5 + t_r14_c27_6;
  assign t_r14_c27_10 = t_r14_c27_7 + t_r14_c27_8;
  assign t_r14_c27_11 = t_r14_c27_9 + t_r14_c27_10;
  assign t_r14_c27_12 = t_r14_c27_11 + p_15_28;
  assign out_14_27 = t_r14_c27_12 >> 4;

  assign t_r14_c28_0 = p_13_28 << 1;
  assign t_r14_c28_1 = p_14_27 << 1;
  assign t_r14_c28_2 = p_14_28 << 2;
  assign t_r14_c28_3 = p_14_29 << 1;
  assign t_r14_c28_4 = p_15_28 << 1;
  assign t_r14_c28_5 = t_r14_c28_0 + p_13_27;
  assign t_r14_c28_6 = t_r14_c28_1 + p_13_29;
  assign t_r14_c28_7 = t_r14_c28_2 + t_r14_c28_3;
  assign t_r14_c28_8 = t_r14_c28_4 + p_15_27;
  assign t_r14_c28_9 = t_r14_c28_5 + t_r14_c28_6;
  assign t_r14_c28_10 = t_r14_c28_7 + t_r14_c28_8;
  assign t_r14_c28_11 = t_r14_c28_9 + t_r14_c28_10;
  assign t_r14_c28_12 = t_r14_c28_11 + p_15_29;
  assign out_14_28 = t_r14_c28_12 >> 4;

  assign t_r14_c29_0 = p_13_29 << 1;
  assign t_r14_c29_1 = p_14_28 << 1;
  assign t_r14_c29_2 = p_14_29 << 2;
  assign t_r14_c29_3 = p_14_30 << 1;
  assign t_r14_c29_4 = p_15_29 << 1;
  assign t_r14_c29_5 = t_r14_c29_0 + p_13_28;
  assign t_r14_c29_6 = t_r14_c29_1 + p_13_30;
  assign t_r14_c29_7 = t_r14_c29_2 + t_r14_c29_3;
  assign t_r14_c29_8 = t_r14_c29_4 + p_15_28;
  assign t_r14_c29_9 = t_r14_c29_5 + t_r14_c29_6;
  assign t_r14_c29_10 = t_r14_c29_7 + t_r14_c29_8;
  assign t_r14_c29_11 = t_r14_c29_9 + t_r14_c29_10;
  assign t_r14_c29_12 = t_r14_c29_11 + p_15_30;
  assign out_14_29 = t_r14_c29_12 >> 4;

  assign t_r14_c30_0 = p_13_30 << 1;
  assign t_r14_c30_1 = p_14_29 << 1;
  assign t_r14_c30_2 = p_14_30 << 2;
  assign t_r14_c30_3 = p_14_31 << 1;
  assign t_r14_c30_4 = p_15_30 << 1;
  assign t_r14_c30_5 = t_r14_c30_0 + p_13_29;
  assign t_r14_c30_6 = t_r14_c30_1 + p_13_31;
  assign t_r14_c30_7 = t_r14_c30_2 + t_r14_c30_3;
  assign t_r14_c30_8 = t_r14_c30_4 + p_15_29;
  assign t_r14_c30_9 = t_r14_c30_5 + t_r14_c30_6;
  assign t_r14_c30_10 = t_r14_c30_7 + t_r14_c30_8;
  assign t_r14_c30_11 = t_r14_c30_9 + t_r14_c30_10;
  assign t_r14_c30_12 = t_r14_c30_11 + p_15_31;
  assign out_14_30 = t_r14_c30_12 >> 4;

  assign t_r14_c31_0 = p_13_31 << 1;
  assign t_r14_c31_1 = p_14_30 << 1;
  assign t_r14_c31_2 = p_14_31 << 2;
  assign t_r14_c31_3 = p_14_32 << 1;
  assign t_r14_c31_4 = p_15_31 << 1;
  assign t_r14_c31_5 = t_r14_c31_0 + p_13_30;
  assign t_r14_c31_6 = t_r14_c31_1 + p_13_32;
  assign t_r14_c31_7 = t_r14_c31_2 + t_r14_c31_3;
  assign t_r14_c31_8 = t_r14_c31_4 + p_15_30;
  assign t_r14_c31_9 = t_r14_c31_5 + t_r14_c31_6;
  assign t_r14_c31_10 = t_r14_c31_7 + t_r14_c31_8;
  assign t_r14_c31_11 = t_r14_c31_9 + t_r14_c31_10;
  assign t_r14_c31_12 = t_r14_c31_11 + p_15_32;
  assign out_14_31 = t_r14_c31_12 >> 4;

  assign t_r14_c32_0 = p_13_32 << 1;
  assign t_r14_c32_1 = p_14_31 << 1;
  assign t_r14_c32_2 = p_14_32 << 2;
  assign t_r14_c32_3 = p_14_33 << 1;
  assign t_r14_c32_4 = p_15_32 << 1;
  assign t_r14_c32_5 = t_r14_c32_0 + p_13_31;
  assign t_r14_c32_6 = t_r14_c32_1 + p_13_33;
  assign t_r14_c32_7 = t_r14_c32_2 + t_r14_c32_3;
  assign t_r14_c32_8 = t_r14_c32_4 + p_15_31;
  assign t_r14_c32_9 = t_r14_c32_5 + t_r14_c32_6;
  assign t_r14_c32_10 = t_r14_c32_7 + t_r14_c32_8;
  assign t_r14_c32_11 = t_r14_c32_9 + t_r14_c32_10;
  assign t_r14_c32_12 = t_r14_c32_11 + p_15_33;
  assign out_14_32 = t_r14_c32_12 >> 4;

  assign t_r14_c33_0 = p_13_33 << 1;
  assign t_r14_c33_1 = p_14_32 << 1;
  assign t_r14_c33_2 = p_14_33 << 2;
  assign t_r14_c33_3 = p_14_34 << 1;
  assign t_r14_c33_4 = p_15_33 << 1;
  assign t_r14_c33_5 = t_r14_c33_0 + p_13_32;
  assign t_r14_c33_6 = t_r14_c33_1 + p_13_34;
  assign t_r14_c33_7 = t_r14_c33_2 + t_r14_c33_3;
  assign t_r14_c33_8 = t_r14_c33_4 + p_15_32;
  assign t_r14_c33_9 = t_r14_c33_5 + t_r14_c33_6;
  assign t_r14_c33_10 = t_r14_c33_7 + t_r14_c33_8;
  assign t_r14_c33_11 = t_r14_c33_9 + t_r14_c33_10;
  assign t_r14_c33_12 = t_r14_c33_11 + p_15_34;
  assign out_14_33 = t_r14_c33_12 >> 4;

  assign t_r14_c34_0 = p_13_34 << 1;
  assign t_r14_c34_1 = p_14_33 << 1;
  assign t_r14_c34_2 = p_14_34 << 2;
  assign t_r14_c34_3 = p_14_35 << 1;
  assign t_r14_c34_4 = p_15_34 << 1;
  assign t_r14_c34_5 = t_r14_c34_0 + p_13_33;
  assign t_r14_c34_6 = t_r14_c34_1 + p_13_35;
  assign t_r14_c34_7 = t_r14_c34_2 + t_r14_c34_3;
  assign t_r14_c34_8 = t_r14_c34_4 + p_15_33;
  assign t_r14_c34_9 = t_r14_c34_5 + t_r14_c34_6;
  assign t_r14_c34_10 = t_r14_c34_7 + t_r14_c34_8;
  assign t_r14_c34_11 = t_r14_c34_9 + t_r14_c34_10;
  assign t_r14_c34_12 = t_r14_c34_11 + p_15_35;
  assign out_14_34 = t_r14_c34_12 >> 4;

  assign t_r14_c35_0 = p_13_35 << 1;
  assign t_r14_c35_1 = p_14_34 << 1;
  assign t_r14_c35_2 = p_14_35 << 2;
  assign t_r14_c35_3 = p_14_36 << 1;
  assign t_r14_c35_4 = p_15_35 << 1;
  assign t_r14_c35_5 = t_r14_c35_0 + p_13_34;
  assign t_r14_c35_6 = t_r14_c35_1 + p_13_36;
  assign t_r14_c35_7 = t_r14_c35_2 + t_r14_c35_3;
  assign t_r14_c35_8 = t_r14_c35_4 + p_15_34;
  assign t_r14_c35_9 = t_r14_c35_5 + t_r14_c35_6;
  assign t_r14_c35_10 = t_r14_c35_7 + t_r14_c35_8;
  assign t_r14_c35_11 = t_r14_c35_9 + t_r14_c35_10;
  assign t_r14_c35_12 = t_r14_c35_11 + p_15_36;
  assign out_14_35 = t_r14_c35_12 >> 4;

  assign t_r14_c36_0 = p_13_36 << 1;
  assign t_r14_c36_1 = p_14_35 << 1;
  assign t_r14_c36_2 = p_14_36 << 2;
  assign t_r14_c36_3 = p_14_37 << 1;
  assign t_r14_c36_4 = p_15_36 << 1;
  assign t_r14_c36_5 = t_r14_c36_0 + p_13_35;
  assign t_r14_c36_6 = t_r14_c36_1 + p_13_37;
  assign t_r14_c36_7 = t_r14_c36_2 + t_r14_c36_3;
  assign t_r14_c36_8 = t_r14_c36_4 + p_15_35;
  assign t_r14_c36_9 = t_r14_c36_5 + t_r14_c36_6;
  assign t_r14_c36_10 = t_r14_c36_7 + t_r14_c36_8;
  assign t_r14_c36_11 = t_r14_c36_9 + t_r14_c36_10;
  assign t_r14_c36_12 = t_r14_c36_11 + p_15_37;
  assign out_14_36 = t_r14_c36_12 >> 4;

  assign t_r14_c37_0 = p_13_37 << 1;
  assign t_r14_c37_1 = p_14_36 << 1;
  assign t_r14_c37_2 = p_14_37 << 2;
  assign t_r14_c37_3 = p_14_38 << 1;
  assign t_r14_c37_4 = p_15_37 << 1;
  assign t_r14_c37_5 = t_r14_c37_0 + p_13_36;
  assign t_r14_c37_6 = t_r14_c37_1 + p_13_38;
  assign t_r14_c37_7 = t_r14_c37_2 + t_r14_c37_3;
  assign t_r14_c37_8 = t_r14_c37_4 + p_15_36;
  assign t_r14_c37_9 = t_r14_c37_5 + t_r14_c37_6;
  assign t_r14_c37_10 = t_r14_c37_7 + t_r14_c37_8;
  assign t_r14_c37_11 = t_r14_c37_9 + t_r14_c37_10;
  assign t_r14_c37_12 = t_r14_c37_11 + p_15_38;
  assign out_14_37 = t_r14_c37_12 >> 4;

  assign t_r14_c38_0 = p_13_38 << 1;
  assign t_r14_c38_1 = p_14_37 << 1;
  assign t_r14_c38_2 = p_14_38 << 2;
  assign t_r14_c38_3 = p_14_39 << 1;
  assign t_r14_c38_4 = p_15_38 << 1;
  assign t_r14_c38_5 = t_r14_c38_0 + p_13_37;
  assign t_r14_c38_6 = t_r14_c38_1 + p_13_39;
  assign t_r14_c38_7 = t_r14_c38_2 + t_r14_c38_3;
  assign t_r14_c38_8 = t_r14_c38_4 + p_15_37;
  assign t_r14_c38_9 = t_r14_c38_5 + t_r14_c38_6;
  assign t_r14_c38_10 = t_r14_c38_7 + t_r14_c38_8;
  assign t_r14_c38_11 = t_r14_c38_9 + t_r14_c38_10;
  assign t_r14_c38_12 = t_r14_c38_11 + p_15_39;
  assign out_14_38 = t_r14_c38_12 >> 4;

  assign t_r14_c39_0 = p_13_39 << 1;
  assign t_r14_c39_1 = p_14_38 << 1;
  assign t_r14_c39_2 = p_14_39 << 2;
  assign t_r14_c39_3 = p_14_40 << 1;
  assign t_r14_c39_4 = p_15_39 << 1;
  assign t_r14_c39_5 = t_r14_c39_0 + p_13_38;
  assign t_r14_c39_6 = t_r14_c39_1 + p_13_40;
  assign t_r14_c39_7 = t_r14_c39_2 + t_r14_c39_3;
  assign t_r14_c39_8 = t_r14_c39_4 + p_15_38;
  assign t_r14_c39_9 = t_r14_c39_5 + t_r14_c39_6;
  assign t_r14_c39_10 = t_r14_c39_7 + t_r14_c39_8;
  assign t_r14_c39_11 = t_r14_c39_9 + t_r14_c39_10;
  assign t_r14_c39_12 = t_r14_c39_11 + p_15_40;
  assign out_14_39 = t_r14_c39_12 >> 4;

  assign t_r14_c40_0 = p_13_40 << 1;
  assign t_r14_c40_1 = p_14_39 << 1;
  assign t_r14_c40_2 = p_14_40 << 2;
  assign t_r14_c40_3 = p_14_41 << 1;
  assign t_r14_c40_4 = p_15_40 << 1;
  assign t_r14_c40_5 = t_r14_c40_0 + p_13_39;
  assign t_r14_c40_6 = t_r14_c40_1 + p_13_41;
  assign t_r14_c40_7 = t_r14_c40_2 + t_r14_c40_3;
  assign t_r14_c40_8 = t_r14_c40_4 + p_15_39;
  assign t_r14_c40_9 = t_r14_c40_5 + t_r14_c40_6;
  assign t_r14_c40_10 = t_r14_c40_7 + t_r14_c40_8;
  assign t_r14_c40_11 = t_r14_c40_9 + t_r14_c40_10;
  assign t_r14_c40_12 = t_r14_c40_11 + p_15_41;
  assign out_14_40 = t_r14_c40_12 >> 4;

  assign t_r14_c41_0 = p_13_41 << 1;
  assign t_r14_c41_1 = p_14_40 << 1;
  assign t_r14_c41_2 = p_14_41 << 2;
  assign t_r14_c41_3 = p_14_42 << 1;
  assign t_r14_c41_4 = p_15_41 << 1;
  assign t_r14_c41_5 = t_r14_c41_0 + p_13_40;
  assign t_r14_c41_6 = t_r14_c41_1 + p_13_42;
  assign t_r14_c41_7 = t_r14_c41_2 + t_r14_c41_3;
  assign t_r14_c41_8 = t_r14_c41_4 + p_15_40;
  assign t_r14_c41_9 = t_r14_c41_5 + t_r14_c41_6;
  assign t_r14_c41_10 = t_r14_c41_7 + t_r14_c41_8;
  assign t_r14_c41_11 = t_r14_c41_9 + t_r14_c41_10;
  assign t_r14_c41_12 = t_r14_c41_11 + p_15_42;
  assign out_14_41 = t_r14_c41_12 >> 4;

  assign t_r14_c42_0 = p_13_42 << 1;
  assign t_r14_c42_1 = p_14_41 << 1;
  assign t_r14_c42_2 = p_14_42 << 2;
  assign t_r14_c42_3 = p_14_43 << 1;
  assign t_r14_c42_4 = p_15_42 << 1;
  assign t_r14_c42_5 = t_r14_c42_0 + p_13_41;
  assign t_r14_c42_6 = t_r14_c42_1 + p_13_43;
  assign t_r14_c42_7 = t_r14_c42_2 + t_r14_c42_3;
  assign t_r14_c42_8 = t_r14_c42_4 + p_15_41;
  assign t_r14_c42_9 = t_r14_c42_5 + t_r14_c42_6;
  assign t_r14_c42_10 = t_r14_c42_7 + t_r14_c42_8;
  assign t_r14_c42_11 = t_r14_c42_9 + t_r14_c42_10;
  assign t_r14_c42_12 = t_r14_c42_11 + p_15_43;
  assign out_14_42 = t_r14_c42_12 >> 4;

  assign t_r14_c43_0 = p_13_43 << 1;
  assign t_r14_c43_1 = p_14_42 << 1;
  assign t_r14_c43_2 = p_14_43 << 2;
  assign t_r14_c43_3 = p_14_44 << 1;
  assign t_r14_c43_4 = p_15_43 << 1;
  assign t_r14_c43_5 = t_r14_c43_0 + p_13_42;
  assign t_r14_c43_6 = t_r14_c43_1 + p_13_44;
  assign t_r14_c43_7 = t_r14_c43_2 + t_r14_c43_3;
  assign t_r14_c43_8 = t_r14_c43_4 + p_15_42;
  assign t_r14_c43_9 = t_r14_c43_5 + t_r14_c43_6;
  assign t_r14_c43_10 = t_r14_c43_7 + t_r14_c43_8;
  assign t_r14_c43_11 = t_r14_c43_9 + t_r14_c43_10;
  assign t_r14_c43_12 = t_r14_c43_11 + p_15_44;
  assign out_14_43 = t_r14_c43_12 >> 4;

  assign t_r14_c44_0 = p_13_44 << 1;
  assign t_r14_c44_1 = p_14_43 << 1;
  assign t_r14_c44_2 = p_14_44 << 2;
  assign t_r14_c44_3 = p_14_45 << 1;
  assign t_r14_c44_4 = p_15_44 << 1;
  assign t_r14_c44_5 = t_r14_c44_0 + p_13_43;
  assign t_r14_c44_6 = t_r14_c44_1 + p_13_45;
  assign t_r14_c44_7 = t_r14_c44_2 + t_r14_c44_3;
  assign t_r14_c44_8 = t_r14_c44_4 + p_15_43;
  assign t_r14_c44_9 = t_r14_c44_5 + t_r14_c44_6;
  assign t_r14_c44_10 = t_r14_c44_7 + t_r14_c44_8;
  assign t_r14_c44_11 = t_r14_c44_9 + t_r14_c44_10;
  assign t_r14_c44_12 = t_r14_c44_11 + p_15_45;
  assign out_14_44 = t_r14_c44_12 >> 4;

  assign t_r14_c45_0 = p_13_45 << 1;
  assign t_r14_c45_1 = p_14_44 << 1;
  assign t_r14_c45_2 = p_14_45 << 2;
  assign t_r14_c45_3 = p_14_46 << 1;
  assign t_r14_c45_4 = p_15_45 << 1;
  assign t_r14_c45_5 = t_r14_c45_0 + p_13_44;
  assign t_r14_c45_6 = t_r14_c45_1 + p_13_46;
  assign t_r14_c45_7 = t_r14_c45_2 + t_r14_c45_3;
  assign t_r14_c45_8 = t_r14_c45_4 + p_15_44;
  assign t_r14_c45_9 = t_r14_c45_5 + t_r14_c45_6;
  assign t_r14_c45_10 = t_r14_c45_7 + t_r14_c45_8;
  assign t_r14_c45_11 = t_r14_c45_9 + t_r14_c45_10;
  assign t_r14_c45_12 = t_r14_c45_11 + p_15_46;
  assign out_14_45 = t_r14_c45_12 >> 4;

  assign t_r14_c46_0 = p_13_46 << 1;
  assign t_r14_c46_1 = p_14_45 << 1;
  assign t_r14_c46_2 = p_14_46 << 2;
  assign t_r14_c46_3 = p_14_47 << 1;
  assign t_r14_c46_4 = p_15_46 << 1;
  assign t_r14_c46_5 = t_r14_c46_0 + p_13_45;
  assign t_r14_c46_6 = t_r14_c46_1 + p_13_47;
  assign t_r14_c46_7 = t_r14_c46_2 + t_r14_c46_3;
  assign t_r14_c46_8 = t_r14_c46_4 + p_15_45;
  assign t_r14_c46_9 = t_r14_c46_5 + t_r14_c46_6;
  assign t_r14_c46_10 = t_r14_c46_7 + t_r14_c46_8;
  assign t_r14_c46_11 = t_r14_c46_9 + t_r14_c46_10;
  assign t_r14_c46_12 = t_r14_c46_11 + p_15_47;
  assign out_14_46 = t_r14_c46_12 >> 4;

  assign t_r14_c47_0 = p_13_47 << 1;
  assign t_r14_c47_1 = p_14_46 << 1;
  assign t_r14_c47_2 = p_14_47 << 2;
  assign t_r14_c47_3 = p_14_48 << 1;
  assign t_r14_c47_4 = p_15_47 << 1;
  assign t_r14_c47_5 = t_r14_c47_0 + p_13_46;
  assign t_r14_c47_6 = t_r14_c47_1 + p_13_48;
  assign t_r14_c47_7 = t_r14_c47_2 + t_r14_c47_3;
  assign t_r14_c47_8 = t_r14_c47_4 + p_15_46;
  assign t_r14_c47_9 = t_r14_c47_5 + t_r14_c47_6;
  assign t_r14_c47_10 = t_r14_c47_7 + t_r14_c47_8;
  assign t_r14_c47_11 = t_r14_c47_9 + t_r14_c47_10;
  assign t_r14_c47_12 = t_r14_c47_11 + p_15_48;
  assign out_14_47 = t_r14_c47_12 >> 4;

  assign t_r14_c48_0 = p_13_48 << 1;
  assign t_r14_c48_1 = p_14_47 << 1;
  assign t_r14_c48_2 = p_14_48 << 2;
  assign t_r14_c48_3 = p_14_49 << 1;
  assign t_r14_c48_4 = p_15_48 << 1;
  assign t_r14_c48_5 = t_r14_c48_0 + p_13_47;
  assign t_r14_c48_6 = t_r14_c48_1 + p_13_49;
  assign t_r14_c48_7 = t_r14_c48_2 + t_r14_c48_3;
  assign t_r14_c48_8 = t_r14_c48_4 + p_15_47;
  assign t_r14_c48_9 = t_r14_c48_5 + t_r14_c48_6;
  assign t_r14_c48_10 = t_r14_c48_7 + t_r14_c48_8;
  assign t_r14_c48_11 = t_r14_c48_9 + t_r14_c48_10;
  assign t_r14_c48_12 = t_r14_c48_11 + p_15_49;
  assign out_14_48 = t_r14_c48_12 >> 4;

  assign t_r14_c49_0 = p_13_49 << 1;
  assign t_r14_c49_1 = p_14_48 << 1;
  assign t_r14_c49_2 = p_14_49 << 2;
  assign t_r14_c49_3 = p_14_50 << 1;
  assign t_r14_c49_4 = p_15_49 << 1;
  assign t_r14_c49_5 = t_r14_c49_0 + p_13_48;
  assign t_r14_c49_6 = t_r14_c49_1 + p_13_50;
  assign t_r14_c49_7 = t_r14_c49_2 + t_r14_c49_3;
  assign t_r14_c49_8 = t_r14_c49_4 + p_15_48;
  assign t_r14_c49_9 = t_r14_c49_5 + t_r14_c49_6;
  assign t_r14_c49_10 = t_r14_c49_7 + t_r14_c49_8;
  assign t_r14_c49_11 = t_r14_c49_9 + t_r14_c49_10;
  assign t_r14_c49_12 = t_r14_c49_11 + p_15_50;
  assign out_14_49 = t_r14_c49_12 >> 4;

  assign t_r14_c50_0 = p_13_50 << 1;
  assign t_r14_c50_1 = p_14_49 << 1;
  assign t_r14_c50_2 = p_14_50 << 2;
  assign t_r14_c50_3 = p_14_51 << 1;
  assign t_r14_c50_4 = p_15_50 << 1;
  assign t_r14_c50_5 = t_r14_c50_0 + p_13_49;
  assign t_r14_c50_6 = t_r14_c50_1 + p_13_51;
  assign t_r14_c50_7 = t_r14_c50_2 + t_r14_c50_3;
  assign t_r14_c50_8 = t_r14_c50_4 + p_15_49;
  assign t_r14_c50_9 = t_r14_c50_5 + t_r14_c50_6;
  assign t_r14_c50_10 = t_r14_c50_7 + t_r14_c50_8;
  assign t_r14_c50_11 = t_r14_c50_9 + t_r14_c50_10;
  assign t_r14_c50_12 = t_r14_c50_11 + p_15_51;
  assign out_14_50 = t_r14_c50_12 >> 4;

  assign t_r14_c51_0 = p_13_51 << 1;
  assign t_r14_c51_1 = p_14_50 << 1;
  assign t_r14_c51_2 = p_14_51 << 2;
  assign t_r14_c51_3 = p_14_52 << 1;
  assign t_r14_c51_4 = p_15_51 << 1;
  assign t_r14_c51_5 = t_r14_c51_0 + p_13_50;
  assign t_r14_c51_6 = t_r14_c51_1 + p_13_52;
  assign t_r14_c51_7 = t_r14_c51_2 + t_r14_c51_3;
  assign t_r14_c51_8 = t_r14_c51_4 + p_15_50;
  assign t_r14_c51_9 = t_r14_c51_5 + t_r14_c51_6;
  assign t_r14_c51_10 = t_r14_c51_7 + t_r14_c51_8;
  assign t_r14_c51_11 = t_r14_c51_9 + t_r14_c51_10;
  assign t_r14_c51_12 = t_r14_c51_11 + p_15_52;
  assign out_14_51 = t_r14_c51_12 >> 4;

  assign t_r14_c52_0 = p_13_52 << 1;
  assign t_r14_c52_1 = p_14_51 << 1;
  assign t_r14_c52_2 = p_14_52 << 2;
  assign t_r14_c52_3 = p_14_53 << 1;
  assign t_r14_c52_4 = p_15_52 << 1;
  assign t_r14_c52_5 = t_r14_c52_0 + p_13_51;
  assign t_r14_c52_6 = t_r14_c52_1 + p_13_53;
  assign t_r14_c52_7 = t_r14_c52_2 + t_r14_c52_3;
  assign t_r14_c52_8 = t_r14_c52_4 + p_15_51;
  assign t_r14_c52_9 = t_r14_c52_5 + t_r14_c52_6;
  assign t_r14_c52_10 = t_r14_c52_7 + t_r14_c52_8;
  assign t_r14_c52_11 = t_r14_c52_9 + t_r14_c52_10;
  assign t_r14_c52_12 = t_r14_c52_11 + p_15_53;
  assign out_14_52 = t_r14_c52_12 >> 4;

  assign t_r14_c53_0 = p_13_53 << 1;
  assign t_r14_c53_1 = p_14_52 << 1;
  assign t_r14_c53_2 = p_14_53 << 2;
  assign t_r14_c53_3 = p_14_54 << 1;
  assign t_r14_c53_4 = p_15_53 << 1;
  assign t_r14_c53_5 = t_r14_c53_0 + p_13_52;
  assign t_r14_c53_6 = t_r14_c53_1 + p_13_54;
  assign t_r14_c53_7 = t_r14_c53_2 + t_r14_c53_3;
  assign t_r14_c53_8 = t_r14_c53_4 + p_15_52;
  assign t_r14_c53_9 = t_r14_c53_5 + t_r14_c53_6;
  assign t_r14_c53_10 = t_r14_c53_7 + t_r14_c53_8;
  assign t_r14_c53_11 = t_r14_c53_9 + t_r14_c53_10;
  assign t_r14_c53_12 = t_r14_c53_11 + p_15_54;
  assign out_14_53 = t_r14_c53_12 >> 4;

  assign t_r14_c54_0 = p_13_54 << 1;
  assign t_r14_c54_1 = p_14_53 << 1;
  assign t_r14_c54_2 = p_14_54 << 2;
  assign t_r14_c54_3 = p_14_55 << 1;
  assign t_r14_c54_4 = p_15_54 << 1;
  assign t_r14_c54_5 = t_r14_c54_0 + p_13_53;
  assign t_r14_c54_6 = t_r14_c54_1 + p_13_55;
  assign t_r14_c54_7 = t_r14_c54_2 + t_r14_c54_3;
  assign t_r14_c54_8 = t_r14_c54_4 + p_15_53;
  assign t_r14_c54_9 = t_r14_c54_5 + t_r14_c54_6;
  assign t_r14_c54_10 = t_r14_c54_7 + t_r14_c54_8;
  assign t_r14_c54_11 = t_r14_c54_9 + t_r14_c54_10;
  assign t_r14_c54_12 = t_r14_c54_11 + p_15_55;
  assign out_14_54 = t_r14_c54_12 >> 4;

  assign t_r14_c55_0 = p_13_55 << 1;
  assign t_r14_c55_1 = p_14_54 << 1;
  assign t_r14_c55_2 = p_14_55 << 2;
  assign t_r14_c55_3 = p_14_56 << 1;
  assign t_r14_c55_4 = p_15_55 << 1;
  assign t_r14_c55_5 = t_r14_c55_0 + p_13_54;
  assign t_r14_c55_6 = t_r14_c55_1 + p_13_56;
  assign t_r14_c55_7 = t_r14_c55_2 + t_r14_c55_3;
  assign t_r14_c55_8 = t_r14_c55_4 + p_15_54;
  assign t_r14_c55_9 = t_r14_c55_5 + t_r14_c55_6;
  assign t_r14_c55_10 = t_r14_c55_7 + t_r14_c55_8;
  assign t_r14_c55_11 = t_r14_c55_9 + t_r14_c55_10;
  assign t_r14_c55_12 = t_r14_c55_11 + p_15_56;
  assign out_14_55 = t_r14_c55_12 >> 4;

  assign t_r14_c56_0 = p_13_56 << 1;
  assign t_r14_c56_1 = p_14_55 << 1;
  assign t_r14_c56_2 = p_14_56 << 2;
  assign t_r14_c56_3 = p_14_57 << 1;
  assign t_r14_c56_4 = p_15_56 << 1;
  assign t_r14_c56_5 = t_r14_c56_0 + p_13_55;
  assign t_r14_c56_6 = t_r14_c56_1 + p_13_57;
  assign t_r14_c56_7 = t_r14_c56_2 + t_r14_c56_3;
  assign t_r14_c56_8 = t_r14_c56_4 + p_15_55;
  assign t_r14_c56_9 = t_r14_c56_5 + t_r14_c56_6;
  assign t_r14_c56_10 = t_r14_c56_7 + t_r14_c56_8;
  assign t_r14_c56_11 = t_r14_c56_9 + t_r14_c56_10;
  assign t_r14_c56_12 = t_r14_c56_11 + p_15_57;
  assign out_14_56 = t_r14_c56_12 >> 4;

  assign t_r14_c57_0 = p_13_57 << 1;
  assign t_r14_c57_1 = p_14_56 << 1;
  assign t_r14_c57_2 = p_14_57 << 2;
  assign t_r14_c57_3 = p_14_58 << 1;
  assign t_r14_c57_4 = p_15_57 << 1;
  assign t_r14_c57_5 = t_r14_c57_0 + p_13_56;
  assign t_r14_c57_6 = t_r14_c57_1 + p_13_58;
  assign t_r14_c57_7 = t_r14_c57_2 + t_r14_c57_3;
  assign t_r14_c57_8 = t_r14_c57_4 + p_15_56;
  assign t_r14_c57_9 = t_r14_c57_5 + t_r14_c57_6;
  assign t_r14_c57_10 = t_r14_c57_7 + t_r14_c57_8;
  assign t_r14_c57_11 = t_r14_c57_9 + t_r14_c57_10;
  assign t_r14_c57_12 = t_r14_c57_11 + p_15_58;
  assign out_14_57 = t_r14_c57_12 >> 4;

  assign t_r14_c58_0 = p_13_58 << 1;
  assign t_r14_c58_1 = p_14_57 << 1;
  assign t_r14_c58_2 = p_14_58 << 2;
  assign t_r14_c58_3 = p_14_59 << 1;
  assign t_r14_c58_4 = p_15_58 << 1;
  assign t_r14_c58_5 = t_r14_c58_0 + p_13_57;
  assign t_r14_c58_6 = t_r14_c58_1 + p_13_59;
  assign t_r14_c58_7 = t_r14_c58_2 + t_r14_c58_3;
  assign t_r14_c58_8 = t_r14_c58_4 + p_15_57;
  assign t_r14_c58_9 = t_r14_c58_5 + t_r14_c58_6;
  assign t_r14_c58_10 = t_r14_c58_7 + t_r14_c58_8;
  assign t_r14_c58_11 = t_r14_c58_9 + t_r14_c58_10;
  assign t_r14_c58_12 = t_r14_c58_11 + p_15_59;
  assign out_14_58 = t_r14_c58_12 >> 4;

  assign t_r14_c59_0 = p_13_59 << 1;
  assign t_r14_c59_1 = p_14_58 << 1;
  assign t_r14_c59_2 = p_14_59 << 2;
  assign t_r14_c59_3 = p_14_60 << 1;
  assign t_r14_c59_4 = p_15_59 << 1;
  assign t_r14_c59_5 = t_r14_c59_0 + p_13_58;
  assign t_r14_c59_6 = t_r14_c59_1 + p_13_60;
  assign t_r14_c59_7 = t_r14_c59_2 + t_r14_c59_3;
  assign t_r14_c59_8 = t_r14_c59_4 + p_15_58;
  assign t_r14_c59_9 = t_r14_c59_5 + t_r14_c59_6;
  assign t_r14_c59_10 = t_r14_c59_7 + t_r14_c59_8;
  assign t_r14_c59_11 = t_r14_c59_9 + t_r14_c59_10;
  assign t_r14_c59_12 = t_r14_c59_11 + p_15_60;
  assign out_14_59 = t_r14_c59_12 >> 4;

  assign t_r14_c60_0 = p_13_60 << 1;
  assign t_r14_c60_1 = p_14_59 << 1;
  assign t_r14_c60_2 = p_14_60 << 2;
  assign t_r14_c60_3 = p_14_61 << 1;
  assign t_r14_c60_4 = p_15_60 << 1;
  assign t_r14_c60_5 = t_r14_c60_0 + p_13_59;
  assign t_r14_c60_6 = t_r14_c60_1 + p_13_61;
  assign t_r14_c60_7 = t_r14_c60_2 + t_r14_c60_3;
  assign t_r14_c60_8 = t_r14_c60_4 + p_15_59;
  assign t_r14_c60_9 = t_r14_c60_5 + t_r14_c60_6;
  assign t_r14_c60_10 = t_r14_c60_7 + t_r14_c60_8;
  assign t_r14_c60_11 = t_r14_c60_9 + t_r14_c60_10;
  assign t_r14_c60_12 = t_r14_c60_11 + p_15_61;
  assign out_14_60 = t_r14_c60_12 >> 4;

  assign t_r14_c61_0 = p_13_61 << 1;
  assign t_r14_c61_1 = p_14_60 << 1;
  assign t_r14_c61_2 = p_14_61 << 2;
  assign t_r14_c61_3 = p_14_62 << 1;
  assign t_r14_c61_4 = p_15_61 << 1;
  assign t_r14_c61_5 = t_r14_c61_0 + p_13_60;
  assign t_r14_c61_6 = t_r14_c61_1 + p_13_62;
  assign t_r14_c61_7 = t_r14_c61_2 + t_r14_c61_3;
  assign t_r14_c61_8 = t_r14_c61_4 + p_15_60;
  assign t_r14_c61_9 = t_r14_c61_5 + t_r14_c61_6;
  assign t_r14_c61_10 = t_r14_c61_7 + t_r14_c61_8;
  assign t_r14_c61_11 = t_r14_c61_9 + t_r14_c61_10;
  assign t_r14_c61_12 = t_r14_c61_11 + p_15_62;
  assign out_14_61 = t_r14_c61_12 >> 4;

  assign t_r14_c62_0 = p_13_62 << 1;
  assign t_r14_c62_1 = p_14_61 << 1;
  assign t_r14_c62_2 = p_14_62 << 2;
  assign t_r14_c62_3 = p_14_63 << 1;
  assign t_r14_c62_4 = p_15_62 << 1;
  assign t_r14_c62_5 = t_r14_c62_0 + p_13_61;
  assign t_r14_c62_6 = t_r14_c62_1 + p_13_63;
  assign t_r14_c62_7 = t_r14_c62_2 + t_r14_c62_3;
  assign t_r14_c62_8 = t_r14_c62_4 + p_15_61;
  assign t_r14_c62_9 = t_r14_c62_5 + t_r14_c62_6;
  assign t_r14_c62_10 = t_r14_c62_7 + t_r14_c62_8;
  assign t_r14_c62_11 = t_r14_c62_9 + t_r14_c62_10;
  assign t_r14_c62_12 = t_r14_c62_11 + p_15_63;
  assign out_14_62 = t_r14_c62_12 >> 4;

  assign t_r14_c63_0 = p_13_63 << 1;
  assign t_r14_c63_1 = p_14_62 << 1;
  assign t_r14_c63_2 = p_14_63 << 2;
  assign t_r14_c63_3 = p_14_64 << 1;
  assign t_r14_c63_4 = p_15_63 << 1;
  assign t_r14_c63_5 = t_r14_c63_0 + p_13_62;
  assign t_r14_c63_6 = t_r14_c63_1 + p_13_64;
  assign t_r14_c63_7 = t_r14_c63_2 + t_r14_c63_3;
  assign t_r14_c63_8 = t_r14_c63_4 + p_15_62;
  assign t_r14_c63_9 = t_r14_c63_5 + t_r14_c63_6;
  assign t_r14_c63_10 = t_r14_c63_7 + t_r14_c63_8;
  assign t_r14_c63_11 = t_r14_c63_9 + t_r14_c63_10;
  assign t_r14_c63_12 = t_r14_c63_11 + p_15_64;
  assign out_14_63 = t_r14_c63_12 >> 4;

  assign t_r14_c64_0 = p_13_64 << 1;
  assign t_r14_c64_1 = p_14_63 << 1;
  assign t_r14_c64_2 = p_14_64 << 2;
  assign t_r14_c64_3 = p_14_65 << 1;
  assign t_r14_c64_4 = p_15_64 << 1;
  assign t_r14_c64_5 = t_r14_c64_0 + p_13_63;
  assign t_r14_c64_6 = t_r14_c64_1 + p_13_65;
  assign t_r14_c64_7 = t_r14_c64_2 + t_r14_c64_3;
  assign t_r14_c64_8 = t_r14_c64_4 + p_15_63;
  assign t_r14_c64_9 = t_r14_c64_5 + t_r14_c64_6;
  assign t_r14_c64_10 = t_r14_c64_7 + t_r14_c64_8;
  assign t_r14_c64_11 = t_r14_c64_9 + t_r14_c64_10;
  assign t_r14_c64_12 = t_r14_c64_11 + p_15_65;
  assign out_14_64 = t_r14_c64_12 >> 4;

  assign t_r15_c1_0 = p_14_1 << 1;
  assign t_r15_c1_1 = p_15_0 << 1;
  assign t_r15_c1_2 = p_15_1 << 2;
  assign t_r15_c1_3 = p_15_2 << 1;
  assign t_r15_c1_4 = p_16_1 << 1;
  assign t_r15_c1_5 = t_r15_c1_0 + p_14_0;
  assign t_r15_c1_6 = t_r15_c1_1 + p_14_2;
  assign t_r15_c1_7 = t_r15_c1_2 + t_r15_c1_3;
  assign t_r15_c1_8 = t_r15_c1_4 + p_16_0;
  assign t_r15_c1_9 = t_r15_c1_5 + t_r15_c1_6;
  assign t_r15_c1_10 = t_r15_c1_7 + t_r15_c1_8;
  assign t_r15_c1_11 = t_r15_c1_9 + t_r15_c1_10;
  assign t_r15_c1_12 = t_r15_c1_11 + p_16_2;
  assign out_15_1 = t_r15_c1_12 >> 4;

  assign t_r15_c2_0 = p_14_2 << 1;
  assign t_r15_c2_1 = p_15_1 << 1;
  assign t_r15_c2_2 = p_15_2 << 2;
  assign t_r15_c2_3 = p_15_3 << 1;
  assign t_r15_c2_4 = p_16_2 << 1;
  assign t_r15_c2_5 = t_r15_c2_0 + p_14_1;
  assign t_r15_c2_6 = t_r15_c2_1 + p_14_3;
  assign t_r15_c2_7 = t_r15_c2_2 + t_r15_c2_3;
  assign t_r15_c2_8 = t_r15_c2_4 + p_16_1;
  assign t_r15_c2_9 = t_r15_c2_5 + t_r15_c2_6;
  assign t_r15_c2_10 = t_r15_c2_7 + t_r15_c2_8;
  assign t_r15_c2_11 = t_r15_c2_9 + t_r15_c2_10;
  assign t_r15_c2_12 = t_r15_c2_11 + p_16_3;
  assign out_15_2 = t_r15_c2_12 >> 4;

  assign t_r15_c3_0 = p_14_3 << 1;
  assign t_r15_c3_1 = p_15_2 << 1;
  assign t_r15_c3_2 = p_15_3 << 2;
  assign t_r15_c3_3 = p_15_4 << 1;
  assign t_r15_c3_4 = p_16_3 << 1;
  assign t_r15_c3_5 = t_r15_c3_0 + p_14_2;
  assign t_r15_c3_6 = t_r15_c3_1 + p_14_4;
  assign t_r15_c3_7 = t_r15_c3_2 + t_r15_c3_3;
  assign t_r15_c3_8 = t_r15_c3_4 + p_16_2;
  assign t_r15_c3_9 = t_r15_c3_5 + t_r15_c3_6;
  assign t_r15_c3_10 = t_r15_c3_7 + t_r15_c3_8;
  assign t_r15_c3_11 = t_r15_c3_9 + t_r15_c3_10;
  assign t_r15_c3_12 = t_r15_c3_11 + p_16_4;
  assign out_15_3 = t_r15_c3_12 >> 4;

  assign t_r15_c4_0 = p_14_4 << 1;
  assign t_r15_c4_1 = p_15_3 << 1;
  assign t_r15_c4_2 = p_15_4 << 2;
  assign t_r15_c4_3 = p_15_5 << 1;
  assign t_r15_c4_4 = p_16_4 << 1;
  assign t_r15_c4_5 = t_r15_c4_0 + p_14_3;
  assign t_r15_c4_6 = t_r15_c4_1 + p_14_5;
  assign t_r15_c4_7 = t_r15_c4_2 + t_r15_c4_3;
  assign t_r15_c4_8 = t_r15_c4_4 + p_16_3;
  assign t_r15_c4_9 = t_r15_c4_5 + t_r15_c4_6;
  assign t_r15_c4_10 = t_r15_c4_7 + t_r15_c4_8;
  assign t_r15_c4_11 = t_r15_c4_9 + t_r15_c4_10;
  assign t_r15_c4_12 = t_r15_c4_11 + p_16_5;
  assign out_15_4 = t_r15_c4_12 >> 4;

  assign t_r15_c5_0 = p_14_5 << 1;
  assign t_r15_c5_1 = p_15_4 << 1;
  assign t_r15_c5_2 = p_15_5 << 2;
  assign t_r15_c5_3 = p_15_6 << 1;
  assign t_r15_c5_4 = p_16_5 << 1;
  assign t_r15_c5_5 = t_r15_c5_0 + p_14_4;
  assign t_r15_c5_6 = t_r15_c5_1 + p_14_6;
  assign t_r15_c5_7 = t_r15_c5_2 + t_r15_c5_3;
  assign t_r15_c5_8 = t_r15_c5_4 + p_16_4;
  assign t_r15_c5_9 = t_r15_c5_5 + t_r15_c5_6;
  assign t_r15_c5_10 = t_r15_c5_7 + t_r15_c5_8;
  assign t_r15_c5_11 = t_r15_c5_9 + t_r15_c5_10;
  assign t_r15_c5_12 = t_r15_c5_11 + p_16_6;
  assign out_15_5 = t_r15_c5_12 >> 4;

  assign t_r15_c6_0 = p_14_6 << 1;
  assign t_r15_c6_1 = p_15_5 << 1;
  assign t_r15_c6_2 = p_15_6 << 2;
  assign t_r15_c6_3 = p_15_7 << 1;
  assign t_r15_c6_4 = p_16_6 << 1;
  assign t_r15_c6_5 = t_r15_c6_0 + p_14_5;
  assign t_r15_c6_6 = t_r15_c6_1 + p_14_7;
  assign t_r15_c6_7 = t_r15_c6_2 + t_r15_c6_3;
  assign t_r15_c6_8 = t_r15_c6_4 + p_16_5;
  assign t_r15_c6_9 = t_r15_c6_5 + t_r15_c6_6;
  assign t_r15_c6_10 = t_r15_c6_7 + t_r15_c6_8;
  assign t_r15_c6_11 = t_r15_c6_9 + t_r15_c6_10;
  assign t_r15_c6_12 = t_r15_c6_11 + p_16_7;
  assign out_15_6 = t_r15_c6_12 >> 4;

  assign t_r15_c7_0 = p_14_7 << 1;
  assign t_r15_c7_1 = p_15_6 << 1;
  assign t_r15_c7_2 = p_15_7 << 2;
  assign t_r15_c7_3 = p_15_8 << 1;
  assign t_r15_c7_4 = p_16_7 << 1;
  assign t_r15_c7_5 = t_r15_c7_0 + p_14_6;
  assign t_r15_c7_6 = t_r15_c7_1 + p_14_8;
  assign t_r15_c7_7 = t_r15_c7_2 + t_r15_c7_3;
  assign t_r15_c7_8 = t_r15_c7_4 + p_16_6;
  assign t_r15_c7_9 = t_r15_c7_5 + t_r15_c7_6;
  assign t_r15_c7_10 = t_r15_c7_7 + t_r15_c7_8;
  assign t_r15_c7_11 = t_r15_c7_9 + t_r15_c7_10;
  assign t_r15_c7_12 = t_r15_c7_11 + p_16_8;
  assign out_15_7 = t_r15_c7_12 >> 4;

  assign t_r15_c8_0 = p_14_8 << 1;
  assign t_r15_c8_1 = p_15_7 << 1;
  assign t_r15_c8_2 = p_15_8 << 2;
  assign t_r15_c8_3 = p_15_9 << 1;
  assign t_r15_c8_4 = p_16_8 << 1;
  assign t_r15_c8_5 = t_r15_c8_0 + p_14_7;
  assign t_r15_c8_6 = t_r15_c8_1 + p_14_9;
  assign t_r15_c8_7 = t_r15_c8_2 + t_r15_c8_3;
  assign t_r15_c8_8 = t_r15_c8_4 + p_16_7;
  assign t_r15_c8_9 = t_r15_c8_5 + t_r15_c8_6;
  assign t_r15_c8_10 = t_r15_c8_7 + t_r15_c8_8;
  assign t_r15_c8_11 = t_r15_c8_9 + t_r15_c8_10;
  assign t_r15_c8_12 = t_r15_c8_11 + p_16_9;
  assign out_15_8 = t_r15_c8_12 >> 4;

  assign t_r15_c9_0 = p_14_9 << 1;
  assign t_r15_c9_1 = p_15_8 << 1;
  assign t_r15_c9_2 = p_15_9 << 2;
  assign t_r15_c9_3 = p_15_10 << 1;
  assign t_r15_c9_4 = p_16_9 << 1;
  assign t_r15_c9_5 = t_r15_c9_0 + p_14_8;
  assign t_r15_c9_6 = t_r15_c9_1 + p_14_10;
  assign t_r15_c9_7 = t_r15_c9_2 + t_r15_c9_3;
  assign t_r15_c9_8 = t_r15_c9_4 + p_16_8;
  assign t_r15_c9_9 = t_r15_c9_5 + t_r15_c9_6;
  assign t_r15_c9_10 = t_r15_c9_7 + t_r15_c9_8;
  assign t_r15_c9_11 = t_r15_c9_9 + t_r15_c9_10;
  assign t_r15_c9_12 = t_r15_c9_11 + p_16_10;
  assign out_15_9 = t_r15_c9_12 >> 4;

  assign t_r15_c10_0 = p_14_10 << 1;
  assign t_r15_c10_1 = p_15_9 << 1;
  assign t_r15_c10_2 = p_15_10 << 2;
  assign t_r15_c10_3 = p_15_11 << 1;
  assign t_r15_c10_4 = p_16_10 << 1;
  assign t_r15_c10_5 = t_r15_c10_0 + p_14_9;
  assign t_r15_c10_6 = t_r15_c10_1 + p_14_11;
  assign t_r15_c10_7 = t_r15_c10_2 + t_r15_c10_3;
  assign t_r15_c10_8 = t_r15_c10_4 + p_16_9;
  assign t_r15_c10_9 = t_r15_c10_5 + t_r15_c10_6;
  assign t_r15_c10_10 = t_r15_c10_7 + t_r15_c10_8;
  assign t_r15_c10_11 = t_r15_c10_9 + t_r15_c10_10;
  assign t_r15_c10_12 = t_r15_c10_11 + p_16_11;
  assign out_15_10 = t_r15_c10_12 >> 4;

  assign t_r15_c11_0 = p_14_11 << 1;
  assign t_r15_c11_1 = p_15_10 << 1;
  assign t_r15_c11_2 = p_15_11 << 2;
  assign t_r15_c11_3 = p_15_12 << 1;
  assign t_r15_c11_4 = p_16_11 << 1;
  assign t_r15_c11_5 = t_r15_c11_0 + p_14_10;
  assign t_r15_c11_6 = t_r15_c11_1 + p_14_12;
  assign t_r15_c11_7 = t_r15_c11_2 + t_r15_c11_3;
  assign t_r15_c11_8 = t_r15_c11_4 + p_16_10;
  assign t_r15_c11_9 = t_r15_c11_5 + t_r15_c11_6;
  assign t_r15_c11_10 = t_r15_c11_7 + t_r15_c11_8;
  assign t_r15_c11_11 = t_r15_c11_9 + t_r15_c11_10;
  assign t_r15_c11_12 = t_r15_c11_11 + p_16_12;
  assign out_15_11 = t_r15_c11_12 >> 4;

  assign t_r15_c12_0 = p_14_12 << 1;
  assign t_r15_c12_1 = p_15_11 << 1;
  assign t_r15_c12_2 = p_15_12 << 2;
  assign t_r15_c12_3 = p_15_13 << 1;
  assign t_r15_c12_4 = p_16_12 << 1;
  assign t_r15_c12_5 = t_r15_c12_0 + p_14_11;
  assign t_r15_c12_6 = t_r15_c12_1 + p_14_13;
  assign t_r15_c12_7 = t_r15_c12_2 + t_r15_c12_3;
  assign t_r15_c12_8 = t_r15_c12_4 + p_16_11;
  assign t_r15_c12_9 = t_r15_c12_5 + t_r15_c12_6;
  assign t_r15_c12_10 = t_r15_c12_7 + t_r15_c12_8;
  assign t_r15_c12_11 = t_r15_c12_9 + t_r15_c12_10;
  assign t_r15_c12_12 = t_r15_c12_11 + p_16_13;
  assign out_15_12 = t_r15_c12_12 >> 4;

  assign t_r15_c13_0 = p_14_13 << 1;
  assign t_r15_c13_1 = p_15_12 << 1;
  assign t_r15_c13_2 = p_15_13 << 2;
  assign t_r15_c13_3 = p_15_14 << 1;
  assign t_r15_c13_4 = p_16_13 << 1;
  assign t_r15_c13_5 = t_r15_c13_0 + p_14_12;
  assign t_r15_c13_6 = t_r15_c13_1 + p_14_14;
  assign t_r15_c13_7 = t_r15_c13_2 + t_r15_c13_3;
  assign t_r15_c13_8 = t_r15_c13_4 + p_16_12;
  assign t_r15_c13_9 = t_r15_c13_5 + t_r15_c13_6;
  assign t_r15_c13_10 = t_r15_c13_7 + t_r15_c13_8;
  assign t_r15_c13_11 = t_r15_c13_9 + t_r15_c13_10;
  assign t_r15_c13_12 = t_r15_c13_11 + p_16_14;
  assign out_15_13 = t_r15_c13_12 >> 4;

  assign t_r15_c14_0 = p_14_14 << 1;
  assign t_r15_c14_1 = p_15_13 << 1;
  assign t_r15_c14_2 = p_15_14 << 2;
  assign t_r15_c14_3 = p_15_15 << 1;
  assign t_r15_c14_4 = p_16_14 << 1;
  assign t_r15_c14_5 = t_r15_c14_0 + p_14_13;
  assign t_r15_c14_6 = t_r15_c14_1 + p_14_15;
  assign t_r15_c14_7 = t_r15_c14_2 + t_r15_c14_3;
  assign t_r15_c14_8 = t_r15_c14_4 + p_16_13;
  assign t_r15_c14_9 = t_r15_c14_5 + t_r15_c14_6;
  assign t_r15_c14_10 = t_r15_c14_7 + t_r15_c14_8;
  assign t_r15_c14_11 = t_r15_c14_9 + t_r15_c14_10;
  assign t_r15_c14_12 = t_r15_c14_11 + p_16_15;
  assign out_15_14 = t_r15_c14_12 >> 4;

  assign t_r15_c15_0 = p_14_15 << 1;
  assign t_r15_c15_1 = p_15_14 << 1;
  assign t_r15_c15_2 = p_15_15 << 2;
  assign t_r15_c15_3 = p_15_16 << 1;
  assign t_r15_c15_4 = p_16_15 << 1;
  assign t_r15_c15_5 = t_r15_c15_0 + p_14_14;
  assign t_r15_c15_6 = t_r15_c15_1 + p_14_16;
  assign t_r15_c15_7 = t_r15_c15_2 + t_r15_c15_3;
  assign t_r15_c15_8 = t_r15_c15_4 + p_16_14;
  assign t_r15_c15_9 = t_r15_c15_5 + t_r15_c15_6;
  assign t_r15_c15_10 = t_r15_c15_7 + t_r15_c15_8;
  assign t_r15_c15_11 = t_r15_c15_9 + t_r15_c15_10;
  assign t_r15_c15_12 = t_r15_c15_11 + p_16_16;
  assign out_15_15 = t_r15_c15_12 >> 4;

  assign t_r15_c16_0 = p_14_16 << 1;
  assign t_r15_c16_1 = p_15_15 << 1;
  assign t_r15_c16_2 = p_15_16 << 2;
  assign t_r15_c16_3 = p_15_17 << 1;
  assign t_r15_c16_4 = p_16_16 << 1;
  assign t_r15_c16_5 = t_r15_c16_0 + p_14_15;
  assign t_r15_c16_6 = t_r15_c16_1 + p_14_17;
  assign t_r15_c16_7 = t_r15_c16_2 + t_r15_c16_3;
  assign t_r15_c16_8 = t_r15_c16_4 + p_16_15;
  assign t_r15_c16_9 = t_r15_c16_5 + t_r15_c16_6;
  assign t_r15_c16_10 = t_r15_c16_7 + t_r15_c16_8;
  assign t_r15_c16_11 = t_r15_c16_9 + t_r15_c16_10;
  assign t_r15_c16_12 = t_r15_c16_11 + p_16_17;
  assign out_15_16 = t_r15_c16_12 >> 4;

  assign t_r15_c17_0 = p_14_17 << 1;
  assign t_r15_c17_1 = p_15_16 << 1;
  assign t_r15_c17_2 = p_15_17 << 2;
  assign t_r15_c17_3 = p_15_18 << 1;
  assign t_r15_c17_4 = p_16_17 << 1;
  assign t_r15_c17_5 = t_r15_c17_0 + p_14_16;
  assign t_r15_c17_6 = t_r15_c17_1 + p_14_18;
  assign t_r15_c17_7 = t_r15_c17_2 + t_r15_c17_3;
  assign t_r15_c17_8 = t_r15_c17_4 + p_16_16;
  assign t_r15_c17_9 = t_r15_c17_5 + t_r15_c17_6;
  assign t_r15_c17_10 = t_r15_c17_7 + t_r15_c17_8;
  assign t_r15_c17_11 = t_r15_c17_9 + t_r15_c17_10;
  assign t_r15_c17_12 = t_r15_c17_11 + p_16_18;
  assign out_15_17 = t_r15_c17_12 >> 4;

  assign t_r15_c18_0 = p_14_18 << 1;
  assign t_r15_c18_1 = p_15_17 << 1;
  assign t_r15_c18_2 = p_15_18 << 2;
  assign t_r15_c18_3 = p_15_19 << 1;
  assign t_r15_c18_4 = p_16_18 << 1;
  assign t_r15_c18_5 = t_r15_c18_0 + p_14_17;
  assign t_r15_c18_6 = t_r15_c18_1 + p_14_19;
  assign t_r15_c18_7 = t_r15_c18_2 + t_r15_c18_3;
  assign t_r15_c18_8 = t_r15_c18_4 + p_16_17;
  assign t_r15_c18_9 = t_r15_c18_5 + t_r15_c18_6;
  assign t_r15_c18_10 = t_r15_c18_7 + t_r15_c18_8;
  assign t_r15_c18_11 = t_r15_c18_9 + t_r15_c18_10;
  assign t_r15_c18_12 = t_r15_c18_11 + p_16_19;
  assign out_15_18 = t_r15_c18_12 >> 4;

  assign t_r15_c19_0 = p_14_19 << 1;
  assign t_r15_c19_1 = p_15_18 << 1;
  assign t_r15_c19_2 = p_15_19 << 2;
  assign t_r15_c19_3 = p_15_20 << 1;
  assign t_r15_c19_4 = p_16_19 << 1;
  assign t_r15_c19_5 = t_r15_c19_0 + p_14_18;
  assign t_r15_c19_6 = t_r15_c19_1 + p_14_20;
  assign t_r15_c19_7 = t_r15_c19_2 + t_r15_c19_3;
  assign t_r15_c19_8 = t_r15_c19_4 + p_16_18;
  assign t_r15_c19_9 = t_r15_c19_5 + t_r15_c19_6;
  assign t_r15_c19_10 = t_r15_c19_7 + t_r15_c19_8;
  assign t_r15_c19_11 = t_r15_c19_9 + t_r15_c19_10;
  assign t_r15_c19_12 = t_r15_c19_11 + p_16_20;
  assign out_15_19 = t_r15_c19_12 >> 4;

  assign t_r15_c20_0 = p_14_20 << 1;
  assign t_r15_c20_1 = p_15_19 << 1;
  assign t_r15_c20_2 = p_15_20 << 2;
  assign t_r15_c20_3 = p_15_21 << 1;
  assign t_r15_c20_4 = p_16_20 << 1;
  assign t_r15_c20_5 = t_r15_c20_0 + p_14_19;
  assign t_r15_c20_6 = t_r15_c20_1 + p_14_21;
  assign t_r15_c20_7 = t_r15_c20_2 + t_r15_c20_3;
  assign t_r15_c20_8 = t_r15_c20_4 + p_16_19;
  assign t_r15_c20_9 = t_r15_c20_5 + t_r15_c20_6;
  assign t_r15_c20_10 = t_r15_c20_7 + t_r15_c20_8;
  assign t_r15_c20_11 = t_r15_c20_9 + t_r15_c20_10;
  assign t_r15_c20_12 = t_r15_c20_11 + p_16_21;
  assign out_15_20 = t_r15_c20_12 >> 4;

  assign t_r15_c21_0 = p_14_21 << 1;
  assign t_r15_c21_1 = p_15_20 << 1;
  assign t_r15_c21_2 = p_15_21 << 2;
  assign t_r15_c21_3 = p_15_22 << 1;
  assign t_r15_c21_4 = p_16_21 << 1;
  assign t_r15_c21_5 = t_r15_c21_0 + p_14_20;
  assign t_r15_c21_6 = t_r15_c21_1 + p_14_22;
  assign t_r15_c21_7 = t_r15_c21_2 + t_r15_c21_3;
  assign t_r15_c21_8 = t_r15_c21_4 + p_16_20;
  assign t_r15_c21_9 = t_r15_c21_5 + t_r15_c21_6;
  assign t_r15_c21_10 = t_r15_c21_7 + t_r15_c21_8;
  assign t_r15_c21_11 = t_r15_c21_9 + t_r15_c21_10;
  assign t_r15_c21_12 = t_r15_c21_11 + p_16_22;
  assign out_15_21 = t_r15_c21_12 >> 4;

  assign t_r15_c22_0 = p_14_22 << 1;
  assign t_r15_c22_1 = p_15_21 << 1;
  assign t_r15_c22_2 = p_15_22 << 2;
  assign t_r15_c22_3 = p_15_23 << 1;
  assign t_r15_c22_4 = p_16_22 << 1;
  assign t_r15_c22_5 = t_r15_c22_0 + p_14_21;
  assign t_r15_c22_6 = t_r15_c22_1 + p_14_23;
  assign t_r15_c22_7 = t_r15_c22_2 + t_r15_c22_3;
  assign t_r15_c22_8 = t_r15_c22_4 + p_16_21;
  assign t_r15_c22_9 = t_r15_c22_5 + t_r15_c22_6;
  assign t_r15_c22_10 = t_r15_c22_7 + t_r15_c22_8;
  assign t_r15_c22_11 = t_r15_c22_9 + t_r15_c22_10;
  assign t_r15_c22_12 = t_r15_c22_11 + p_16_23;
  assign out_15_22 = t_r15_c22_12 >> 4;

  assign t_r15_c23_0 = p_14_23 << 1;
  assign t_r15_c23_1 = p_15_22 << 1;
  assign t_r15_c23_2 = p_15_23 << 2;
  assign t_r15_c23_3 = p_15_24 << 1;
  assign t_r15_c23_4 = p_16_23 << 1;
  assign t_r15_c23_5 = t_r15_c23_0 + p_14_22;
  assign t_r15_c23_6 = t_r15_c23_1 + p_14_24;
  assign t_r15_c23_7 = t_r15_c23_2 + t_r15_c23_3;
  assign t_r15_c23_8 = t_r15_c23_4 + p_16_22;
  assign t_r15_c23_9 = t_r15_c23_5 + t_r15_c23_6;
  assign t_r15_c23_10 = t_r15_c23_7 + t_r15_c23_8;
  assign t_r15_c23_11 = t_r15_c23_9 + t_r15_c23_10;
  assign t_r15_c23_12 = t_r15_c23_11 + p_16_24;
  assign out_15_23 = t_r15_c23_12 >> 4;

  assign t_r15_c24_0 = p_14_24 << 1;
  assign t_r15_c24_1 = p_15_23 << 1;
  assign t_r15_c24_2 = p_15_24 << 2;
  assign t_r15_c24_3 = p_15_25 << 1;
  assign t_r15_c24_4 = p_16_24 << 1;
  assign t_r15_c24_5 = t_r15_c24_0 + p_14_23;
  assign t_r15_c24_6 = t_r15_c24_1 + p_14_25;
  assign t_r15_c24_7 = t_r15_c24_2 + t_r15_c24_3;
  assign t_r15_c24_8 = t_r15_c24_4 + p_16_23;
  assign t_r15_c24_9 = t_r15_c24_5 + t_r15_c24_6;
  assign t_r15_c24_10 = t_r15_c24_7 + t_r15_c24_8;
  assign t_r15_c24_11 = t_r15_c24_9 + t_r15_c24_10;
  assign t_r15_c24_12 = t_r15_c24_11 + p_16_25;
  assign out_15_24 = t_r15_c24_12 >> 4;

  assign t_r15_c25_0 = p_14_25 << 1;
  assign t_r15_c25_1 = p_15_24 << 1;
  assign t_r15_c25_2 = p_15_25 << 2;
  assign t_r15_c25_3 = p_15_26 << 1;
  assign t_r15_c25_4 = p_16_25 << 1;
  assign t_r15_c25_5 = t_r15_c25_0 + p_14_24;
  assign t_r15_c25_6 = t_r15_c25_1 + p_14_26;
  assign t_r15_c25_7 = t_r15_c25_2 + t_r15_c25_3;
  assign t_r15_c25_8 = t_r15_c25_4 + p_16_24;
  assign t_r15_c25_9 = t_r15_c25_5 + t_r15_c25_6;
  assign t_r15_c25_10 = t_r15_c25_7 + t_r15_c25_8;
  assign t_r15_c25_11 = t_r15_c25_9 + t_r15_c25_10;
  assign t_r15_c25_12 = t_r15_c25_11 + p_16_26;
  assign out_15_25 = t_r15_c25_12 >> 4;

  assign t_r15_c26_0 = p_14_26 << 1;
  assign t_r15_c26_1 = p_15_25 << 1;
  assign t_r15_c26_2 = p_15_26 << 2;
  assign t_r15_c26_3 = p_15_27 << 1;
  assign t_r15_c26_4 = p_16_26 << 1;
  assign t_r15_c26_5 = t_r15_c26_0 + p_14_25;
  assign t_r15_c26_6 = t_r15_c26_1 + p_14_27;
  assign t_r15_c26_7 = t_r15_c26_2 + t_r15_c26_3;
  assign t_r15_c26_8 = t_r15_c26_4 + p_16_25;
  assign t_r15_c26_9 = t_r15_c26_5 + t_r15_c26_6;
  assign t_r15_c26_10 = t_r15_c26_7 + t_r15_c26_8;
  assign t_r15_c26_11 = t_r15_c26_9 + t_r15_c26_10;
  assign t_r15_c26_12 = t_r15_c26_11 + p_16_27;
  assign out_15_26 = t_r15_c26_12 >> 4;

  assign t_r15_c27_0 = p_14_27 << 1;
  assign t_r15_c27_1 = p_15_26 << 1;
  assign t_r15_c27_2 = p_15_27 << 2;
  assign t_r15_c27_3 = p_15_28 << 1;
  assign t_r15_c27_4 = p_16_27 << 1;
  assign t_r15_c27_5 = t_r15_c27_0 + p_14_26;
  assign t_r15_c27_6 = t_r15_c27_1 + p_14_28;
  assign t_r15_c27_7 = t_r15_c27_2 + t_r15_c27_3;
  assign t_r15_c27_8 = t_r15_c27_4 + p_16_26;
  assign t_r15_c27_9 = t_r15_c27_5 + t_r15_c27_6;
  assign t_r15_c27_10 = t_r15_c27_7 + t_r15_c27_8;
  assign t_r15_c27_11 = t_r15_c27_9 + t_r15_c27_10;
  assign t_r15_c27_12 = t_r15_c27_11 + p_16_28;
  assign out_15_27 = t_r15_c27_12 >> 4;

  assign t_r15_c28_0 = p_14_28 << 1;
  assign t_r15_c28_1 = p_15_27 << 1;
  assign t_r15_c28_2 = p_15_28 << 2;
  assign t_r15_c28_3 = p_15_29 << 1;
  assign t_r15_c28_4 = p_16_28 << 1;
  assign t_r15_c28_5 = t_r15_c28_0 + p_14_27;
  assign t_r15_c28_6 = t_r15_c28_1 + p_14_29;
  assign t_r15_c28_7 = t_r15_c28_2 + t_r15_c28_3;
  assign t_r15_c28_8 = t_r15_c28_4 + p_16_27;
  assign t_r15_c28_9 = t_r15_c28_5 + t_r15_c28_6;
  assign t_r15_c28_10 = t_r15_c28_7 + t_r15_c28_8;
  assign t_r15_c28_11 = t_r15_c28_9 + t_r15_c28_10;
  assign t_r15_c28_12 = t_r15_c28_11 + p_16_29;
  assign out_15_28 = t_r15_c28_12 >> 4;

  assign t_r15_c29_0 = p_14_29 << 1;
  assign t_r15_c29_1 = p_15_28 << 1;
  assign t_r15_c29_2 = p_15_29 << 2;
  assign t_r15_c29_3 = p_15_30 << 1;
  assign t_r15_c29_4 = p_16_29 << 1;
  assign t_r15_c29_5 = t_r15_c29_0 + p_14_28;
  assign t_r15_c29_6 = t_r15_c29_1 + p_14_30;
  assign t_r15_c29_7 = t_r15_c29_2 + t_r15_c29_3;
  assign t_r15_c29_8 = t_r15_c29_4 + p_16_28;
  assign t_r15_c29_9 = t_r15_c29_5 + t_r15_c29_6;
  assign t_r15_c29_10 = t_r15_c29_7 + t_r15_c29_8;
  assign t_r15_c29_11 = t_r15_c29_9 + t_r15_c29_10;
  assign t_r15_c29_12 = t_r15_c29_11 + p_16_30;
  assign out_15_29 = t_r15_c29_12 >> 4;

  assign t_r15_c30_0 = p_14_30 << 1;
  assign t_r15_c30_1 = p_15_29 << 1;
  assign t_r15_c30_2 = p_15_30 << 2;
  assign t_r15_c30_3 = p_15_31 << 1;
  assign t_r15_c30_4 = p_16_30 << 1;
  assign t_r15_c30_5 = t_r15_c30_0 + p_14_29;
  assign t_r15_c30_6 = t_r15_c30_1 + p_14_31;
  assign t_r15_c30_7 = t_r15_c30_2 + t_r15_c30_3;
  assign t_r15_c30_8 = t_r15_c30_4 + p_16_29;
  assign t_r15_c30_9 = t_r15_c30_5 + t_r15_c30_6;
  assign t_r15_c30_10 = t_r15_c30_7 + t_r15_c30_8;
  assign t_r15_c30_11 = t_r15_c30_9 + t_r15_c30_10;
  assign t_r15_c30_12 = t_r15_c30_11 + p_16_31;
  assign out_15_30 = t_r15_c30_12 >> 4;

  assign t_r15_c31_0 = p_14_31 << 1;
  assign t_r15_c31_1 = p_15_30 << 1;
  assign t_r15_c31_2 = p_15_31 << 2;
  assign t_r15_c31_3 = p_15_32 << 1;
  assign t_r15_c31_4 = p_16_31 << 1;
  assign t_r15_c31_5 = t_r15_c31_0 + p_14_30;
  assign t_r15_c31_6 = t_r15_c31_1 + p_14_32;
  assign t_r15_c31_7 = t_r15_c31_2 + t_r15_c31_3;
  assign t_r15_c31_8 = t_r15_c31_4 + p_16_30;
  assign t_r15_c31_9 = t_r15_c31_5 + t_r15_c31_6;
  assign t_r15_c31_10 = t_r15_c31_7 + t_r15_c31_8;
  assign t_r15_c31_11 = t_r15_c31_9 + t_r15_c31_10;
  assign t_r15_c31_12 = t_r15_c31_11 + p_16_32;
  assign out_15_31 = t_r15_c31_12 >> 4;

  assign t_r15_c32_0 = p_14_32 << 1;
  assign t_r15_c32_1 = p_15_31 << 1;
  assign t_r15_c32_2 = p_15_32 << 2;
  assign t_r15_c32_3 = p_15_33 << 1;
  assign t_r15_c32_4 = p_16_32 << 1;
  assign t_r15_c32_5 = t_r15_c32_0 + p_14_31;
  assign t_r15_c32_6 = t_r15_c32_1 + p_14_33;
  assign t_r15_c32_7 = t_r15_c32_2 + t_r15_c32_3;
  assign t_r15_c32_8 = t_r15_c32_4 + p_16_31;
  assign t_r15_c32_9 = t_r15_c32_5 + t_r15_c32_6;
  assign t_r15_c32_10 = t_r15_c32_7 + t_r15_c32_8;
  assign t_r15_c32_11 = t_r15_c32_9 + t_r15_c32_10;
  assign t_r15_c32_12 = t_r15_c32_11 + p_16_33;
  assign out_15_32 = t_r15_c32_12 >> 4;

  assign t_r15_c33_0 = p_14_33 << 1;
  assign t_r15_c33_1 = p_15_32 << 1;
  assign t_r15_c33_2 = p_15_33 << 2;
  assign t_r15_c33_3 = p_15_34 << 1;
  assign t_r15_c33_4 = p_16_33 << 1;
  assign t_r15_c33_5 = t_r15_c33_0 + p_14_32;
  assign t_r15_c33_6 = t_r15_c33_1 + p_14_34;
  assign t_r15_c33_7 = t_r15_c33_2 + t_r15_c33_3;
  assign t_r15_c33_8 = t_r15_c33_4 + p_16_32;
  assign t_r15_c33_9 = t_r15_c33_5 + t_r15_c33_6;
  assign t_r15_c33_10 = t_r15_c33_7 + t_r15_c33_8;
  assign t_r15_c33_11 = t_r15_c33_9 + t_r15_c33_10;
  assign t_r15_c33_12 = t_r15_c33_11 + p_16_34;
  assign out_15_33 = t_r15_c33_12 >> 4;

  assign t_r15_c34_0 = p_14_34 << 1;
  assign t_r15_c34_1 = p_15_33 << 1;
  assign t_r15_c34_2 = p_15_34 << 2;
  assign t_r15_c34_3 = p_15_35 << 1;
  assign t_r15_c34_4 = p_16_34 << 1;
  assign t_r15_c34_5 = t_r15_c34_0 + p_14_33;
  assign t_r15_c34_6 = t_r15_c34_1 + p_14_35;
  assign t_r15_c34_7 = t_r15_c34_2 + t_r15_c34_3;
  assign t_r15_c34_8 = t_r15_c34_4 + p_16_33;
  assign t_r15_c34_9 = t_r15_c34_5 + t_r15_c34_6;
  assign t_r15_c34_10 = t_r15_c34_7 + t_r15_c34_8;
  assign t_r15_c34_11 = t_r15_c34_9 + t_r15_c34_10;
  assign t_r15_c34_12 = t_r15_c34_11 + p_16_35;
  assign out_15_34 = t_r15_c34_12 >> 4;

  assign t_r15_c35_0 = p_14_35 << 1;
  assign t_r15_c35_1 = p_15_34 << 1;
  assign t_r15_c35_2 = p_15_35 << 2;
  assign t_r15_c35_3 = p_15_36 << 1;
  assign t_r15_c35_4 = p_16_35 << 1;
  assign t_r15_c35_5 = t_r15_c35_0 + p_14_34;
  assign t_r15_c35_6 = t_r15_c35_1 + p_14_36;
  assign t_r15_c35_7 = t_r15_c35_2 + t_r15_c35_3;
  assign t_r15_c35_8 = t_r15_c35_4 + p_16_34;
  assign t_r15_c35_9 = t_r15_c35_5 + t_r15_c35_6;
  assign t_r15_c35_10 = t_r15_c35_7 + t_r15_c35_8;
  assign t_r15_c35_11 = t_r15_c35_9 + t_r15_c35_10;
  assign t_r15_c35_12 = t_r15_c35_11 + p_16_36;
  assign out_15_35 = t_r15_c35_12 >> 4;

  assign t_r15_c36_0 = p_14_36 << 1;
  assign t_r15_c36_1 = p_15_35 << 1;
  assign t_r15_c36_2 = p_15_36 << 2;
  assign t_r15_c36_3 = p_15_37 << 1;
  assign t_r15_c36_4 = p_16_36 << 1;
  assign t_r15_c36_5 = t_r15_c36_0 + p_14_35;
  assign t_r15_c36_6 = t_r15_c36_1 + p_14_37;
  assign t_r15_c36_7 = t_r15_c36_2 + t_r15_c36_3;
  assign t_r15_c36_8 = t_r15_c36_4 + p_16_35;
  assign t_r15_c36_9 = t_r15_c36_5 + t_r15_c36_6;
  assign t_r15_c36_10 = t_r15_c36_7 + t_r15_c36_8;
  assign t_r15_c36_11 = t_r15_c36_9 + t_r15_c36_10;
  assign t_r15_c36_12 = t_r15_c36_11 + p_16_37;
  assign out_15_36 = t_r15_c36_12 >> 4;

  assign t_r15_c37_0 = p_14_37 << 1;
  assign t_r15_c37_1 = p_15_36 << 1;
  assign t_r15_c37_2 = p_15_37 << 2;
  assign t_r15_c37_3 = p_15_38 << 1;
  assign t_r15_c37_4 = p_16_37 << 1;
  assign t_r15_c37_5 = t_r15_c37_0 + p_14_36;
  assign t_r15_c37_6 = t_r15_c37_1 + p_14_38;
  assign t_r15_c37_7 = t_r15_c37_2 + t_r15_c37_3;
  assign t_r15_c37_8 = t_r15_c37_4 + p_16_36;
  assign t_r15_c37_9 = t_r15_c37_5 + t_r15_c37_6;
  assign t_r15_c37_10 = t_r15_c37_7 + t_r15_c37_8;
  assign t_r15_c37_11 = t_r15_c37_9 + t_r15_c37_10;
  assign t_r15_c37_12 = t_r15_c37_11 + p_16_38;
  assign out_15_37 = t_r15_c37_12 >> 4;

  assign t_r15_c38_0 = p_14_38 << 1;
  assign t_r15_c38_1 = p_15_37 << 1;
  assign t_r15_c38_2 = p_15_38 << 2;
  assign t_r15_c38_3 = p_15_39 << 1;
  assign t_r15_c38_4 = p_16_38 << 1;
  assign t_r15_c38_5 = t_r15_c38_0 + p_14_37;
  assign t_r15_c38_6 = t_r15_c38_1 + p_14_39;
  assign t_r15_c38_7 = t_r15_c38_2 + t_r15_c38_3;
  assign t_r15_c38_8 = t_r15_c38_4 + p_16_37;
  assign t_r15_c38_9 = t_r15_c38_5 + t_r15_c38_6;
  assign t_r15_c38_10 = t_r15_c38_7 + t_r15_c38_8;
  assign t_r15_c38_11 = t_r15_c38_9 + t_r15_c38_10;
  assign t_r15_c38_12 = t_r15_c38_11 + p_16_39;
  assign out_15_38 = t_r15_c38_12 >> 4;

  assign t_r15_c39_0 = p_14_39 << 1;
  assign t_r15_c39_1 = p_15_38 << 1;
  assign t_r15_c39_2 = p_15_39 << 2;
  assign t_r15_c39_3 = p_15_40 << 1;
  assign t_r15_c39_4 = p_16_39 << 1;
  assign t_r15_c39_5 = t_r15_c39_0 + p_14_38;
  assign t_r15_c39_6 = t_r15_c39_1 + p_14_40;
  assign t_r15_c39_7 = t_r15_c39_2 + t_r15_c39_3;
  assign t_r15_c39_8 = t_r15_c39_4 + p_16_38;
  assign t_r15_c39_9 = t_r15_c39_5 + t_r15_c39_6;
  assign t_r15_c39_10 = t_r15_c39_7 + t_r15_c39_8;
  assign t_r15_c39_11 = t_r15_c39_9 + t_r15_c39_10;
  assign t_r15_c39_12 = t_r15_c39_11 + p_16_40;
  assign out_15_39 = t_r15_c39_12 >> 4;

  assign t_r15_c40_0 = p_14_40 << 1;
  assign t_r15_c40_1 = p_15_39 << 1;
  assign t_r15_c40_2 = p_15_40 << 2;
  assign t_r15_c40_3 = p_15_41 << 1;
  assign t_r15_c40_4 = p_16_40 << 1;
  assign t_r15_c40_5 = t_r15_c40_0 + p_14_39;
  assign t_r15_c40_6 = t_r15_c40_1 + p_14_41;
  assign t_r15_c40_7 = t_r15_c40_2 + t_r15_c40_3;
  assign t_r15_c40_8 = t_r15_c40_4 + p_16_39;
  assign t_r15_c40_9 = t_r15_c40_5 + t_r15_c40_6;
  assign t_r15_c40_10 = t_r15_c40_7 + t_r15_c40_8;
  assign t_r15_c40_11 = t_r15_c40_9 + t_r15_c40_10;
  assign t_r15_c40_12 = t_r15_c40_11 + p_16_41;
  assign out_15_40 = t_r15_c40_12 >> 4;

  assign t_r15_c41_0 = p_14_41 << 1;
  assign t_r15_c41_1 = p_15_40 << 1;
  assign t_r15_c41_2 = p_15_41 << 2;
  assign t_r15_c41_3 = p_15_42 << 1;
  assign t_r15_c41_4 = p_16_41 << 1;
  assign t_r15_c41_5 = t_r15_c41_0 + p_14_40;
  assign t_r15_c41_6 = t_r15_c41_1 + p_14_42;
  assign t_r15_c41_7 = t_r15_c41_2 + t_r15_c41_3;
  assign t_r15_c41_8 = t_r15_c41_4 + p_16_40;
  assign t_r15_c41_9 = t_r15_c41_5 + t_r15_c41_6;
  assign t_r15_c41_10 = t_r15_c41_7 + t_r15_c41_8;
  assign t_r15_c41_11 = t_r15_c41_9 + t_r15_c41_10;
  assign t_r15_c41_12 = t_r15_c41_11 + p_16_42;
  assign out_15_41 = t_r15_c41_12 >> 4;

  assign t_r15_c42_0 = p_14_42 << 1;
  assign t_r15_c42_1 = p_15_41 << 1;
  assign t_r15_c42_2 = p_15_42 << 2;
  assign t_r15_c42_3 = p_15_43 << 1;
  assign t_r15_c42_4 = p_16_42 << 1;
  assign t_r15_c42_5 = t_r15_c42_0 + p_14_41;
  assign t_r15_c42_6 = t_r15_c42_1 + p_14_43;
  assign t_r15_c42_7 = t_r15_c42_2 + t_r15_c42_3;
  assign t_r15_c42_8 = t_r15_c42_4 + p_16_41;
  assign t_r15_c42_9 = t_r15_c42_5 + t_r15_c42_6;
  assign t_r15_c42_10 = t_r15_c42_7 + t_r15_c42_8;
  assign t_r15_c42_11 = t_r15_c42_9 + t_r15_c42_10;
  assign t_r15_c42_12 = t_r15_c42_11 + p_16_43;
  assign out_15_42 = t_r15_c42_12 >> 4;

  assign t_r15_c43_0 = p_14_43 << 1;
  assign t_r15_c43_1 = p_15_42 << 1;
  assign t_r15_c43_2 = p_15_43 << 2;
  assign t_r15_c43_3 = p_15_44 << 1;
  assign t_r15_c43_4 = p_16_43 << 1;
  assign t_r15_c43_5 = t_r15_c43_0 + p_14_42;
  assign t_r15_c43_6 = t_r15_c43_1 + p_14_44;
  assign t_r15_c43_7 = t_r15_c43_2 + t_r15_c43_3;
  assign t_r15_c43_8 = t_r15_c43_4 + p_16_42;
  assign t_r15_c43_9 = t_r15_c43_5 + t_r15_c43_6;
  assign t_r15_c43_10 = t_r15_c43_7 + t_r15_c43_8;
  assign t_r15_c43_11 = t_r15_c43_9 + t_r15_c43_10;
  assign t_r15_c43_12 = t_r15_c43_11 + p_16_44;
  assign out_15_43 = t_r15_c43_12 >> 4;

  assign t_r15_c44_0 = p_14_44 << 1;
  assign t_r15_c44_1 = p_15_43 << 1;
  assign t_r15_c44_2 = p_15_44 << 2;
  assign t_r15_c44_3 = p_15_45 << 1;
  assign t_r15_c44_4 = p_16_44 << 1;
  assign t_r15_c44_5 = t_r15_c44_0 + p_14_43;
  assign t_r15_c44_6 = t_r15_c44_1 + p_14_45;
  assign t_r15_c44_7 = t_r15_c44_2 + t_r15_c44_3;
  assign t_r15_c44_8 = t_r15_c44_4 + p_16_43;
  assign t_r15_c44_9 = t_r15_c44_5 + t_r15_c44_6;
  assign t_r15_c44_10 = t_r15_c44_7 + t_r15_c44_8;
  assign t_r15_c44_11 = t_r15_c44_9 + t_r15_c44_10;
  assign t_r15_c44_12 = t_r15_c44_11 + p_16_45;
  assign out_15_44 = t_r15_c44_12 >> 4;

  assign t_r15_c45_0 = p_14_45 << 1;
  assign t_r15_c45_1 = p_15_44 << 1;
  assign t_r15_c45_2 = p_15_45 << 2;
  assign t_r15_c45_3 = p_15_46 << 1;
  assign t_r15_c45_4 = p_16_45 << 1;
  assign t_r15_c45_5 = t_r15_c45_0 + p_14_44;
  assign t_r15_c45_6 = t_r15_c45_1 + p_14_46;
  assign t_r15_c45_7 = t_r15_c45_2 + t_r15_c45_3;
  assign t_r15_c45_8 = t_r15_c45_4 + p_16_44;
  assign t_r15_c45_9 = t_r15_c45_5 + t_r15_c45_6;
  assign t_r15_c45_10 = t_r15_c45_7 + t_r15_c45_8;
  assign t_r15_c45_11 = t_r15_c45_9 + t_r15_c45_10;
  assign t_r15_c45_12 = t_r15_c45_11 + p_16_46;
  assign out_15_45 = t_r15_c45_12 >> 4;

  assign t_r15_c46_0 = p_14_46 << 1;
  assign t_r15_c46_1 = p_15_45 << 1;
  assign t_r15_c46_2 = p_15_46 << 2;
  assign t_r15_c46_3 = p_15_47 << 1;
  assign t_r15_c46_4 = p_16_46 << 1;
  assign t_r15_c46_5 = t_r15_c46_0 + p_14_45;
  assign t_r15_c46_6 = t_r15_c46_1 + p_14_47;
  assign t_r15_c46_7 = t_r15_c46_2 + t_r15_c46_3;
  assign t_r15_c46_8 = t_r15_c46_4 + p_16_45;
  assign t_r15_c46_9 = t_r15_c46_5 + t_r15_c46_6;
  assign t_r15_c46_10 = t_r15_c46_7 + t_r15_c46_8;
  assign t_r15_c46_11 = t_r15_c46_9 + t_r15_c46_10;
  assign t_r15_c46_12 = t_r15_c46_11 + p_16_47;
  assign out_15_46 = t_r15_c46_12 >> 4;

  assign t_r15_c47_0 = p_14_47 << 1;
  assign t_r15_c47_1 = p_15_46 << 1;
  assign t_r15_c47_2 = p_15_47 << 2;
  assign t_r15_c47_3 = p_15_48 << 1;
  assign t_r15_c47_4 = p_16_47 << 1;
  assign t_r15_c47_5 = t_r15_c47_0 + p_14_46;
  assign t_r15_c47_6 = t_r15_c47_1 + p_14_48;
  assign t_r15_c47_7 = t_r15_c47_2 + t_r15_c47_3;
  assign t_r15_c47_8 = t_r15_c47_4 + p_16_46;
  assign t_r15_c47_9 = t_r15_c47_5 + t_r15_c47_6;
  assign t_r15_c47_10 = t_r15_c47_7 + t_r15_c47_8;
  assign t_r15_c47_11 = t_r15_c47_9 + t_r15_c47_10;
  assign t_r15_c47_12 = t_r15_c47_11 + p_16_48;
  assign out_15_47 = t_r15_c47_12 >> 4;

  assign t_r15_c48_0 = p_14_48 << 1;
  assign t_r15_c48_1 = p_15_47 << 1;
  assign t_r15_c48_2 = p_15_48 << 2;
  assign t_r15_c48_3 = p_15_49 << 1;
  assign t_r15_c48_4 = p_16_48 << 1;
  assign t_r15_c48_5 = t_r15_c48_0 + p_14_47;
  assign t_r15_c48_6 = t_r15_c48_1 + p_14_49;
  assign t_r15_c48_7 = t_r15_c48_2 + t_r15_c48_3;
  assign t_r15_c48_8 = t_r15_c48_4 + p_16_47;
  assign t_r15_c48_9 = t_r15_c48_5 + t_r15_c48_6;
  assign t_r15_c48_10 = t_r15_c48_7 + t_r15_c48_8;
  assign t_r15_c48_11 = t_r15_c48_9 + t_r15_c48_10;
  assign t_r15_c48_12 = t_r15_c48_11 + p_16_49;
  assign out_15_48 = t_r15_c48_12 >> 4;

  assign t_r15_c49_0 = p_14_49 << 1;
  assign t_r15_c49_1 = p_15_48 << 1;
  assign t_r15_c49_2 = p_15_49 << 2;
  assign t_r15_c49_3 = p_15_50 << 1;
  assign t_r15_c49_4 = p_16_49 << 1;
  assign t_r15_c49_5 = t_r15_c49_0 + p_14_48;
  assign t_r15_c49_6 = t_r15_c49_1 + p_14_50;
  assign t_r15_c49_7 = t_r15_c49_2 + t_r15_c49_3;
  assign t_r15_c49_8 = t_r15_c49_4 + p_16_48;
  assign t_r15_c49_9 = t_r15_c49_5 + t_r15_c49_6;
  assign t_r15_c49_10 = t_r15_c49_7 + t_r15_c49_8;
  assign t_r15_c49_11 = t_r15_c49_9 + t_r15_c49_10;
  assign t_r15_c49_12 = t_r15_c49_11 + p_16_50;
  assign out_15_49 = t_r15_c49_12 >> 4;

  assign t_r15_c50_0 = p_14_50 << 1;
  assign t_r15_c50_1 = p_15_49 << 1;
  assign t_r15_c50_2 = p_15_50 << 2;
  assign t_r15_c50_3 = p_15_51 << 1;
  assign t_r15_c50_4 = p_16_50 << 1;
  assign t_r15_c50_5 = t_r15_c50_0 + p_14_49;
  assign t_r15_c50_6 = t_r15_c50_1 + p_14_51;
  assign t_r15_c50_7 = t_r15_c50_2 + t_r15_c50_3;
  assign t_r15_c50_8 = t_r15_c50_4 + p_16_49;
  assign t_r15_c50_9 = t_r15_c50_5 + t_r15_c50_6;
  assign t_r15_c50_10 = t_r15_c50_7 + t_r15_c50_8;
  assign t_r15_c50_11 = t_r15_c50_9 + t_r15_c50_10;
  assign t_r15_c50_12 = t_r15_c50_11 + p_16_51;
  assign out_15_50 = t_r15_c50_12 >> 4;

  assign t_r15_c51_0 = p_14_51 << 1;
  assign t_r15_c51_1 = p_15_50 << 1;
  assign t_r15_c51_2 = p_15_51 << 2;
  assign t_r15_c51_3 = p_15_52 << 1;
  assign t_r15_c51_4 = p_16_51 << 1;
  assign t_r15_c51_5 = t_r15_c51_0 + p_14_50;
  assign t_r15_c51_6 = t_r15_c51_1 + p_14_52;
  assign t_r15_c51_7 = t_r15_c51_2 + t_r15_c51_3;
  assign t_r15_c51_8 = t_r15_c51_4 + p_16_50;
  assign t_r15_c51_9 = t_r15_c51_5 + t_r15_c51_6;
  assign t_r15_c51_10 = t_r15_c51_7 + t_r15_c51_8;
  assign t_r15_c51_11 = t_r15_c51_9 + t_r15_c51_10;
  assign t_r15_c51_12 = t_r15_c51_11 + p_16_52;
  assign out_15_51 = t_r15_c51_12 >> 4;

  assign t_r15_c52_0 = p_14_52 << 1;
  assign t_r15_c52_1 = p_15_51 << 1;
  assign t_r15_c52_2 = p_15_52 << 2;
  assign t_r15_c52_3 = p_15_53 << 1;
  assign t_r15_c52_4 = p_16_52 << 1;
  assign t_r15_c52_5 = t_r15_c52_0 + p_14_51;
  assign t_r15_c52_6 = t_r15_c52_1 + p_14_53;
  assign t_r15_c52_7 = t_r15_c52_2 + t_r15_c52_3;
  assign t_r15_c52_8 = t_r15_c52_4 + p_16_51;
  assign t_r15_c52_9 = t_r15_c52_5 + t_r15_c52_6;
  assign t_r15_c52_10 = t_r15_c52_7 + t_r15_c52_8;
  assign t_r15_c52_11 = t_r15_c52_9 + t_r15_c52_10;
  assign t_r15_c52_12 = t_r15_c52_11 + p_16_53;
  assign out_15_52 = t_r15_c52_12 >> 4;

  assign t_r15_c53_0 = p_14_53 << 1;
  assign t_r15_c53_1 = p_15_52 << 1;
  assign t_r15_c53_2 = p_15_53 << 2;
  assign t_r15_c53_3 = p_15_54 << 1;
  assign t_r15_c53_4 = p_16_53 << 1;
  assign t_r15_c53_5 = t_r15_c53_0 + p_14_52;
  assign t_r15_c53_6 = t_r15_c53_1 + p_14_54;
  assign t_r15_c53_7 = t_r15_c53_2 + t_r15_c53_3;
  assign t_r15_c53_8 = t_r15_c53_4 + p_16_52;
  assign t_r15_c53_9 = t_r15_c53_5 + t_r15_c53_6;
  assign t_r15_c53_10 = t_r15_c53_7 + t_r15_c53_8;
  assign t_r15_c53_11 = t_r15_c53_9 + t_r15_c53_10;
  assign t_r15_c53_12 = t_r15_c53_11 + p_16_54;
  assign out_15_53 = t_r15_c53_12 >> 4;

  assign t_r15_c54_0 = p_14_54 << 1;
  assign t_r15_c54_1 = p_15_53 << 1;
  assign t_r15_c54_2 = p_15_54 << 2;
  assign t_r15_c54_3 = p_15_55 << 1;
  assign t_r15_c54_4 = p_16_54 << 1;
  assign t_r15_c54_5 = t_r15_c54_0 + p_14_53;
  assign t_r15_c54_6 = t_r15_c54_1 + p_14_55;
  assign t_r15_c54_7 = t_r15_c54_2 + t_r15_c54_3;
  assign t_r15_c54_8 = t_r15_c54_4 + p_16_53;
  assign t_r15_c54_9 = t_r15_c54_5 + t_r15_c54_6;
  assign t_r15_c54_10 = t_r15_c54_7 + t_r15_c54_8;
  assign t_r15_c54_11 = t_r15_c54_9 + t_r15_c54_10;
  assign t_r15_c54_12 = t_r15_c54_11 + p_16_55;
  assign out_15_54 = t_r15_c54_12 >> 4;

  assign t_r15_c55_0 = p_14_55 << 1;
  assign t_r15_c55_1 = p_15_54 << 1;
  assign t_r15_c55_2 = p_15_55 << 2;
  assign t_r15_c55_3 = p_15_56 << 1;
  assign t_r15_c55_4 = p_16_55 << 1;
  assign t_r15_c55_5 = t_r15_c55_0 + p_14_54;
  assign t_r15_c55_6 = t_r15_c55_1 + p_14_56;
  assign t_r15_c55_7 = t_r15_c55_2 + t_r15_c55_3;
  assign t_r15_c55_8 = t_r15_c55_4 + p_16_54;
  assign t_r15_c55_9 = t_r15_c55_5 + t_r15_c55_6;
  assign t_r15_c55_10 = t_r15_c55_7 + t_r15_c55_8;
  assign t_r15_c55_11 = t_r15_c55_9 + t_r15_c55_10;
  assign t_r15_c55_12 = t_r15_c55_11 + p_16_56;
  assign out_15_55 = t_r15_c55_12 >> 4;

  assign t_r15_c56_0 = p_14_56 << 1;
  assign t_r15_c56_1 = p_15_55 << 1;
  assign t_r15_c56_2 = p_15_56 << 2;
  assign t_r15_c56_3 = p_15_57 << 1;
  assign t_r15_c56_4 = p_16_56 << 1;
  assign t_r15_c56_5 = t_r15_c56_0 + p_14_55;
  assign t_r15_c56_6 = t_r15_c56_1 + p_14_57;
  assign t_r15_c56_7 = t_r15_c56_2 + t_r15_c56_3;
  assign t_r15_c56_8 = t_r15_c56_4 + p_16_55;
  assign t_r15_c56_9 = t_r15_c56_5 + t_r15_c56_6;
  assign t_r15_c56_10 = t_r15_c56_7 + t_r15_c56_8;
  assign t_r15_c56_11 = t_r15_c56_9 + t_r15_c56_10;
  assign t_r15_c56_12 = t_r15_c56_11 + p_16_57;
  assign out_15_56 = t_r15_c56_12 >> 4;

  assign t_r15_c57_0 = p_14_57 << 1;
  assign t_r15_c57_1 = p_15_56 << 1;
  assign t_r15_c57_2 = p_15_57 << 2;
  assign t_r15_c57_3 = p_15_58 << 1;
  assign t_r15_c57_4 = p_16_57 << 1;
  assign t_r15_c57_5 = t_r15_c57_0 + p_14_56;
  assign t_r15_c57_6 = t_r15_c57_1 + p_14_58;
  assign t_r15_c57_7 = t_r15_c57_2 + t_r15_c57_3;
  assign t_r15_c57_8 = t_r15_c57_4 + p_16_56;
  assign t_r15_c57_9 = t_r15_c57_5 + t_r15_c57_6;
  assign t_r15_c57_10 = t_r15_c57_7 + t_r15_c57_8;
  assign t_r15_c57_11 = t_r15_c57_9 + t_r15_c57_10;
  assign t_r15_c57_12 = t_r15_c57_11 + p_16_58;
  assign out_15_57 = t_r15_c57_12 >> 4;

  assign t_r15_c58_0 = p_14_58 << 1;
  assign t_r15_c58_1 = p_15_57 << 1;
  assign t_r15_c58_2 = p_15_58 << 2;
  assign t_r15_c58_3 = p_15_59 << 1;
  assign t_r15_c58_4 = p_16_58 << 1;
  assign t_r15_c58_5 = t_r15_c58_0 + p_14_57;
  assign t_r15_c58_6 = t_r15_c58_1 + p_14_59;
  assign t_r15_c58_7 = t_r15_c58_2 + t_r15_c58_3;
  assign t_r15_c58_8 = t_r15_c58_4 + p_16_57;
  assign t_r15_c58_9 = t_r15_c58_5 + t_r15_c58_6;
  assign t_r15_c58_10 = t_r15_c58_7 + t_r15_c58_8;
  assign t_r15_c58_11 = t_r15_c58_9 + t_r15_c58_10;
  assign t_r15_c58_12 = t_r15_c58_11 + p_16_59;
  assign out_15_58 = t_r15_c58_12 >> 4;

  assign t_r15_c59_0 = p_14_59 << 1;
  assign t_r15_c59_1 = p_15_58 << 1;
  assign t_r15_c59_2 = p_15_59 << 2;
  assign t_r15_c59_3 = p_15_60 << 1;
  assign t_r15_c59_4 = p_16_59 << 1;
  assign t_r15_c59_5 = t_r15_c59_0 + p_14_58;
  assign t_r15_c59_6 = t_r15_c59_1 + p_14_60;
  assign t_r15_c59_7 = t_r15_c59_2 + t_r15_c59_3;
  assign t_r15_c59_8 = t_r15_c59_4 + p_16_58;
  assign t_r15_c59_9 = t_r15_c59_5 + t_r15_c59_6;
  assign t_r15_c59_10 = t_r15_c59_7 + t_r15_c59_8;
  assign t_r15_c59_11 = t_r15_c59_9 + t_r15_c59_10;
  assign t_r15_c59_12 = t_r15_c59_11 + p_16_60;
  assign out_15_59 = t_r15_c59_12 >> 4;

  assign t_r15_c60_0 = p_14_60 << 1;
  assign t_r15_c60_1 = p_15_59 << 1;
  assign t_r15_c60_2 = p_15_60 << 2;
  assign t_r15_c60_3 = p_15_61 << 1;
  assign t_r15_c60_4 = p_16_60 << 1;
  assign t_r15_c60_5 = t_r15_c60_0 + p_14_59;
  assign t_r15_c60_6 = t_r15_c60_1 + p_14_61;
  assign t_r15_c60_7 = t_r15_c60_2 + t_r15_c60_3;
  assign t_r15_c60_8 = t_r15_c60_4 + p_16_59;
  assign t_r15_c60_9 = t_r15_c60_5 + t_r15_c60_6;
  assign t_r15_c60_10 = t_r15_c60_7 + t_r15_c60_8;
  assign t_r15_c60_11 = t_r15_c60_9 + t_r15_c60_10;
  assign t_r15_c60_12 = t_r15_c60_11 + p_16_61;
  assign out_15_60 = t_r15_c60_12 >> 4;

  assign t_r15_c61_0 = p_14_61 << 1;
  assign t_r15_c61_1 = p_15_60 << 1;
  assign t_r15_c61_2 = p_15_61 << 2;
  assign t_r15_c61_3 = p_15_62 << 1;
  assign t_r15_c61_4 = p_16_61 << 1;
  assign t_r15_c61_5 = t_r15_c61_0 + p_14_60;
  assign t_r15_c61_6 = t_r15_c61_1 + p_14_62;
  assign t_r15_c61_7 = t_r15_c61_2 + t_r15_c61_3;
  assign t_r15_c61_8 = t_r15_c61_4 + p_16_60;
  assign t_r15_c61_9 = t_r15_c61_5 + t_r15_c61_6;
  assign t_r15_c61_10 = t_r15_c61_7 + t_r15_c61_8;
  assign t_r15_c61_11 = t_r15_c61_9 + t_r15_c61_10;
  assign t_r15_c61_12 = t_r15_c61_11 + p_16_62;
  assign out_15_61 = t_r15_c61_12 >> 4;

  assign t_r15_c62_0 = p_14_62 << 1;
  assign t_r15_c62_1 = p_15_61 << 1;
  assign t_r15_c62_2 = p_15_62 << 2;
  assign t_r15_c62_3 = p_15_63 << 1;
  assign t_r15_c62_4 = p_16_62 << 1;
  assign t_r15_c62_5 = t_r15_c62_0 + p_14_61;
  assign t_r15_c62_6 = t_r15_c62_1 + p_14_63;
  assign t_r15_c62_7 = t_r15_c62_2 + t_r15_c62_3;
  assign t_r15_c62_8 = t_r15_c62_4 + p_16_61;
  assign t_r15_c62_9 = t_r15_c62_5 + t_r15_c62_6;
  assign t_r15_c62_10 = t_r15_c62_7 + t_r15_c62_8;
  assign t_r15_c62_11 = t_r15_c62_9 + t_r15_c62_10;
  assign t_r15_c62_12 = t_r15_c62_11 + p_16_63;
  assign out_15_62 = t_r15_c62_12 >> 4;

  assign t_r15_c63_0 = p_14_63 << 1;
  assign t_r15_c63_1 = p_15_62 << 1;
  assign t_r15_c63_2 = p_15_63 << 2;
  assign t_r15_c63_3 = p_15_64 << 1;
  assign t_r15_c63_4 = p_16_63 << 1;
  assign t_r15_c63_5 = t_r15_c63_0 + p_14_62;
  assign t_r15_c63_6 = t_r15_c63_1 + p_14_64;
  assign t_r15_c63_7 = t_r15_c63_2 + t_r15_c63_3;
  assign t_r15_c63_8 = t_r15_c63_4 + p_16_62;
  assign t_r15_c63_9 = t_r15_c63_5 + t_r15_c63_6;
  assign t_r15_c63_10 = t_r15_c63_7 + t_r15_c63_8;
  assign t_r15_c63_11 = t_r15_c63_9 + t_r15_c63_10;
  assign t_r15_c63_12 = t_r15_c63_11 + p_16_64;
  assign out_15_63 = t_r15_c63_12 >> 4;

  assign t_r15_c64_0 = p_14_64 << 1;
  assign t_r15_c64_1 = p_15_63 << 1;
  assign t_r15_c64_2 = p_15_64 << 2;
  assign t_r15_c64_3 = p_15_65 << 1;
  assign t_r15_c64_4 = p_16_64 << 1;
  assign t_r15_c64_5 = t_r15_c64_0 + p_14_63;
  assign t_r15_c64_6 = t_r15_c64_1 + p_14_65;
  assign t_r15_c64_7 = t_r15_c64_2 + t_r15_c64_3;
  assign t_r15_c64_8 = t_r15_c64_4 + p_16_63;
  assign t_r15_c64_9 = t_r15_c64_5 + t_r15_c64_6;
  assign t_r15_c64_10 = t_r15_c64_7 + t_r15_c64_8;
  assign t_r15_c64_11 = t_r15_c64_9 + t_r15_c64_10;
  assign t_r15_c64_12 = t_r15_c64_11 + p_16_65;
  assign out_15_64 = t_r15_c64_12 >> 4;

  assign t_r16_c1_0 = p_15_1 << 1;
  assign t_r16_c1_1 = p_16_0 << 1;
  assign t_r16_c1_2 = p_16_1 << 2;
  assign t_r16_c1_3 = p_16_2 << 1;
  assign t_r16_c1_4 = p_17_1 << 1;
  assign t_r16_c1_5 = t_r16_c1_0 + p_15_0;
  assign t_r16_c1_6 = t_r16_c1_1 + p_15_2;
  assign t_r16_c1_7 = t_r16_c1_2 + t_r16_c1_3;
  assign t_r16_c1_8 = t_r16_c1_4 + p_17_0;
  assign t_r16_c1_9 = t_r16_c1_5 + t_r16_c1_6;
  assign t_r16_c1_10 = t_r16_c1_7 + t_r16_c1_8;
  assign t_r16_c1_11 = t_r16_c1_9 + t_r16_c1_10;
  assign t_r16_c1_12 = t_r16_c1_11 + p_17_2;
  assign out_16_1 = t_r16_c1_12 >> 4;

  assign t_r16_c2_0 = p_15_2 << 1;
  assign t_r16_c2_1 = p_16_1 << 1;
  assign t_r16_c2_2 = p_16_2 << 2;
  assign t_r16_c2_3 = p_16_3 << 1;
  assign t_r16_c2_4 = p_17_2 << 1;
  assign t_r16_c2_5 = t_r16_c2_0 + p_15_1;
  assign t_r16_c2_6 = t_r16_c2_1 + p_15_3;
  assign t_r16_c2_7 = t_r16_c2_2 + t_r16_c2_3;
  assign t_r16_c2_8 = t_r16_c2_4 + p_17_1;
  assign t_r16_c2_9 = t_r16_c2_5 + t_r16_c2_6;
  assign t_r16_c2_10 = t_r16_c2_7 + t_r16_c2_8;
  assign t_r16_c2_11 = t_r16_c2_9 + t_r16_c2_10;
  assign t_r16_c2_12 = t_r16_c2_11 + p_17_3;
  assign out_16_2 = t_r16_c2_12 >> 4;

  assign t_r16_c3_0 = p_15_3 << 1;
  assign t_r16_c3_1 = p_16_2 << 1;
  assign t_r16_c3_2 = p_16_3 << 2;
  assign t_r16_c3_3 = p_16_4 << 1;
  assign t_r16_c3_4 = p_17_3 << 1;
  assign t_r16_c3_5 = t_r16_c3_0 + p_15_2;
  assign t_r16_c3_6 = t_r16_c3_1 + p_15_4;
  assign t_r16_c3_7 = t_r16_c3_2 + t_r16_c3_3;
  assign t_r16_c3_8 = t_r16_c3_4 + p_17_2;
  assign t_r16_c3_9 = t_r16_c3_5 + t_r16_c3_6;
  assign t_r16_c3_10 = t_r16_c3_7 + t_r16_c3_8;
  assign t_r16_c3_11 = t_r16_c3_9 + t_r16_c3_10;
  assign t_r16_c3_12 = t_r16_c3_11 + p_17_4;
  assign out_16_3 = t_r16_c3_12 >> 4;

  assign t_r16_c4_0 = p_15_4 << 1;
  assign t_r16_c4_1 = p_16_3 << 1;
  assign t_r16_c4_2 = p_16_4 << 2;
  assign t_r16_c4_3 = p_16_5 << 1;
  assign t_r16_c4_4 = p_17_4 << 1;
  assign t_r16_c4_5 = t_r16_c4_0 + p_15_3;
  assign t_r16_c4_6 = t_r16_c4_1 + p_15_5;
  assign t_r16_c4_7 = t_r16_c4_2 + t_r16_c4_3;
  assign t_r16_c4_8 = t_r16_c4_4 + p_17_3;
  assign t_r16_c4_9 = t_r16_c4_5 + t_r16_c4_6;
  assign t_r16_c4_10 = t_r16_c4_7 + t_r16_c4_8;
  assign t_r16_c4_11 = t_r16_c4_9 + t_r16_c4_10;
  assign t_r16_c4_12 = t_r16_c4_11 + p_17_5;
  assign out_16_4 = t_r16_c4_12 >> 4;

  assign t_r16_c5_0 = p_15_5 << 1;
  assign t_r16_c5_1 = p_16_4 << 1;
  assign t_r16_c5_2 = p_16_5 << 2;
  assign t_r16_c5_3 = p_16_6 << 1;
  assign t_r16_c5_4 = p_17_5 << 1;
  assign t_r16_c5_5 = t_r16_c5_0 + p_15_4;
  assign t_r16_c5_6 = t_r16_c5_1 + p_15_6;
  assign t_r16_c5_7 = t_r16_c5_2 + t_r16_c5_3;
  assign t_r16_c5_8 = t_r16_c5_4 + p_17_4;
  assign t_r16_c5_9 = t_r16_c5_5 + t_r16_c5_6;
  assign t_r16_c5_10 = t_r16_c5_7 + t_r16_c5_8;
  assign t_r16_c5_11 = t_r16_c5_9 + t_r16_c5_10;
  assign t_r16_c5_12 = t_r16_c5_11 + p_17_6;
  assign out_16_5 = t_r16_c5_12 >> 4;

  assign t_r16_c6_0 = p_15_6 << 1;
  assign t_r16_c6_1 = p_16_5 << 1;
  assign t_r16_c6_2 = p_16_6 << 2;
  assign t_r16_c6_3 = p_16_7 << 1;
  assign t_r16_c6_4 = p_17_6 << 1;
  assign t_r16_c6_5 = t_r16_c6_0 + p_15_5;
  assign t_r16_c6_6 = t_r16_c6_1 + p_15_7;
  assign t_r16_c6_7 = t_r16_c6_2 + t_r16_c6_3;
  assign t_r16_c6_8 = t_r16_c6_4 + p_17_5;
  assign t_r16_c6_9 = t_r16_c6_5 + t_r16_c6_6;
  assign t_r16_c6_10 = t_r16_c6_7 + t_r16_c6_8;
  assign t_r16_c6_11 = t_r16_c6_9 + t_r16_c6_10;
  assign t_r16_c6_12 = t_r16_c6_11 + p_17_7;
  assign out_16_6 = t_r16_c6_12 >> 4;

  assign t_r16_c7_0 = p_15_7 << 1;
  assign t_r16_c7_1 = p_16_6 << 1;
  assign t_r16_c7_2 = p_16_7 << 2;
  assign t_r16_c7_3 = p_16_8 << 1;
  assign t_r16_c7_4 = p_17_7 << 1;
  assign t_r16_c7_5 = t_r16_c7_0 + p_15_6;
  assign t_r16_c7_6 = t_r16_c7_1 + p_15_8;
  assign t_r16_c7_7 = t_r16_c7_2 + t_r16_c7_3;
  assign t_r16_c7_8 = t_r16_c7_4 + p_17_6;
  assign t_r16_c7_9 = t_r16_c7_5 + t_r16_c7_6;
  assign t_r16_c7_10 = t_r16_c7_7 + t_r16_c7_8;
  assign t_r16_c7_11 = t_r16_c7_9 + t_r16_c7_10;
  assign t_r16_c7_12 = t_r16_c7_11 + p_17_8;
  assign out_16_7 = t_r16_c7_12 >> 4;

  assign t_r16_c8_0 = p_15_8 << 1;
  assign t_r16_c8_1 = p_16_7 << 1;
  assign t_r16_c8_2 = p_16_8 << 2;
  assign t_r16_c8_3 = p_16_9 << 1;
  assign t_r16_c8_4 = p_17_8 << 1;
  assign t_r16_c8_5 = t_r16_c8_0 + p_15_7;
  assign t_r16_c8_6 = t_r16_c8_1 + p_15_9;
  assign t_r16_c8_7 = t_r16_c8_2 + t_r16_c8_3;
  assign t_r16_c8_8 = t_r16_c8_4 + p_17_7;
  assign t_r16_c8_9 = t_r16_c8_5 + t_r16_c8_6;
  assign t_r16_c8_10 = t_r16_c8_7 + t_r16_c8_8;
  assign t_r16_c8_11 = t_r16_c8_9 + t_r16_c8_10;
  assign t_r16_c8_12 = t_r16_c8_11 + p_17_9;
  assign out_16_8 = t_r16_c8_12 >> 4;

  assign t_r16_c9_0 = p_15_9 << 1;
  assign t_r16_c9_1 = p_16_8 << 1;
  assign t_r16_c9_2 = p_16_9 << 2;
  assign t_r16_c9_3 = p_16_10 << 1;
  assign t_r16_c9_4 = p_17_9 << 1;
  assign t_r16_c9_5 = t_r16_c9_0 + p_15_8;
  assign t_r16_c9_6 = t_r16_c9_1 + p_15_10;
  assign t_r16_c9_7 = t_r16_c9_2 + t_r16_c9_3;
  assign t_r16_c9_8 = t_r16_c9_4 + p_17_8;
  assign t_r16_c9_9 = t_r16_c9_5 + t_r16_c9_6;
  assign t_r16_c9_10 = t_r16_c9_7 + t_r16_c9_8;
  assign t_r16_c9_11 = t_r16_c9_9 + t_r16_c9_10;
  assign t_r16_c9_12 = t_r16_c9_11 + p_17_10;
  assign out_16_9 = t_r16_c9_12 >> 4;

  assign t_r16_c10_0 = p_15_10 << 1;
  assign t_r16_c10_1 = p_16_9 << 1;
  assign t_r16_c10_2 = p_16_10 << 2;
  assign t_r16_c10_3 = p_16_11 << 1;
  assign t_r16_c10_4 = p_17_10 << 1;
  assign t_r16_c10_5 = t_r16_c10_0 + p_15_9;
  assign t_r16_c10_6 = t_r16_c10_1 + p_15_11;
  assign t_r16_c10_7 = t_r16_c10_2 + t_r16_c10_3;
  assign t_r16_c10_8 = t_r16_c10_4 + p_17_9;
  assign t_r16_c10_9 = t_r16_c10_5 + t_r16_c10_6;
  assign t_r16_c10_10 = t_r16_c10_7 + t_r16_c10_8;
  assign t_r16_c10_11 = t_r16_c10_9 + t_r16_c10_10;
  assign t_r16_c10_12 = t_r16_c10_11 + p_17_11;
  assign out_16_10 = t_r16_c10_12 >> 4;

  assign t_r16_c11_0 = p_15_11 << 1;
  assign t_r16_c11_1 = p_16_10 << 1;
  assign t_r16_c11_2 = p_16_11 << 2;
  assign t_r16_c11_3 = p_16_12 << 1;
  assign t_r16_c11_4 = p_17_11 << 1;
  assign t_r16_c11_5 = t_r16_c11_0 + p_15_10;
  assign t_r16_c11_6 = t_r16_c11_1 + p_15_12;
  assign t_r16_c11_7 = t_r16_c11_2 + t_r16_c11_3;
  assign t_r16_c11_8 = t_r16_c11_4 + p_17_10;
  assign t_r16_c11_9 = t_r16_c11_5 + t_r16_c11_6;
  assign t_r16_c11_10 = t_r16_c11_7 + t_r16_c11_8;
  assign t_r16_c11_11 = t_r16_c11_9 + t_r16_c11_10;
  assign t_r16_c11_12 = t_r16_c11_11 + p_17_12;
  assign out_16_11 = t_r16_c11_12 >> 4;

  assign t_r16_c12_0 = p_15_12 << 1;
  assign t_r16_c12_1 = p_16_11 << 1;
  assign t_r16_c12_2 = p_16_12 << 2;
  assign t_r16_c12_3 = p_16_13 << 1;
  assign t_r16_c12_4 = p_17_12 << 1;
  assign t_r16_c12_5 = t_r16_c12_0 + p_15_11;
  assign t_r16_c12_6 = t_r16_c12_1 + p_15_13;
  assign t_r16_c12_7 = t_r16_c12_2 + t_r16_c12_3;
  assign t_r16_c12_8 = t_r16_c12_4 + p_17_11;
  assign t_r16_c12_9 = t_r16_c12_5 + t_r16_c12_6;
  assign t_r16_c12_10 = t_r16_c12_7 + t_r16_c12_8;
  assign t_r16_c12_11 = t_r16_c12_9 + t_r16_c12_10;
  assign t_r16_c12_12 = t_r16_c12_11 + p_17_13;
  assign out_16_12 = t_r16_c12_12 >> 4;

  assign t_r16_c13_0 = p_15_13 << 1;
  assign t_r16_c13_1 = p_16_12 << 1;
  assign t_r16_c13_2 = p_16_13 << 2;
  assign t_r16_c13_3 = p_16_14 << 1;
  assign t_r16_c13_4 = p_17_13 << 1;
  assign t_r16_c13_5 = t_r16_c13_0 + p_15_12;
  assign t_r16_c13_6 = t_r16_c13_1 + p_15_14;
  assign t_r16_c13_7 = t_r16_c13_2 + t_r16_c13_3;
  assign t_r16_c13_8 = t_r16_c13_4 + p_17_12;
  assign t_r16_c13_9 = t_r16_c13_5 + t_r16_c13_6;
  assign t_r16_c13_10 = t_r16_c13_7 + t_r16_c13_8;
  assign t_r16_c13_11 = t_r16_c13_9 + t_r16_c13_10;
  assign t_r16_c13_12 = t_r16_c13_11 + p_17_14;
  assign out_16_13 = t_r16_c13_12 >> 4;

  assign t_r16_c14_0 = p_15_14 << 1;
  assign t_r16_c14_1 = p_16_13 << 1;
  assign t_r16_c14_2 = p_16_14 << 2;
  assign t_r16_c14_3 = p_16_15 << 1;
  assign t_r16_c14_4 = p_17_14 << 1;
  assign t_r16_c14_5 = t_r16_c14_0 + p_15_13;
  assign t_r16_c14_6 = t_r16_c14_1 + p_15_15;
  assign t_r16_c14_7 = t_r16_c14_2 + t_r16_c14_3;
  assign t_r16_c14_8 = t_r16_c14_4 + p_17_13;
  assign t_r16_c14_9 = t_r16_c14_5 + t_r16_c14_6;
  assign t_r16_c14_10 = t_r16_c14_7 + t_r16_c14_8;
  assign t_r16_c14_11 = t_r16_c14_9 + t_r16_c14_10;
  assign t_r16_c14_12 = t_r16_c14_11 + p_17_15;
  assign out_16_14 = t_r16_c14_12 >> 4;

  assign t_r16_c15_0 = p_15_15 << 1;
  assign t_r16_c15_1 = p_16_14 << 1;
  assign t_r16_c15_2 = p_16_15 << 2;
  assign t_r16_c15_3 = p_16_16 << 1;
  assign t_r16_c15_4 = p_17_15 << 1;
  assign t_r16_c15_5 = t_r16_c15_0 + p_15_14;
  assign t_r16_c15_6 = t_r16_c15_1 + p_15_16;
  assign t_r16_c15_7 = t_r16_c15_2 + t_r16_c15_3;
  assign t_r16_c15_8 = t_r16_c15_4 + p_17_14;
  assign t_r16_c15_9 = t_r16_c15_5 + t_r16_c15_6;
  assign t_r16_c15_10 = t_r16_c15_7 + t_r16_c15_8;
  assign t_r16_c15_11 = t_r16_c15_9 + t_r16_c15_10;
  assign t_r16_c15_12 = t_r16_c15_11 + p_17_16;
  assign out_16_15 = t_r16_c15_12 >> 4;

  assign t_r16_c16_0 = p_15_16 << 1;
  assign t_r16_c16_1 = p_16_15 << 1;
  assign t_r16_c16_2 = p_16_16 << 2;
  assign t_r16_c16_3 = p_16_17 << 1;
  assign t_r16_c16_4 = p_17_16 << 1;
  assign t_r16_c16_5 = t_r16_c16_0 + p_15_15;
  assign t_r16_c16_6 = t_r16_c16_1 + p_15_17;
  assign t_r16_c16_7 = t_r16_c16_2 + t_r16_c16_3;
  assign t_r16_c16_8 = t_r16_c16_4 + p_17_15;
  assign t_r16_c16_9 = t_r16_c16_5 + t_r16_c16_6;
  assign t_r16_c16_10 = t_r16_c16_7 + t_r16_c16_8;
  assign t_r16_c16_11 = t_r16_c16_9 + t_r16_c16_10;
  assign t_r16_c16_12 = t_r16_c16_11 + p_17_17;
  assign out_16_16 = t_r16_c16_12 >> 4;

  assign t_r16_c17_0 = p_15_17 << 1;
  assign t_r16_c17_1 = p_16_16 << 1;
  assign t_r16_c17_2 = p_16_17 << 2;
  assign t_r16_c17_3 = p_16_18 << 1;
  assign t_r16_c17_4 = p_17_17 << 1;
  assign t_r16_c17_5 = t_r16_c17_0 + p_15_16;
  assign t_r16_c17_6 = t_r16_c17_1 + p_15_18;
  assign t_r16_c17_7 = t_r16_c17_2 + t_r16_c17_3;
  assign t_r16_c17_8 = t_r16_c17_4 + p_17_16;
  assign t_r16_c17_9 = t_r16_c17_5 + t_r16_c17_6;
  assign t_r16_c17_10 = t_r16_c17_7 + t_r16_c17_8;
  assign t_r16_c17_11 = t_r16_c17_9 + t_r16_c17_10;
  assign t_r16_c17_12 = t_r16_c17_11 + p_17_18;
  assign out_16_17 = t_r16_c17_12 >> 4;

  assign t_r16_c18_0 = p_15_18 << 1;
  assign t_r16_c18_1 = p_16_17 << 1;
  assign t_r16_c18_2 = p_16_18 << 2;
  assign t_r16_c18_3 = p_16_19 << 1;
  assign t_r16_c18_4 = p_17_18 << 1;
  assign t_r16_c18_5 = t_r16_c18_0 + p_15_17;
  assign t_r16_c18_6 = t_r16_c18_1 + p_15_19;
  assign t_r16_c18_7 = t_r16_c18_2 + t_r16_c18_3;
  assign t_r16_c18_8 = t_r16_c18_4 + p_17_17;
  assign t_r16_c18_9 = t_r16_c18_5 + t_r16_c18_6;
  assign t_r16_c18_10 = t_r16_c18_7 + t_r16_c18_8;
  assign t_r16_c18_11 = t_r16_c18_9 + t_r16_c18_10;
  assign t_r16_c18_12 = t_r16_c18_11 + p_17_19;
  assign out_16_18 = t_r16_c18_12 >> 4;

  assign t_r16_c19_0 = p_15_19 << 1;
  assign t_r16_c19_1 = p_16_18 << 1;
  assign t_r16_c19_2 = p_16_19 << 2;
  assign t_r16_c19_3 = p_16_20 << 1;
  assign t_r16_c19_4 = p_17_19 << 1;
  assign t_r16_c19_5 = t_r16_c19_0 + p_15_18;
  assign t_r16_c19_6 = t_r16_c19_1 + p_15_20;
  assign t_r16_c19_7 = t_r16_c19_2 + t_r16_c19_3;
  assign t_r16_c19_8 = t_r16_c19_4 + p_17_18;
  assign t_r16_c19_9 = t_r16_c19_5 + t_r16_c19_6;
  assign t_r16_c19_10 = t_r16_c19_7 + t_r16_c19_8;
  assign t_r16_c19_11 = t_r16_c19_9 + t_r16_c19_10;
  assign t_r16_c19_12 = t_r16_c19_11 + p_17_20;
  assign out_16_19 = t_r16_c19_12 >> 4;

  assign t_r16_c20_0 = p_15_20 << 1;
  assign t_r16_c20_1 = p_16_19 << 1;
  assign t_r16_c20_2 = p_16_20 << 2;
  assign t_r16_c20_3 = p_16_21 << 1;
  assign t_r16_c20_4 = p_17_20 << 1;
  assign t_r16_c20_5 = t_r16_c20_0 + p_15_19;
  assign t_r16_c20_6 = t_r16_c20_1 + p_15_21;
  assign t_r16_c20_7 = t_r16_c20_2 + t_r16_c20_3;
  assign t_r16_c20_8 = t_r16_c20_4 + p_17_19;
  assign t_r16_c20_9 = t_r16_c20_5 + t_r16_c20_6;
  assign t_r16_c20_10 = t_r16_c20_7 + t_r16_c20_8;
  assign t_r16_c20_11 = t_r16_c20_9 + t_r16_c20_10;
  assign t_r16_c20_12 = t_r16_c20_11 + p_17_21;
  assign out_16_20 = t_r16_c20_12 >> 4;

  assign t_r16_c21_0 = p_15_21 << 1;
  assign t_r16_c21_1 = p_16_20 << 1;
  assign t_r16_c21_2 = p_16_21 << 2;
  assign t_r16_c21_3 = p_16_22 << 1;
  assign t_r16_c21_4 = p_17_21 << 1;
  assign t_r16_c21_5 = t_r16_c21_0 + p_15_20;
  assign t_r16_c21_6 = t_r16_c21_1 + p_15_22;
  assign t_r16_c21_7 = t_r16_c21_2 + t_r16_c21_3;
  assign t_r16_c21_8 = t_r16_c21_4 + p_17_20;
  assign t_r16_c21_9 = t_r16_c21_5 + t_r16_c21_6;
  assign t_r16_c21_10 = t_r16_c21_7 + t_r16_c21_8;
  assign t_r16_c21_11 = t_r16_c21_9 + t_r16_c21_10;
  assign t_r16_c21_12 = t_r16_c21_11 + p_17_22;
  assign out_16_21 = t_r16_c21_12 >> 4;

  assign t_r16_c22_0 = p_15_22 << 1;
  assign t_r16_c22_1 = p_16_21 << 1;
  assign t_r16_c22_2 = p_16_22 << 2;
  assign t_r16_c22_3 = p_16_23 << 1;
  assign t_r16_c22_4 = p_17_22 << 1;
  assign t_r16_c22_5 = t_r16_c22_0 + p_15_21;
  assign t_r16_c22_6 = t_r16_c22_1 + p_15_23;
  assign t_r16_c22_7 = t_r16_c22_2 + t_r16_c22_3;
  assign t_r16_c22_8 = t_r16_c22_4 + p_17_21;
  assign t_r16_c22_9 = t_r16_c22_5 + t_r16_c22_6;
  assign t_r16_c22_10 = t_r16_c22_7 + t_r16_c22_8;
  assign t_r16_c22_11 = t_r16_c22_9 + t_r16_c22_10;
  assign t_r16_c22_12 = t_r16_c22_11 + p_17_23;
  assign out_16_22 = t_r16_c22_12 >> 4;

  assign t_r16_c23_0 = p_15_23 << 1;
  assign t_r16_c23_1 = p_16_22 << 1;
  assign t_r16_c23_2 = p_16_23 << 2;
  assign t_r16_c23_3 = p_16_24 << 1;
  assign t_r16_c23_4 = p_17_23 << 1;
  assign t_r16_c23_5 = t_r16_c23_0 + p_15_22;
  assign t_r16_c23_6 = t_r16_c23_1 + p_15_24;
  assign t_r16_c23_7 = t_r16_c23_2 + t_r16_c23_3;
  assign t_r16_c23_8 = t_r16_c23_4 + p_17_22;
  assign t_r16_c23_9 = t_r16_c23_5 + t_r16_c23_6;
  assign t_r16_c23_10 = t_r16_c23_7 + t_r16_c23_8;
  assign t_r16_c23_11 = t_r16_c23_9 + t_r16_c23_10;
  assign t_r16_c23_12 = t_r16_c23_11 + p_17_24;
  assign out_16_23 = t_r16_c23_12 >> 4;

  assign t_r16_c24_0 = p_15_24 << 1;
  assign t_r16_c24_1 = p_16_23 << 1;
  assign t_r16_c24_2 = p_16_24 << 2;
  assign t_r16_c24_3 = p_16_25 << 1;
  assign t_r16_c24_4 = p_17_24 << 1;
  assign t_r16_c24_5 = t_r16_c24_0 + p_15_23;
  assign t_r16_c24_6 = t_r16_c24_1 + p_15_25;
  assign t_r16_c24_7 = t_r16_c24_2 + t_r16_c24_3;
  assign t_r16_c24_8 = t_r16_c24_4 + p_17_23;
  assign t_r16_c24_9 = t_r16_c24_5 + t_r16_c24_6;
  assign t_r16_c24_10 = t_r16_c24_7 + t_r16_c24_8;
  assign t_r16_c24_11 = t_r16_c24_9 + t_r16_c24_10;
  assign t_r16_c24_12 = t_r16_c24_11 + p_17_25;
  assign out_16_24 = t_r16_c24_12 >> 4;

  assign t_r16_c25_0 = p_15_25 << 1;
  assign t_r16_c25_1 = p_16_24 << 1;
  assign t_r16_c25_2 = p_16_25 << 2;
  assign t_r16_c25_3 = p_16_26 << 1;
  assign t_r16_c25_4 = p_17_25 << 1;
  assign t_r16_c25_5 = t_r16_c25_0 + p_15_24;
  assign t_r16_c25_6 = t_r16_c25_1 + p_15_26;
  assign t_r16_c25_7 = t_r16_c25_2 + t_r16_c25_3;
  assign t_r16_c25_8 = t_r16_c25_4 + p_17_24;
  assign t_r16_c25_9 = t_r16_c25_5 + t_r16_c25_6;
  assign t_r16_c25_10 = t_r16_c25_7 + t_r16_c25_8;
  assign t_r16_c25_11 = t_r16_c25_9 + t_r16_c25_10;
  assign t_r16_c25_12 = t_r16_c25_11 + p_17_26;
  assign out_16_25 = t_r16_c25_12 >> 4;

  assign t_r16_c26_0 = p_15_26 << 1;
  assign t_r16_c26_1 = p_16_25 << 1;
  assign t_r16_c26_2 = p_16_26 << 2;
  assign t_r16_c26_3 = p_16_27 << 1;
  assign t_r16_c26_4 = p_17_26 << 1;
  assign t_r16_c26_5 = t_r16_c26_0 + p_15_25;
  assign t_r16_c26_6 = t_r16_c26_1 + p_15_27;
  assign t_r16_c26_7 = t_r16_c26_2 + t_r16_c26_3;
  assign t_r16_c26_8 = t_r16_c26_4 + p_17_25;
  assign t_r16_c26_9 = t_r16_c26_5 + t_r16_c26_6;
  assign t_r16_c26_10 = t_r16_c26_7 + t_r16_c26_8;
  assign t_r16_c26_11 = t_r16_c26_9 + t_r16_c26_10;
  assign t_r16_c26_12 = t_r16_c26_11 + p_17_27;
  assign out_16_26 = t_r16_c26_12 >> 4;

  assign t_r16_c27_0 = p_15_27 << 1;
  assign t_r16_c27_1 = p_16_26 << 1;
  assign t_r16_c27_2 = p_16_27 << 2;
  assign t_r16_c27_3 = p_16_28 << 1;
  assign t_r16_c27_4 = p_17_27 << 1;
  assign t_r16_c27_5 = t_r16_c27_0 + p_15_26;
  assign t_r16_c27_6 = t_r16_c27_1 + p_15_28;
  assign t_r16_c27_7 = t_r16_c27_2 + t_r16_c27_3;
  assign t_r16_c27_8 = t_r16_c27_4 + p_17_26;
  assign t_r16_c27_9 = t_r16_c27_5 + t_r16_c27_6;
  assign t_r16_c27_10 = t_r16_c27_7 + t_r16_c27_8;
  assign t_r16_c27_11 = t_r16_c27_9 + t_r16_c27_10;
  assign t_r16_c27_12 = t_r16_c27_11 + p_17_28;
  assign out_16_27 = t_r16_c27_12 >> 4;

  assign t_r16_c28_0 = p_15_28 << 1;
  assign t_r16_c28_1 = p_16_27 << 1;
  assign t_r16_c28_2 = p_16_28 << 2;
  assign t_r16_c28_3 = p_16_29 << 1;
  assign t_r16_c28_4 = p_17_28 << 1;
  assign t_r16_c28_5 = t_r16_c28_0 + p_15_27;
  assign t_r16_c28_6 = t_r16_c28_1 + p_15_29;
  assign t_r16_c28_7 = t_r16_c28_2 + t_r16_c28_3;
  assign t_r16_c28_8 = t_r16_c28_4 + p_17_27;
  assign t_r16_c28_9 = t_r16_c28_5 + t_r16_c28_6;
  assign t_r16_c28_10 = t_r16_c28_7 + t_r16_c28_8;
  assign t_r16_c28_11 = t_r16_c28_9 + t_r16_c28_10;
  assign t_r16_c28_12 = t_r16_c28_11 + p_17_29;
  assign out_16_28 = t_r16_c28_12 >> 4;

  assign t_r16_c29_0 = p_15_29 << 1;
  assign t_r16_c29_1 = p_16_28 << 1;
  assign t_r16_c29_2 = p_16_29 << 2;
  assign t_r16_c29_3 = p_16_30 << 1;
  assign t_r16_c29_4 = p_17_29 << 1;
  assign t_r16_c29_5 = t_r16_c29_0 + p_15_28;
  assign t_r16_c29_6 = t_r16_c29_1 + p_15_30;
  assign t_r16_c29_7 = t_r16_c29_2 + t_r16_c29_3;
  assign t_r16_c29_8 = t_r16_c29_4 + p_17_28;
  assign t_r16_c29_9 = t_r16_c29_5 + t_r16_c29_6;
  assign t_r16_c29_10 = t_r16_c29_7 + t_r16_c29_8;
  assign t_r16_c29_11 = t_r16_c29_9 + t_r16_c29_10;
  assign t_r16_c29_12 = t_r16_c29_11 + p_17_30;
  assign out_16_29 = t_r16_c29_12 >> 4;

  assign t_r16_c30_0 = p_15_30 << 1;
  assign t_r16_c30_1 = p_16_29 << 1;
  assign t_r16_c30_2 = p_16_30 << 2;
  assign t_r16_c30_3 = p_16_31 << 1;
  assign t_r16_c30_4 = p_17_30 << 1;
  assign t_r16_c30_5 = t_r16_c30_0 + p_15_29;
  assign t_r16_c30_6 = t_r16_c30_1 + p_15_31;
  assign t_r16_c30_7 = t_r16_c30_2 + t_r16_c30_3;
  assign t_r16_c30_8 = t_r16_c30_4 + p_17_29;
  assign t_r16_c30_9 = t_r16_c30_5 + t_r16_c30_6;
  assign t_r16_c30_10 = t_r16_c30_7 + t_r16_c30_8;
  assign t_r16_c30_11 = t_r16_c30_9 + t_r16_c30_10;
  assign t_r16_c30_12 = t_r16_c30_11 + p_17_31;
  assign out_16_30 = t_r16_c30_12 >> 4;

  assign t_r16_c31_0 = p_15_31 << 1;
  assign t_r16_c31_1 = p_16_30 << 1;
  assign t_r16_c31_2 = p_16_31 << 2;
  assign t_r16_c31_3 = p_16_32 << 1;
  assign t_r16_c31_4 = p_17_31 << 1;
  assign t_r16_c31_5 = t_r16_c31_0 + p_15_30;
  assign t_r16_c31_6 = t_r16_c31_1 + p_15_32;
  assign t_r16_c31_7 = t_r16_c31_2 + t_r16_c31_3;
  assign t_r16_c31_8 = t_r16_c31_4 + p_17_30;
  assign t_r16_c31_9 = t_r16_c31_5 + t_r16_c31_6;
  assign t_r16_c31_10 = t_r16_c31_7 + t_r16_c31_8;
  assign t_r16_c31_11 = t_r16_c31_9 + t_r16_c31_10;
  assign t_r16_c31_12 = t_r16_c31_11 + p_17_32;
  assign out_16_31 = t_r16_c31_12 >> 4;

  assign t_r16_c32_0 = p_15_32 << 1;
  assign t_r16_c32_1 = p_16_31 << 1;
  assign t_r16_c32_2 = p_16_32 << 2;
  assign t_r16_c32_3 = p_16_33 << 1;
  assign t_r16_c32_4 = p_17_32 << 1;
  assign t_r16_c32_5 = t_r16_c32_0 + p_15_31;
  assign t_r16_c32_6 = t_r16_c32_1 + p_15_33;
  assign t_r16_c32_7 = t_r16_c32_2 + t_r16_c32_3;
  assign t_r16_c32_8 = t_r16_c32_4 + p_17_31;
  assign t_r16_c32_9 = t_r16_c32_5 + t_r16_c32_6;
  assign t_r16_c32_10 = t_r16_c32_7 + t_r16_c32_8;
  assign t_r16_c32_11 = t_r16_c32_9 + t_r16_c32_10;
  assign t_r16_c32_12 = t_r16_c32_11 + p_17_33;
  assign out_16_32 = t_r16_c32_12 >> 4;

  assign t_r16_c33_0 = p_15_33 << 1;
  assign t_r16_c33_1 = p_16_32 << 1;
  assign t_r16_c33_2 = p_16_33 << 2;
  assign t_r16_c33_3 = p_16_34 << 1;
  assign t_r16_c33_4 = p_17_33 << 1;
  assign t_r16_c33_5 = t_r16_c33_0 + p_15_32;
  assign t_r16_c33_6 = t_r16_c33_1 + p_15_34;
  assign t_r16_c33_7 = t_r16_c33_2 + t_r16_c33_3;
  assign t_r16_c33_8 = t_r16_c33_4 + p_17_32;
  assign t_r16_c33_9 = t_r16_c33_5 + t_r16_c33_6;
  assign t_r16_c33_10 = t_r16_c33_7 + t_r16_c33_8;
  assign t_r16_c33_11 = t_r16_c33_9 + t_r16_c33_10;
  assign t_r16_c33_12 = t_r16_c33_11 + p_17_34;
  assign out_16_33 = t_r16_c33_12 >> 4;

  assign t_r16_c34_0 = p_15_34 << 1;
  assign t_r16_c34_1 = p_16_33 << 1;
  assign t_r16_c34_2 = p_16_34 << 2;
  assign t_r16_c34_3 = p_16_35 << 1;
  assign t_r16_c34_4 = p_17_34 << 1;
  assign t_r16_c34_5 = t_r16_c34_0 + p_15_33;
  assign t_r16_c34_6 = t_r16_c34_1 + p_15_35;
  assign t_r16_c34_7 = t_r16_c34_2 + t_r16_c34_3;
  assign t_r16_c34_8 = t_r16_c34_4 + p_17_33;
  assign t_r16_c34_9 = t_r16_c34_5 + t_r16_c34_6;
  assign t_r16_c34_10 = t_r16_c34_7 + t_r16_c34_8;
  assign t_r16_c34_11 = t_r16_c34_9 + t_r16_c34_10;
  assign t_r16_c34_12 = t_r16_c34_11 + p_17_35;
  assign out_16_34 = t_r16_c34_12 >> 4;

  assign t_r16_c35_0 = p_15_35 << 1;
  assign t_r16_c35_1 = p_16_34 << 1;
  assign t_r16_c35_2 = p_16_35 << 2;
  assign t_r16_c35_3 = p_16_36 << 1;
  assign t_r16_c35_4 = p_17_35 << 1;
  assign t_r16_c35_5 = t_r16_c35_0 + p_15_34;
  assign t_r16_c35_6 = t_r16_c35_1 + p_15_36;
  assign t_r16_c35_7 = t_r16_c35_2 + t_r16_c35_3;
  assign t_r16_c35_8 = t_r16_c35_4 + p_17_34;
  assign t_r16_c35_9 = t_r16_c35_5 + t_r16_c35_6;
  assign t_r16_c35_10 = t_r16_c35_7 + t_r16_c35_8;
  assign t_r16_c35_11 = t_r16_c35_9 + t_r16_c35_10;
  assign t_r16_c35_12 = t_r16_c35_11 + p_17_36;
  assign out_16_35 = t_r16_c35_12 >> 4;

  assign t_r16_c36_0 = p_15_36 << 1;
  assign t_r16_c36_1 = p_16_35 << 1;
  assign t_r16_c36_2 = p_16_36 << 2;
  assign t_r16_c36_3 = p_16_37 << 1;
  assign t_r16_c36_4 = p_17_36 << 1;
  assign t_r16_c36_5 = t_r16_c36_0 + p_15_35;
  assign t_r16_c36_6 = t_r16_c36_1 + p_15_37;
  assign t_r16_c36_7 = t_r16_c36_2 + t_r16_c36_3;
  assign t_r16_c36_8 = t_r16_c36_4 + p_17_35;
  assign t_r16_c36_9 = t_r16_c36_5 + t_r16_c36_6;
  assign t_r16_c36_10 = t_r16_c36_7 + t_r16_c36_8;
  assign t_r16_c36_11 = t_r16_c36_9 + t_r16_c36_10;
  assign t_r16_c36_12 = t_r16_c36_11 + p_17_37;
  assign out_16_36 = t_r16_c36_12 >> 4;

  assign t_r16_c37_0 = p_15_37 << 1;
  assign t_r16_c37_1 = p_16_36 << 1;
  assign t_r16_c37_2 = p_16_37 << 2;
  assign t_r16_c37_3 = p_16_38 << 1;
  assign t_r16_c37_4 = p_17_37 << 1;
  assign t_r16_c37_5 = t_r16_c37_0 + p_15_36;
  assign t_r16_c37_6 = t_r16_c37_1 + p_15_38;
  assign t_r16_c37_7 = t_r16_c37_2 + t_r16_c37_3;
  assign t_r16_c37_8 = t_r16_c37_4 + p_17_36;
  assign t_r16_c37_9 = t_r16_c37_5 + t_r16_c37_6;
  assign t_r16_c37_10 = t_r16_c37_7 + t_r16_c37_8;
  assign t_r16_c37_11 = t_r16_c37_9 + t_r16_c37_10;
  assign t_r16_c37_12 = t_r16_c37_11 + p_17_38;
  assign out_16_37 = t_r16_c37_12 >> 4;

  assign t_r16_c38_0 = p_15_38 << 1;
  assign t_r16_c38_1 = p_16_37 << 1;
  assign t_r16_c38_2 = p_16_38 << 2;
  assign t_r16_c38_3 = p_16_39 << 1;
  assign t_r16_c38_4 = p_17_38 << 1;
  assign t_r16_c38_5 = t_r16_c38_0 + p_15_37;
  assign t_r16_c38_6 = t_r16_c38_1 + p_15_39;
  assign t_r16_c38_7 = t_r16_c38_2 + t_r16_c38_3;
  assign t_r16_c38_8 = t_r16_c38_4 + p_17_37;
  assign t_r16_c38_9 = t_r16_c38_5 + t_r16_c38_6;
  assign t_r16_c38_10 = t_r16_c38_7 + t_r16_c38_8;
  assign t_r16_c38_11 = t_r16_c38_9 + t_r16_c38_10;
  assign t_r16_c38_12 = t_r16_c38_11 + p_17_39;
  assign out_16_38 = t_r16_c38_12 >> 4;

  assign t_r16_c39_0 = p_15_39 << 1;
  assign t_r16_c39_1 = p_16_38 << 1;
  assign t_r16_c39_2 = p_16_39 << 2;
  assign t_r16_c39_3 = p_16_40 << 1;
  assign t_r16_c39_4 = p_17_39 << 1;
  assign t_r16_c39_5 = t_r16_c39_0 + p_15_38;
  assign t_r16_c39_6 = t_r16_c39_1 + p_15_40;
  assign t_r16_c39_7 = t_r16_c39_2 + t_r16_c39_3;
  assign t_r16_c39_8 = t_r16_c39_4 + p_17_38;
  assign t_r16_c39_9 = t_r16_c39_5 + t_r16_c39_6;
  assign t_r16_c39_10 = t_r16_c39_7 + t_r16_c39_8;
  assign t_r16_c39_11 = t_r16_c39_9 + t_r16_c39_10;
  assign t_r16_c39_12 = t_r16_c39_11 + p_17_40;
  assign out_16_39 = t_r16_c39_12 >> 4;

  assign t_r16_c40_0 = p_15_40 << 1;
  assign t_r16_c40_1 = p_16_39 << 1;
  assign t_r16_c40_2 = p_16_40 << 2;
  assign t_r16_c40_3 = p_16_41 << 1;
  assign t_r16_c40_4 = p_17_40 << 1;
  assign t_r16_c40_5 = t_r16_c40_0 + p_15_39;
  assign t_r16_c40_6 = t_r16_c40_1 + p_15_41;
  assign t_r16_c40_7 = t_r16_c40_2 + t_r16_c40_3;
  assign t_r16_c40_8 = t_r16_c40_4 + p_17_39;
  assign t_r16_c40_9 = t_r16_c40_5 + t_r16_c40_6;
  assign t_r16_c40_10 = t_r16_c40_7 + t_r16_c40_8;
  assign t_r16_c40_11 = t_r16_c40_9 + t_r16_c40_10;
  assign t_r16_c40_12 = t_r16_c40_11 + p_17_41;
  assign out_16_40 = t_r16_c40_12 >> 4;

  assign t_r16_c41_0 = p_15_41 << 1;
  assign t_r16_c41_1 = p_16_40 << 1;
  assign t_r16_c41_2 = p_16_41 << 2;
  assign t_r16_c41_3 = p_16_42 << 1;
  assign t_r16_c41_4 = p_17_41 << 1;
  assign t_r16_c41_5 = t_r16_c41_0 + p_15_40;
  assign t_r16_c41_6 = t_r16_c41_1 + p_15_42;
  assign t_r16_c41_7 = t_r16_c41_2 + t_r16_c41_3;
  assign t_r16_c41_8 = t_r16_c41_4 + p_17_40;
  assign t_r16_c41_9 = t_r16_c41_5 + t_r16_c41_6;
  assign t_r16_c41_10 = t_r16_c41_7 + t_r16_c41_8;
  assign t_r16_c41_11 = t_r16_c41_9 + t_r16_c41_10;
  assign t_r16_c41_12 = t_r16_c41_11 + p_17_42;
  assign out_16_41 = t_r16_c41_12 >> 4;

  assign t_r16_c42_0 = p_15_42 << 1;
  assign t_r16_c42_1 = p_16_41 << 1;
  assign t_r16_c42_2 = p_16_42 << 2;
  assign t_r16_c42_3 = p_16_43 << 1;
  assign t_r16_c42_4 = p_17_42 << 1;
  assign t_r16_c42_5 = t_r16_c42_0 + p_15_41;
  assign t_r16_c42_6 = t_r16_c42_1 + p_15_43;
  assign t_r16_c42_7 = t_r16_c42_2 + t_r16_c42_3;
  assign t_r16_c42_8 = t_r16_c42_4 + p_17_41;
  assign t_r16_c42_9 = t_r16_c42_5 + t_r16_c42_6;
  assign t_r16_c42_10 = t_r16_c42_7 + t_r16_c42_8;
  assign t_r16_c42_11 = t_r16_c42_9 + t_r16_c42_10;
  assign t_r16_c42_12 = t_r16_c42_11 + p_17_43;
  assign out_16_42 = t_r16_c42_12 >> 4;

  assign t_r16_c43_0 = p_15_43 << 1;
  assign t_r16_c43_1 = p_16_42 << 1;
  assign t_r16_c43_2 = p_16_43 << 2;
  assign t_r16_c43_3 = p_16_44 << 1;
  assign t_r16_c43_4 = p_17_43 << 1;
  assign t_r16_c43_5 = t_r16_c43_0 + p_15_42;
  assign t_r16_c43_6 = t_r16_c43_1 + p_15_44;
  assign t_r16_c43_7 = t_r16_c43_2 + t_r16_c43_3;
  assign t_r16_c43_8 = t_r16_c43_4 + p_17_42;
  assign t_r16_c43_9 = t_r16_c43_5 + t_r16_c43_6;
  assign t_r16_c43_10 = t_r16_c43_7 + t_r16_c43_8;
  assign t_r16_c43_11 = t_r16_c43_9 + t_r16_c43_10;
  assign t_r16_c43_12 = t_r16_c43_11 + p_17_44;
  assign out_16_43 = t_r16_c43_12 >> 4;

  assign t_r16_c44_0 = p_15_44 << 1;
  assign t_r16_c44_1 = p_16_43 << 1;
  assign t_r16_c44_2 = p_16_44 << 2;
  assign t_r16_c44_3 = p_16_45 << 1;
  assign t_r16_c44_4 = p_17_44 << 1;
  assign t_r16_c44_5 = t_r16_c44_0 + p_15_43;
  assign t_r16_c44_6 = t_r16_c44_1 + p_15_45;
  assign t_r16_c44_7 = t_r16_c44_2 + t_r16_c44_3;
  assign t_r16_c44_8 = t_r16_c44_4 + p_17_43;
  assign t_r16_c44_9 = t_r16_c44_5 + t_r16_c44_6;
  assign t_r16_c44_10 = t_r16_c44_7 + t_r16_c44_8;
  assign t_r16_c44_11 = t_r16_c44_9 + t_r16_c44_10;
  assign t_r16_c44_12 = t_r16_c44_11 + p_17_45;
  assign out_16_44 = t_r16_c44_12 >> 4;

  assign t_r16_c45_0 = p_15_45 << 1;
  assign t_r16_c45_1 = p_16_44 << 1;
  assign t_r16_c45_2 = p_16_45 << 2;
  assign t_r16_c45_3 = p_16_46 << 1;
  assign t_r16_c45_4 = p_17_45 << 1;
  assign t_r16_c45_5 = t_r16_c45_0 + p_15_44;
  assign t_r16_c45_6 = t_r16_c45_1 + p_15_46;
  assign t_r16_c45_7 = t_r16_c45_2 + t_r16_c45_3;
  assign t_r16_c45_8 = t_r16_c45_4 + p_17_44;
  assign t_r16_c45_9 = t_r16_c45_5 + t_r16_c45_6;
  assign t_r16_c45_10 = t_r16_c45_7 + t_r16_c45_8;
  assign t_r16_c45_11 = t_r16_c45_9 + t_r16_c45_10;
  assign t_r16_c45_12 = t_r16_c45_11 + p_17_46;
  assign out_16_45 = t_r16_c45_12 >> 4;

  assign t_r16_c46_0 = p_15_46 << 1;
  assign t_r16_c46_1 = p_16_45 << 1;
  assign t_r16_c46_2 = p_16_46 << 2;
  assign t_r16_c46_3 = p_16_47 << 1;
  assign t_r16_c46_4 = p_17_46 << 1;
  assign t_r16_c46_5 = t_r16_c46_0 + p_15_45;
  assign t_r16_c46_6 = t_r16_c46_1 + p_15_47;
  assign t_r16_c46_7 = t_r16_c46_2 + t_r16_c46_3;
  assign t_r16_c46_8 = t_r16_c46_4 + p_17_45;
  assign t_r16_c46_9 = t_r16_c46_5 + t_r16_c46_6;
  assign t_r16_c46_10 = t_r16_c46_7 + t_r16_c46_8;
  assign t_r16_c46_11 = t_r16_c46_9 + t_r16_c46_10;
  assign t_r16_c46_12 = t_r16_c46_11 + p_17_47;
  assign out_16_46 = t_r16_c46_12 >> 4;

  assign t_r16_c47_0 = p_15_47 << 1;
  assign t_r16_c47_1 = p_16_46 << 1;
  assign t_r16_c47_2 = p_16_47 << 2;
  assign t_r16_c47_3 = p_16_48 << 1;
  assign t_r16_c47_4 = p_17_47 << 1;
  assign t_r16_c47_5 = t_r16_c47_0 + p_15_46;
  assign t_r16_c47_6 = t_r16_c47_1 + p_15_48;
  assign t_r16_c47_7 = t_r16_c47_2 + t_r16_c47_3;
  assign t_r16_c47_8 = t_r16_c47_4 + p_17_46;
  assign t_r16_c47_9 = t_r16_c47_5 + t_r16_c47_6;
  assign t_r16_c47_10 = t_r16_c47_7 + t_r16_c47_8;
  assign t_r16_c47_11 = t_r16_c47_9 + t_r16_c47_10;
  assign t_r16_c47_12 = t_r16_c47_11 + p_17_48;
  assign out_16_47 = t_r16_c47_12 >> 4;

  assign t_r16_c48_0 = p_15_48 << 1;
  assign t_r16_c48_1 = p_16_47 << 1;
  assign t_r16_c48_2 = p_16_48 << 2;
  assign t_r16_c48_3 = p_16_49 << 1;
  assign t_r16_c48_4 = p_17_48 << 1;
  assign t_r16_c48_5 = t_r16_c48_0 + p_15_47;
  assign t_r16_c48_6 = t_r16_c48_1 + p_15_49;
  assign t_r16_c48_7 = t_r16_c48_2 + t_r16_c48_3;
  assign t_r16_c48_8 = t_r16_c48_4 + p_17_47;
  assign t_r16_c48_9 = t_r16_c48_5 + t_r16_c48_6;
  assign t_r16_c48_10 = t_r16_c48_7 + t_r16_c48_8;
  assign t_r16_c48_11 = t_r16_c48_9 + t_r16_c48_10;
  assign t_r16_c48_12 = t_r16_c48_11 + p_17_49;
  assign out_16_48 = t_r16_c48_12 >> 4;

  assign t_r16_c49_0 = p_15_49 << 1;
  assign t_r16_c49_1 = p_16_48 << 1;
  assign t_r16_c49_2 = p_16_49 << 2;
  assign t_r16_c49_3 = p_16_50 << 1;
  assign t_r16_c49_4 = p_17_49 << 1;
  assign t_r16_c49_5 = t_r16_c49_0 + p_15_48;
  assign t_r16_c49_6 = t_r16_c49_1 + p_15_50;
  assign t_r16_c49_7 = t_r16_c49_2 + t_r16_c49_3;
  assign t_r16_c49_8 = t_r16_c49_4 + p_17_48;
  assign t_r16_c49_9 = t_r16_c49_5 + t_r16_c49_6;
  assign t_r16_c49_10 = t_r16_c49_7 + t_r16_c49_8;
  assign t_r16_c49_11 = t_r16_c49_9 + t_r16_c49_10;
  assign t_r16_c49_12 = t_r16_c49_11 + p_17_50;
  assign out_16_49 = t_r16_c49_12 >> 4;

  assign t_r16_c50_0 = p_15_50 << 1;
  assign t_r16_c50_1 = p_16_49 << 1;
  assign t_r16_c50_2 = p_16_50 << 2;
  assign t_r16_c50_3 = p_16_51 << 1;
  assign t_r16_c50_4 = p_17_50 << 1;
  assign t_r16_c50_5 = t_r16_c50_0 + p_15_49;
  assign t_r16_c50_6 = t_r16_c50_1 + p_15_51;
  assign t_r16_c50_7 = t_r16_c50_2 + t_r16_c50_3;
  assign t_r16_c50_8 = t_r16_c50_4 + p_17_49;
  assign t_r16_c50_9 = t_r16_c50_5 + t_r16_c50_6;
  assign t_r16_c50_10 = t_r16_c50_7 + t_r16_c50_8;
  assign t_r16_c50_11 = t_r16_c50_9 + t_r16_c50_10;
  assign t_r16_c50_12 = t_r16_c50_11 + p_17_51;
  assign out_16_50 = t_r16_c50_12 >> 4;

  assign t_r16_c51_0 = p_15_51 << 1;
  assign t_r16_c51_1 = p_16_50 << 1;
  assign t_r16_c51_2 = p_16_51 << 2;
  assign t_r16_c51_3 = p_16_52 << 1;
  assign t_r16_c51_4 = p_17_51 << 1;
  assign t_r16_c51_5 = t_r16_c51_0 + p_15_50;
  assign t_r16_c51_6 = t_r16_c51_1 + p_15_52;
  assign t_r16_c51_7 = t_r16_c51_2 + t_r16_c51_3;
  assign t_r16_c51_8 = t_r16_c51_4 + p_17_50;
  assign t_r16_c51_9 = t_r16_c51_5 + t_r16_c51_6;
  assign t_r16_c51_10 = t_r16_c51_7 + t_r16_c51_8;
  assign t_r16_c51_11 = t_r16_c51_9 + t_r16_c51_10;
  assign t_r16_c51_12 = t_r16_c51_11 + p_17_52;
  assign out_16_51 = t_r16_c51_12 >> 4;

  assign t_r16_c52_0 = p_15_52 << 1;
  assign t_r16_c52_1 = p_16_51 << 1;
  assign t_r16_c52_2 = p_16_52 << 2;
  assign t_r16_c52_3 = p_16_53 << 1;
  assign t_r16_c52_4 = p_17_52 << 1;
  assign t_r16_c52_5 = t_r16_c52_0 + p_15_51;
  assign t_r16_c52_6 = t_r16_c52_1 + p_15_53;
  assign t_r16_c52_7 = t_r16_c52_2 + t_r16_c52_3;
  assign t_r16_c52_8 = t_r16_c52_4 + p_17_51;
  assign t_r16_c52_9 = t_r16_c52_5 + t_r16_c52_6;
  assign t_r16_c52_10 = t_r16_c52_7 + t_r16_c52_8;
  assign t_r16_c52_11 = t_r16_c52_9 + t_r16_c52_10;
  assign t_r16_c52_12 = t_r16_c52_11 + p_17_53;
  assign out_16_52 = t_r16_c52_12 >> 4;

  assign t_r16_c53_0 = p_15_53 << 1;
  assign t_r16_c53_1 = p_16_52 << 1;
  assign t_r16_c53_2 = p_16_53 << 2;
  assign t_r16_c53_3 = p_16_54 << 1;
  assign t_r16_c53_4 = p_17_53 << 1;
  assign t_r16_c53_5 = t_r16_c53_0 + p_15_52;
  assign t_r16_c53_6 = t_r16_c53_1 + p_15_54;
  assign t_r16_c53_7 = t_r16_c53_2 + t_r16_c53_3;
  assign t_r16_c53_8 = t_r16_c53_4 + p_17_52;
  assign t_r16_c53_9 = t_r16_c53_5 + t_r16_c53_6;
  assign t_r16_c53_10 = t_r16_c53_7 + t_r16_c53_8;
  assign t_r16_c53_11 = t_r16_c53_9 + t_r16_c53_10;
  assign t_r16_c53_12 = t_r16_c53_11 + p_17_54;
  assign out_16_53 = t_r16_c53_12 >> 4;

  assign t_r16_c54_0 = p_15_54 << 1;
  assign t_r16_c54_1 = p_16_53 << 1;
  assign t_r16_c54_2 = p_16_54 << 2;
  assign t_r16_c54_3 = p_16_55 << 1;
  assign t_r16_c54_4 = p_17_54 << 1;
  assign t_r16_c54_5 = t_r16_c54_0 + p_15_53;
  assign t_r16_c54_6 = t_r16_c54_1 + p_15_55;
  assign t_r16_c54_7 = t_r16_c54_2 + t_r16_c54_3;
  assign t_r16_c54_8 = t_r16_c54_4 + p_17_53;
  assign t_r16_c54_9 = t_r16_c54_5 + t_r16_c54_6;
  assign t_r16_c54_10 = t_r16_c54_7 + t_r16_c54_8;
  assign t_r16_c54_11 = t_r16_c54_9 + t_r16_c54_10;
  assign t_r16_c54_12 = t_r16_c54_11 + p_17_55;
  assign out_16_54 = t_r16_c54_12 >> 4;

  assign t_r16_c55_0 = p_15_55 << 1;
  assign t_r16_c55_1 = p_16_54 << 1;
  assign t_r16_c55_2 = p_16_55 << 2;
  assign t_r16_c55_3 = p_16_56 << 1;
  assign t_r16_c55_4 = p_17_55 << 1;
  assign t_r16_c55_5 = t_r16_c55_0 + p_15_54;
  assign t_r16_c55_6 = t_r16_c55_1 + p_15_56;
  assign t_r16_c55_7 = t_r16_c55_2 + t_r16_c55_3;
  assign t_r16_c55_8 = t_r16_c55_4 + p_17_54;
  assign t_r16_c55_9 = t_r16_c55_5 + t_r16_c55_6;
  assign t_r16_c55_10 = t_r16_c55_7 + t_r16_c55_8;
  assign t_r16_c55_11 = t_r16_c55_9 + t_r16_c55_10;
  assign t_r16_c55_12 = t_r16_c55_11 + p_17_56;
  assign out_16_55 = t_r16_c55_12 >> 4;

  assign t_r16_c56_0 = p_15_56 << 1;
  assign t_r16_c56_1 = p_16_55 << 1;
  assign t_r16_c56_2 = p_16_56 << 2;
  assign t_r16_c56_3 = p_16_57 << 1;
  assign t_r16_c56_4 = p_17_56 << 1;
  assign t_r16_c56_5 = t_r16_c56_0 + p_15_55;
  assign t_r16_c56_6 = t_r16_c56_1 + p_15_57;
  assign t_r16_c56_7 = t_r16_c56_2 + t_r16_c56_3;
  assign t_r16_c56_8 = t_r16_c56_4 + p_17_55;
  assign t_r16_c56_9 = t_r16_c56_5 + t_r16_c56_6;
  assign t_r16_c56_10 = t_r16_c56_7 + t_r16_c56_8;
  assign t_r16_c56_11 = t_r16_c56_9 + t_r16_c56_10;
  assign t_r16_c56_12 = t_r16_c56_11 + p_17_57;
  assign out_16_56 = t_r16_c56_12 >> 4;

  assign t_r16_c57_0 = p_15_57 << 1;
  assign t_r16_c57_1 = p_16_56 << 1;
  assign t_r16_c57_2 = p_16_57 << 2;
  assign t_r16_c57_3 = p_16_58 << 1;
  assign t_r16_c57_4 = p_17_57 << 1;
  assign t_r16_c57_5 = t_r16_c57_0 + p_15_56;
  assign t_r16_c57_6 = t_r16_c57_1 + p_15_58;
  assign t_r16_c57_7 = t_r16_c57_2 + t_r16_c57_3;
  assign t_r16_c57_8 = t_r16_c57_4 + p_17_56;
  assign t_r16_c57_9 = t_r16_c57_5 + t_r16_c57_6;
  assign t_r16_c57_10 = t_r16_c57_7 + t_r16_c57_8;
  assign t_r16_c57_11 = t_r16_c57_9 + t_r16_c57_10;
  assign t_r16_c57_12 = t_r16_c57_11 + p_17_58;
  assign out_16_57 = t_r16_c57_12 >> 4;

  assign t_r16_c58_0 = p_15_58 << 1;
  assign t_r16_c58_1 = p_16_57 << 1;
  assign t_r16_c58_2 = p_16_58 << 2;
  assign t_r16_c58_3 = p_16_59 << 1;
  assign t_r16_c58_4 = p_17_58 << 1;
  assign t_r16_c58_5 = t_r16_c58_0 + p_15_57;
  assign t_r16_c58_6 = t_r16_c58_1 + p_15_59;
  assign t_r16_c58_7 = t_r16_c58_2 + t_r16_c58_3;
  assign t_r16_c58_8 = t_r16_c58_4 + p_17_57;
  assign t_r16_c58_9 = t_r16_c58_5 + t_r16_c58_6;
  assign t_r16_c58_10 = t_r16_c58_7 + t_r16_c58_8;
  assign t_r16_c58_11 = t_r16_c58_9 + t_r16_c58_10;
  assign t_r16_c58_12 = t_r16_c58_11 + p_17_59;
  assign out_16_58 = t_r16_c58_12 >> 4;

  assign t_r16_c59_0 = p_15_59 << 1;
  assign t_r16_c59_1 = p_16_58 << 1;
  assign t_r16_c59_2 = p_16_59 << 2;
  assign t_r16_c59_3 = p_16_60 << 1;
  assign t_r16_c59_4 = p_17_59 << 1;
  assign t_r16_c59_5 = t_r16_c59_0 + p_15_58;
  assign t_r16_c59_6 = t_r16_c59_1 + p_15_60;
  assign t_r16_c59_7 = t_r16_c59_2 + t_r16_c59_3;
  assign t_r16_c59_8 = t_r16_c59_4 + p_17_58;
  assign t_r16_c59_9 = t_r16_c59_5 + t_r16_c59_6;
  assign t_r16_c59_10 = t_r16_c59_7 + t_r16_c59_8;
  assign t_r16_c59_11 = t_r16_c59_9 + t_r16_c59_10;
  assign t_r16_c59_12 = t_r16_c59_11 + p_17_60;
  assign out_16_59 = t_r16_c59_12 >> 4;

  assign t_r16_c60_0 = p_15_60 << 1;
  assign t_r16_c60_1 = p_16_59 << 1;
  assign t_r16_c60_2 = p_16_60 << 2;
  assign t_r16_c60_3 = p_16_61 << 1;
  assign t_r16_c60_4 = p_17_60 << 1;
  assign t_r16_c60_5 = t_r16_c60_0 + p_15_59;
  assign t_r16_c60_6 = t_r16_c60_1 + p_15_61;
  assign t_r16_c60_7 = t_r16_c60_2 + t_r16_c60_3;
  assign t_r16_c60_8 = t_r16_c60_4 + p_17_59;
  assign t_r16_c60_9 = t_r16_c60_5 + t_r16_c60_6;
  assign t_r16_c60_10 = t_r16_c60_7 + t_r16_c60_8;
  assign t_r16_c60_11 = t_r16_c60_9 + t_r16_c60_10;
  assign t_r16_c60_12 = t_r16_c60_11 + p_17_61;
  assign out_16_60 = t_r16_c60_12 >> 4;

  assign t_r16_c61_0 = p_15_61 << 1;
  assign t_r16_c61_1 = p_16_60 << 1;
  assign t_r16_c61_2 = p_16_61 << 2;
  assign t_r16_c61_3 = p_16_62 << 1;
  assign t_r16_c61_4 = p_17_61 << 1;
  assign t_r16_c61_5 = t_r16_c61_0 + p_15_60;
  assign t_r16_c61_6 = t_r16_c61_1 + p_15_62;
  assign t_r16_c61_7 = t_r16_c61_2 + t_r16_c61_3;
  assign t_r16_c61_8 = t_r16_c61_4 + p_17_60;
  assign t_r16_c61_9 = t_r16_c61_5 + t_r16_c61_6;
  assign t_r16_c61_10 = t_r16_c61_7 + t_r16_c61_8;
  assign t_r16_c61_11 = t_r16_c61_9 + t_r16_c61_10;
  assign t_r16_c61_12 = t_r16_c61_11 + p_17_62;
  assign out_16_61 = t_r16_c61_12 >> 4;

  assign t_r16_c62_0 = p_15_62 << 1;
  assign t_r16_c62_1 = p_16_61 << 1;
  assign t_r16_c62_2 = p_16_62 << 2;
  assign t_r16_c62_3 = p_16_63 << 1;
  assign t_r16_c62_4 = p_17_62 << 1;
  assign t_r16_c62_5 = t_r16_c62_0 + p_15_61;
  assign t_r16_c62_6 = t_r16_c62_1 + p_15_63;
  assign t_r16_c62_7 = t_r16_c62_2 + t_r16_c62_3;
  assign t_r16_c62_8 = t_r16_c62_4 + p_17_61;
  assign t_r16_c62_9 = t_r16_c62_5 + t_r16_c62_6;
  assign t_r16_c62_10 = t_r16_c62_7 + t_r16_c62_8;
  assign t_r16_c62_11 = t_r16_c62_9 + t_r16_c62_10;
  assign t_r16_c62_12 = t_r16_c62_11 + p_17_63;
  assign out_16_62 = t_r16_c62_12 >> 4;

  assign t_r16_c63_0 = p_15_63 << 1;
  assign t_r16_c63_1 = p_16_62 << 1;
  assign t_r16_c63_2 = p_16_63 << 2;
  assign t_r16_c63_3 = p_16_64 << 1;
  assign t_r16_c63_4 = p_17_63 << 1;
  assign t_r16_c63_5 = t_r16_c63_0 + p_15_62;
  assign t_r16_c63_6 = t_r16_c63_1 + p_15_64;
  assign t_r16_c63_7 = t_r16_c63_2 + t_r16_c63_3;
  assign t_r16_c63_8 = t_r16_c63_4 + p_17_62;
  assign t_r16_c63_9 = t_r16_c63_5 + t_r16_c63_6;
  assign t_r16_c63_10 = t_r16_c63_7 + t_r16_c63_8;
  assign t_r16_c63_11 = t_r16_c63_9 + t_r16_c63_10;
  assign t_r16_c63_12 = t_r16_c63_11 + p_17_64;
  assign out_16_63 = t_r16_c63_12 >> 4;

  assign t_r16_c64_0 = p_15_64 << 1;
  assign t_r16_c64_1 = p_16_63 << 1;
  assign t_r16_c64_2 = p_16_64 << 2;
  assign t_r16_c64_3 = p_16_65 << 1;
  assign t_r16_c64_4 = p_17_64 << 1;
  assign t_r16_c64_5 = t_r16_c64_0 + p_15_63;
  assign t_r16_c64_6 = t_r16_c64_1 + p_15_65;
  assign t_r16_c64_7 = t_r16_c64_2 + t_r16_c64_3;
  assign t_r16_c64_8 = t_r16_c64_4 + p_17_63;
  assign t_r16_c64_9 = t_r16_c64_5 + t_r16_c64_6;
  assign t_r16_c64_10 = t_r16_c64_7 + t_r16_c64_8;
  assign t_r16_c64_11 = t_r16_c64_9 + t_r16_c64_10;
  assign t_r16_c64_12 = t_r16_c64_11 + p_17_65;
  assign out_16_64 = t_r16_c64_12 >> 4;

  assign t_r17_c1_0 = p_16_1 << 1;
  assign t_r17_c1_1 = p_17_0 << 1;
  assign t_r17_c1_2 = p_17_1 << 2;
  assign t_r17_c1_3 = p_17_2 << 1;
  assign t_r17_c1_4 = p_18_1 << 1;
  assign t_r17_c1_5 = t_r17_c1_0 + p_16_0;
  assign t_r17_c1_6 = t_r17_c1_1 + p_16_2;
  assign t_r17_c1_7 = t_r17_c1_2 + t_r17_c1_3;
  assign t_r17_c1_8 = t_r17_c1_4 + p_18_0;
  assign t_r17_c1_9 = t_r17_c1_5 + t_r17_c1_6;
  assign t_r17_c1_10 = t_r17_c1_7 + t_r17_c1_8;
  assign t_r17_c1_11 = t_r17_c1_9 + t_r17_c1_10;
  assign t_r17_c1_12 = t_r17_c1_11 + p_18_2;
  assign out_17_1 = t_r17_c1_12 >> 4;

  assign t_r17_c2_0 = p_16_2 << 1;
  assign t_r17_c2_1 = p_17_1 << 1;
  assign t_r17_c2_2 = p_17_2 << 2;
  assign t_r17_c2_3 = p_17_3 << 1;
  assign t_r17_c2_4 = p_18_2 << 1;
  assign t_r17_c2_5 = t_r17_c2_0 + p_16_1;
  assign t_r17_c2_6 = t_r17_c2_1 + p_16_3;
  assign t_r17_c2_7 = t_r17_c2_2 + t_r17_c2_3;
  assign t_r17_c2_8 = t_r17_c2_4 + p_18_1;
  assign t_r17_c2_9 = t_r17_c2_5 + t_r17_c2_6;
  assign t_r17_c2_10 = t_r17_c2_7 + t_r17_c2_8;
  assign t_r17_c2_11 = t_r17_c2_9 + t_r17_c2_10;
  assign t_r17_c2_12 = t_r17_c2_11 + p_18_3;
  assign out_17_2 = t_r17_c2_12 >> 4;

  assign t_r17_c3_0 = p_16_3 << 1;
  assign t_r17_c3_1 = p_17_2 << 1;
  assign t_r17_c3_2 = p_17_3 << 2;
  assign t_r17_c3_3 = p_17_4 << 1;
  assign t_r17_c3_4 = p_18_3 << 1;
  assign t_r17_c3_5 = t_r17_c3_0 + p_16_2;
  assign t_r17_c3_6 = t_r17_c3_1 + p_16_4;
  assign t_r17_c3_7 = t_r17_c3_2 + t_r17_c3_3;
  assign t_r17_c3_8 = t_r17_c3_4 + p_18_2;
  assign t_r17_c3_9 = t_r17_c3_5 + t_r17_c3_6;
  assign t_r17_c3_10 = t_r17_c3_7 + t_r17_c3_8;
  assign t_r17_c3_11 = t_r17_c3_9 + t_r17_c3_10;
  assign t_r17_c3_12 = t_r17_c3_11 + p_18_4;
  assign out_17_3 = t_r17_c3_12 >> 4;

  assign t_r17_c4_0 = p_16_4 << 1;
  assign t_r17_c4_1 = p_17_3 << 1;
  assign t_r17_c4_2 = p_17_4 << 2;
  assign t_r17_c4_3 = p_17_5 << 1;
  assign t_r17_c4_4 = p_18_4 << 1;
  assign t_r17_c4_5 = t_r17_c4_0 + p_16_3;
  assign t_r17_c4_6 = t_r17_c4_1 + p_16_5;
  assign t_r17_c4_7 = t_r17_c4_2 + t_r17_c4_3;
  assign t_r17_c4_8 = t_r17_c4_4 + p_18_3;
  assign t_r17_c4_9 = t_r17_c4_5 + t_r17_c4_6;
  assign t_r17_c4_10 = t_r17_c4_7 + t_r17_c4_8;
  assign t_r17_c4_11 = t_r17_c4_9 + t_r17_c4_10;
  assign t_r17_c4_12 = t_r17_c4_11 + p_18_5;
  assign out_17_4 = t_r17_c4_12 >> 4;

  assign t_r17_c5_0 = p_16_5 << 1;
  assign t_r17_c5_1 = p_17_4 << 1;
  assign t_r17_c5_2 = p_17_5 << 2;
  assign t_r17_c5_3 = p_17_6 << 1;
  assign t_r17_c5_4 = p_18_5 << 1;
  assign t_r17_c5_5 = t_r17_c5_0 + p_16_4;
  assign t_r17_c5_6 = t_r17_c5_1 + p_16_6;
  assign t_r17_c5_7 = t_r17_c5_2 + t_r17_c5_3;
  assign t_r17_c5_8 = t_r17_c5_4 + p_18_4;
  assign t_r17_c5_9 = t_r17_c5_5 + t_r17_c5_6;
  assign t_r17_c5_10 = t_r17_c5_7 + t_r17_c5_8;
  assign t_r17_c5_11 = t_r17_c5_9 + t_r17_c5_10;
  assign t_r17_c5_12 = t_r17_c5_11 + p_18_6;
  assign out_17_5 = t_r17_c5_12 >> 4;

  assign t_r17_c6_0 = p_16_6 << 1;
  assign t_r17_c6_1 = p_17_5 << 1;
  assign t_r17_c6_2 = p_17_6 << 2;
  assign t_r17_c6_3 = p_17_7 << 1;
  assign t_r17_c6_4 = p_18_6 << 1;
  assign t_r17_c6_5 = t_r17_c6_0 + p_16_5;
  assign t_r17_c6_6 = t_r17_c6_1 + p_16_7;
  assign t_r17_c6_7 = t_r17_c6_2 + t_r17_c6_3;
  assign t_r17_c6_8 = t_r17_c6_4 + p_18_5;
  assign t_r17_c6_9 = t_r17_c6_5 + t_r17_c6_6;
  assign t_r17_c6_10 = t_r17_c6_7 + t_r17_c6_8;
  assign t_r17_c6_11 = t_r17_c6_9 + t_r17_c6_10;
  assign t_r17_c6_12 = t_r17_c6_11 + p_18_7;
  assign out_17_6 = t_r17_c6_12 >> 4;

  assign t_r17_c7_0 = p_16_7 << 1;
  assign t_r17_c7_1 = p_17_6 << 1;
  assign t_r17_c7_2 = p_17_7 << 2;
  assign t_r17_c7_3 = p_17_8 << 1;
  assign t_r17_c7_4 = p_18_7 << 1;
  assign t_r17_c7_5 = t_r17_c7_0 + p_16_6;
  assign t_r17_c7_6 = t_r17_c7_1 + p_16_8;
  assign t_r17_c7_7 = t_r17_c7_2 + t_r17_c7_3;
  assign t_r17_c7_8 = t_r17_c7_4 + p_18_6;
  assign t_r17_c7_9 = t_r17_c7_5 + t_r17_c7_6;
  assign t_r17_c7_10 = t_r17_c7_7 + t_r17_c7_8;
  assign t_r17_c7_11 = t_r17_c7_9 + t_r17_c7_10;
  assign t_r17_c7_12 = t_r17_c7_11 + p_18_8;
  assign out_17_7 = t_r17_c7_12 >> 4;

  assign t_r17_c8_0 = p_16_8 << 1;
  assign t_r17_c8_1 = p_17_7 << 1;
  assign t_r17_c8_2 = p_17_8 << 2;
  assign t_r17_c8_3 = p_17_9 << 1;
  assign t_r17_c8_4 = p_18_8 << 1;
  assign t_r17_c8_5 = t_r17_c8_0 + p_16_7;
  assign t_r17_c8_6 = t_r17_c8_1 + p_16_9;
  assign t_r17_c8_7 = t_r17_c8_2 + t_r17_c8_3;
  assign t_r17_c8_8 = t_r17_c8_4 + p_18_7;
  assign t_r17_c8_9 = t_r17_c8_5 + t_r17_c8_6;
  assign t_r17_c8_10 = t_r17_c8_7 + t_r17_c8_8;
  assign t_r17_c8_11 = t_r17_c8_9 + t_r17_c8_10;
  assign t_r17_c8_12 = t_r17_c8_11 + p_18_9;
  assign out_17_8 = t_r17_c8_12 >> 4;

  assign t_r17_c9_0 = p_16_9 << 1;
  assign t_r17_c9_1 = p_17_8 << 1;
  assign t_r17_c9_2 = p_17_9 << 2;
  assign t_r17_c9_3 = p_17_10 << 1;
  assign t_r17_c9_4 = p_18_9 << 1;
  assign t_r17_c9_5 = t_r17_c9_0 + p_16_8;
  assign t_r17_c9_6 = t_r17_c9_1 + p_16_10;
  assign t_r17_c9_7 = t_r17_c9_2 + t_r17_c9_3;
  assign t_r17_c9_8 = t_r17_c9_4 + p_18_8;
  assign t_r17_c9_9 = t_r17_c9_5 + t_r17_c9_6;
  assign t_r17_c9_10 = t_r17_c9_7 + t_r17_c9_8;
  assign t_r17_c9_11 = t_r17_c9_9 + t_r17_c9_10;
  assign t_r17_c9_12 = t_r17_c9_11 + p_18_10;
  assign out_17_9 = t_r17_c9_12 >> 4;

  assign t_r17_c10_0 = p_16_10 << 1;
  assign t_r17_c10_1 = p_17_9 << 1;
  assign t_r17_c10_2 = p_17_10 << 2;
  assign t_r17_c10_3 = p_17_11 << 1;
  assign t_r17_c10_4 = p_18_10 << 1;
  assign t_r17_c10_5 = t_r17_c10_0 + p_16_9;
  assign t_r17_c10_6 = t_r17_c10_1 + p_16_11;
  assign t_r17_c10_7 = t_r17_c10_2 + t_r17_c10_3;
  assign t_r17_c10_8 = t_r17_c10_4 + p_18_9;
  assign t_r17_c10_9 = t_r17_c10_5 + t_r17_c10_6;
  assign t_r17_c10_10 = t_r17_c10_7 + t_r17_c10_8;
  assign t_r17_c10_11 = t_r17_c10_9 + t_r17_c10_10;
  assign t_r17_c10_12 = t_r17_c10_11 + p_18_11;
  assign out_17_10 = t_r17_c10_12 >> 4;

  assign t_r17_c11_0 = p_16_11 << 1;
  assign t_r17_c11_1 = p_17_10 << 1;
  assign t_r17_c11_2 = p_17_11 << 2;
  assign t_r17_c11_3 = p_17_12 << 1;
  assign t_r17_c11_4 = p_18_11 << 1;
  assign t_r17_c11_5 = t_r17_c11_0 + p_16_10;
  assign t_r17_c11_6 = t_r17_c11_1 + p_16_12;
  assign t_r17_c11_7 = t_r17_c11_2 + t_r17_c11_3;
  assign t_r17_c11_8 = t_r17_c11_4 + p_18_10;
  assign t_r17_c11_9 = t_r17_c11_5 + t_r17_c11_6;
  assign t_r17_c11_10 = t_r17_c11_7 + t_r17_c11_8;
  assign t_r17_c11_11 = t_r17_c11_9 + t_r17_c11_10;
  assign t_r17_c11_12 = t_r17_c11_11 + p_18_12;
  assign out_17_11 = t_r17_c11_12 >> 4;

  assign t_r17_c12_0 = p_16_12 << 1;
  assign t_r17_c12_1 = p_17_11 << 1;
  assign t_r17_c12_2 = p_17_12 << 2;
  assign t_r17_c12_3 = p_17_13 << 1;
  assign t_r17_c12_4 = p_18_12 << 1;
  assign t_r17_c12_5 = t_r17_c12_0 + p_16_11;
  assign t_r17_c12_6 = t_r17_c12_1 + p_16_13;
  assign t_r17_c12_7 = t_r17_c12_2 + t_r17_c12_3;
  assign t_r17_c12_8 = t_r17_c12_4 + p_18_11;
  assign t_r17_c12_9 = t_r17_c12_5 + t_r17_c12_6;
  assign t_r17_c12_10 = t_r17_c12_7 + t_r17_c12_8;
  assign t_r17_c12_11 = t_r17_c12_9 + t_r17_c12_10;
  assign t_r17_c12_12 = t_r17_c12_11 + p_18_13;
  assign out_17_12 = t_r17_c12_12 >> 4;

  assign t_r17_c13_0 = p_16_13 << 1;
  assign t_r17_c13_1 = p_17_12 << 1;
  assign t_r17_c13_2 = p_17_13 << 2;
  assign t_r17_c13_3 = p_17_14 << 1;
  assign t_r17_c13_4 = p_18_13 << 1;
  assign t_r17_c13_5 = t_r17_c13_0 + p_16_12;
  assign t_r17_c13_6 = t_r17_c13_1 + p_16_14;
  assign t_r17_c13_7 = t_r17_c13_2 + t_r17_c13_3;
  assign t_r17_c13_8 = t_r17_c13_4 + p_18_12;
  assign t_r17_c13_9 = t_r17_c13_5 + t_r17_c13_6;
  assign t_r17_c13_10 = t_r17_c13_7 + t_r17_c13_8;
  assign t_r17_c13_11 = t_r17_c13_9 + t_r17_c13_10;
  assign t_r17_c13_12 = t_r17_c13_11 + p_18_14;
  assign out_17_13 = t_r17_c13_12 >> 4;

  assign t_r17_c14_0 = p_16_14 << 1;
  assign t_r17_c14_1 = p_17_13 << 1;
  assign t_r17_c14_2 = p_17_14 << 2;
  assign t_r17_c14_3 = p_17_15 << 1;
  assign t_r17_c14_4 = p_18_14 << 1;
  assign t_r17_c14_5 = t_r17_c14_0 + p_16_13;
  assign t_r17_c14_6 = t_r17_c14_1 + p_16_15;
  assign t_r17_c14_7 = t_r17_c14_2 + t_r17_c14_3;
  assign t_r17_c14_8 = t_r17_c14_4 + p_18_13;
  assign t_r17_c14_9 = t_r17_c14_5 + t_r17_c14_6;
  assign t_r17_c14_10 = t_r17_c14_7 + t_r17_c14_8;
  assign t_r17_c14_11 = t_r17_c14_9 + t_r17_c14_10;
  assign t_r17_c14_12 = t_r17_c14_11 + p_18_15;
  assign out_17_14 = t_r17_c14_12 >> 4;

  assign t_r17_c15_0 = p_16_15 << 1;
  assign t_r17_c15_1 = p_17_14 << 1;
  assign t_r17_c15_2 = p_17_15 << 2;
  assign t_r17_c15_3 = p_17_16 << 1;
  assign t_r17_c15_4 = p_18_15 << 1;
  assign t_r17_c15_5 = t_r17_c15_0 + p_16_14;
  assign t_r17_c15_6 = t_r17_c15_1 + p_16_16;
  assign t_r17_c15_7 = t_r17_c15_2 + t_r17_c15_3;
  assign t_r17_c15_8 = t_r17_c15_4 + p_18_14;
  assign t_r17_c15_9 = t_r17_c15_5 + t_r17_c15_6;
  assign t_r17_c15_10 = t_r17_c15_7 + t_r17_c15_8;
  assign t_r17_c15_11 = t_r17_c15_9 + t_r17_c15_10;
  assign t_r17_c15_12 = t_r17_c15_11 + p_18_16;
  assign out_17_15 = t_r17_c15_12 >> 4;

  assign t_r17_c16_0 = p_16_16 << 1;
  assign t_r17_c16_1 = p_17_15 << 1;
  assign t_r17_c16_2 = p_17_16 << 2;
  assign t_r17_c16_3 = p_17_17 << 1;
  assign t_r17_c16_4 = p_18_16 << 1;
  assign t_r17_c16_5 = t_r17_c16_0 + p_16_15;
  assign t_r17_c16_6 = t_r17_c16_1 + p_16_17;
  assign t_r17_c16_7 = t_r17_c16_2 + t_r17_c16_3;
  assign t_r17_c16_8 = t_r17_c16_4 + p_18_15;
  assign t_r17_c16_9 = t_r17_c16_5 + t_r17_c16_6;
  assign t_r17_c16_10 = t_r17_c16_7 + t_r17_c16_8;
  assign t_r17_c16_11 = t_r17_c16_9 + t_r17_c16_10;
  assign t_r17_c16_12 = t_r17_c16_11 + p_18_17;
  assign out_17_16 = t_r17_c16_12 >> 4;

  assign t_r17_c17_0 = p_16_17 << 1;
  assign t_r17_c17_1 = p_17_16 << 1;
  assign t_r17_c17_2 = p_17_17 << 2;
  assign t_r17_c17_3 = p_17_18 << 1;
  assign t_r17_c17_4 = p_18_17 << 1;
  assign t_r17_c17_5 = t_r17_c17_0 + p_16_16;
  assign t_r17_c17_6 = t_r17_c17_1 + p_16_18;
  assign t_r17_c17_7 = t_r17_c17_2 + t_r17_c17_3;
  assign t_r17_c17_8 = t_r17_c17_4 + p_18_16;
  assign t_r17_c17_9 = t_r17_c17_5 + t_r17_c17_6;
  assign t_r17_c17_10 = t_r17_c17_7 + t_r17_c17_8;
  assign t_r17_c17_11 = t_r17_c17_9 + t_r17_c17_10;
  assign t_r17_c17_12 = t_r17_c17_11 + p_18_18;
  assign out_17_17 = t_r17_c17_12 >> 4;

  assign t_r17_c18_0 = p_16_18 << 1;
  assign t_r17_c18_1 = p_17_17 << 1;
  assign t_r17_c18_2 = p_17_18 << 2;
  assign t_r17_c18_3 = p_17_19 << 1;
  assign t_r17_c18_4 = p_18_18 << 1;
  assign t_r17_c18_5 = t_r17_c18_0 + p_16_17;
  assign t_r17_c18_6 = t_r17_c18_1 + p_16_19;
  assign t_r17_c18_7 = t_r17_c18_2 + t_r17_c18_3;
  assign t_r17_c18_8 = t_r17_c18_4 + p_18_17;
  assign t_r17_c18_9 = t_r17_c18_5 + t_r17_c18_6;
  assign t_r17_c18_10 = t_r17_c18_7 + t_r17_c18_8;
  assign t_r17_c18_11 = t_r17_c18_9 + t_r17_c18_10;
  assign t_r17_c18_12 = t_r17_c18_11 + p_18_19;
  assign out_17_18 = t_r17_c18_12 >> 4;

  assign t_r17_c19_0 = p_16_19 << 1;
  assign t_r17_c19_1 = p_17_18 << 1;
  assign t_r17_c19_2 = p_17_19 << 2;
  assign t_r17_c19_3 = p_17_20 << 1;
  assign t_r17_c19_4 = p_18_19 << 1;
  assign t_r17_c19_5 = t_r17_c19_0 + p_16_18;
  assign t_r17_c19_6 = t_r17_c19_1 + p_16_20;
  assign t_r17_c19_7 = t_r17_c19_2 + t_r17_c19_3;
  assign t_r17_c19_8 = t_r17_c19_4 + p_18_18;
  assign t_r17_c19_9 = t_r17_c19_5 + t_r17_c19_6;
  assign t_r17_c19_10 = t_r17_c19_7 + t_r17_c19_8;
  assign t_r17_c19_11 = t_r17_c19_9 + t_r17_c19_10;
  assign t_r17_c19_12 = t_r17_c19_11 + p_18_20;
  assign out_17_19 = t_r17_c19_12 >> 4;

  assign t_r17_c20_0 = p_16_20 << 1;
  assign t_r17_c20_1 = p_17_19 << 1;
  assign t_r17_c20_2 = p_17_20 << 2;
  assign t_r17_c20_3 = p_17_21 << 1;
  assign t_r17_c20_4 = p_18_20 << 1;
  assign t_r17_c20_5 = t_r17_c20_0 + p_16_19;
  assign t_r17_c20_6 = t_r17_c20_1 + p_16_21;
  assign t_r17_c20_7 = t_r17_c20_2 + t_r17_c20_3;
  assign t_r17_c20_8 = t_r17_c20_4 + p_18_19;
  assign t_r17_c20_9 = t_r17_c20_5 + t_r17_c20_6;
  assign t_r17_c20_10 = t_r17_c20_7 + t_r17_c20_8;
  assign t_r17_c20_11 = t_r17_c20_9 + t_r17_c20_10;
  assign t_r17_c20_12 = t_r17_c20_11 + p_18_21;
  assign out_17_20 = t_r17_c20_12 >> 4;

  assign t_r17_c21_0 = p_16_21 << 1;
  assign t_r17_c21_1 = p_17_20 << 1;
  assign t_r17_c21_2 = p_17_21 << 2;
  assign t_r17_c21_3 = p_17_22 << 1;
  assign t_r17_c21_4 = p_18_21 << 1;
  assign t_r17_c21_5 = t_r17_c21_0 + p_16_20;
  assign t_r17_c21_6 = t_r17_c21_1 + p_16_22;
  assign t_r17_c21_7 = t_r17_c21_2 + t_r17_c21_3;
  assign t_r17_c21_8 = t_r17_c21_4 + p_18_20;
  assign t_r17_c21_9 = t_r17_c21_5 + t_r17_c21_6;
  assign t_r17_c21_10 = t_r17_c21_7 + t_r17_c21_8;
  assign t_r17_c21_11 = t_r17_c21_9 + t_r17_c21_10;
  assign t_r17_c21_12 = t_r17_c21_11 + p_18_22;
  assign out_17_21 = t_r17_c21_12 >> 4;

  assign t_r17_c22_0 = p_16_22 << 1;
  assign t_r17_c22_1 = p_17_21 << 1;
  assign t_r17_c22_2 = p_17_22 << 2;
  assign t_r17_c22_3 = p_17_23 << 1;
  assign t_r17_c22_4 = p_18_22 << 1;
  assign t_r17_c22_5 = t_r17_c22_0 + p_16_21;
  assign t_r17_c22_6 = t_r17_c22_1 + p_16_23;
  assign t_r17_c22_7 = t_r17_c22_2 + t_r17_c22_3;
  assign t_r17_c22_8 = t_r17_c22_4 + p_18_21;
  assign t_r17_c22_9 = t_r17_c22_5 + t_r17_c22_6;
  assign t_r17_c22_10 = t_r17_c22_7 + t_r17_c22_8;
  assign t_r17_c22_11 = t_r17_c22_9 + t_r17_c22_10;
  assign t_r17_c22_12 = t_r17_c22_11 + p_18_23;
  assign out_17_22 = t_r17_c22_12 >> 4;

  assign t_r17_c23_0 = p_16_23 << 1;
  assign t_r17_c23_1 = p_17_22 << 1;
  assign t_r17_c23_2 = p_17_23 << 2;
  assign t_r17_c23_3 = p_17_24 << 1;
  assign t_r17_c23_4 = p_18_23 << 1;
  assign t_r17_c23_5 = t_r17_c23_0 + p_16_22;
  assign t_r17_c23_6 = t_r17_c23_1 + p_16_24;
  assign t_r17_c23_7 = t_r17_c23_2 + t_r17_c23_3;
  assign t_r17_c23_8 = t_r17_c23_4 + p_18_22;
  assign t_r17_c23_9 = t_r17_c23_5 + t_r17_c23_6;
  assign t_r17_c23_10 = t_r17_c23_7 + t_r17_c23_8;
  assign t_r17_c23_11 = t_r17_c23_9 + t_r17_c23_10;
  assign t_r17_c23_12 = t_r17_c23_11 + p_18_24;
  assign out_17_23 = t_r17_c23_12 >> 4;

  assign t_r17_c24_0 = p_16_24 << 1;
  assign t_r17_c24_1 = p_17_23 << 1;
  assign t_r17_c24_2 = p_17_24 << 2;
  assign t_r17_c24_3 = p_17_25 << 1;
  assign t_r17_c24_4 = p_18_24 << 1;
  assign t_r17_c24_5 = t_r17_c24_0 + p_16_23;
  assign t_r17_c24_6 = t_r17_c24_1 + p_16_25;
  assign t_r17_c24_7 = t_r17_c24_2 + t_r17_c24_3;
  assign t_r17_c24_8 = t_r17_c24_4 + p_18_23;
  assign t_r17_c24_9 = t_r17_c24_5 + t_r17_c24_6;
  assign t_r17_c24_10 = t_r17_c24_7 + t_r17_c24_8;
  assign t_r17_c24_11 = t_r17_c24_9 + t_r17_c24_10;
  assign t_r17_c24_12 = t_r17_c24_11 + p_18_25;
  assign out_17_24 = t_r17_c24_12 >> 4;

  assign t_r17_c25_0 = p_16_25 << 1;
  assign t_r17_c25_1 = p_17_24 << 1;
  assign t_r17_c25_2 = p_17_25 << 2;
  assign t_r17_c25_3 = p_17_26 << 1;
  assign t_r17_c25_4 = p_18_25 << 1;
  assign t_r17_c25_5 = t_r17_c25_0 + p_16_24;
  assign t_r17_c25_6 = t_r17_c25_1 + p_16_26;
  assign t_r17_c25_7 = t_r17_c25_2 + t_r17_c25_3;
  assign t_r17_c25_8 = t_r17_c25_4 + p_18_24;
  assign t_r17_c25_9 = t_r17_c25_5 + t_r17_c25_6;
  assign t_r17_c25_10 = t_r17_c25_7 + t_r17_c25_8;
  assign t_r17_c25_11 = t_r17_c25_9 + t_r17_c25_10;
  assign t_r17_c25_12 = t_r17_c25_11 + p_18_26;
  assign out_17_25 = t_r17_c25_12 >> 4;

  assign t_r17_c26_0 = p_16_26 << 1;
  assign t_r17_c26_1 = p_17_25 << 1;
  assign t_r17_c26_2 = p_17_26 << 2;
  assign t_r17_c26_3 = p_17_27 << 1;
  assign t_r17_c26_4 = p_18_26 << 1;
  assign t_r17_c26_5 = t_r17_c26_0 + p_16_25;
  assign t_r17_c26_6 = t_r17_c26_1 + p_16_27;
  assign t_r17_c26_7 = t_r17_c26_2 + t_r17_c26_3;
  assign t_r17_c26_8 = t_r17_c26_4 + p_18_25;
  assign t_r17_c26_9 = t_r17_c26_5 + t_r17_c26_6;
  assign t_r17_c26_10 = t_r17_c26_7 + t_r17_c26_8;
  assign t_r17_c26_11 = t_r17_c26_9 + t_r17_c26_10;
  assign t_r17_c26_12 = t_r17_c26_11 + p_18_27;
  assign out_17_26 = t_r17_c26_12 >> 4;

  assign t_r17_c27_0 = p_16_27 << 1;
  assign t_r17_c27_1 = p_17_26 << 1;
  assign t_r17_c27_2 = p_17_27 << 2;
  assign t_r17_c27_3 = p_17_28 << 1;
  assign t_r17_c27_4 = p_18_27 << 1;
  assign t_r17_c27_5 = t_r17_c27_0 + p_16_26;
  assign t_r17_c27_6 = t_r17_c27_1 + p_16_28;
  assign t_r17_c27_7 = t_r17_c27_2 + t_r17_c27_3;
  assign t_r17_c27_8 = t_r17_c27_4 + p_18_26;
  assign t_r17_c27_9 = t_r17_c27_5 + t_r17_c27_6;
  assign t_r17_c27_10 = t_r17_c27_7 + t_r17_c27_8;
  assign t_r17_c27_11 = t_r17_c27_9 + t_r17_c27_10;
  assign t_r17_c27_12 = t_r17_c27_11 + p_18_28;
  assign out_17_27 = t_r17_c27_12 >> 4;

  assign t_r17_c28_0 = p_16_28 << 1;
  assign t_r17_c28_1 = p_17_27 << 1;
  assign t_r17_c28_2 = p_17_28 << 2;
  assign t_r17_c28_3 = p_17_29 << 1;
  assign t_r17_c28_4 = p_18_28 << 1;
  assign t_r17_c28_5 = t_r17_c28_0 + p_16_27;
  assign t_r17_c28_6 = t_r17_c28_1 + p_16_29;
  assign t_r17_c28_7 = t_r17_c28_2 + t_r17_c28_3;
  assign t_r17_c28_8 = t_r17_c28_4 + p_18_27;
  assign t_r17_c28_9 = t_r17_c28_5 + t_r17_c28_6;
  assign t_r17_c28_10 = t_r17_c28_7 + t_r17_c28_8;
  assign t_r17_c28_11 = t_r17_c28_9 + t_r17_c28_10;
  assign t_r17_c28_12 = t_r17_c28_11 + p_18_29;
  assign out_17_28 = t_r17_c28_12 >> 4;

  assign t_r17_c29_0 = p_16_29 << 1;
  assign t_r17_c29_1 = p_17_28 << 1;
  assign t_r17_c29_2 = p_17_29 << 2;
  assign t_r17_c29_3 = p_17_30 << 1;
  assign t_r17_c29_4 = p_18_29 << 1;
  assign t_r17_c29_5 = t_r17_c29_0 + p_16_28;
  assign t_r17_c29_6 = t_r17_c29_1 + p_16_30;
  assign t_r17_c29_7 = t_r17_c29_2 + t_r17_c29_3;
  assign t_r17_c29_8 = t_r17_c29_4 + p_18_28;
  assign t_r17_c29_9 = t_r17_c29_5 + t_r17_c29_6;
  assign t_r17_c29_10 = t_r17_c29_7 + t_r17_c29_8;
  assign t_r17_c29_11 = t_r17_c29_9 + t_r17_c29_10;
  assign t_r17_c29_12 = t_r17_c29_11 + p_18_30;
  assign out_17_29 = t_r17_c29_12 >> 4;

  assign t_r17_c30_0 = p_16_30 << 1;
  assign t_r17_c30_1 = p_17_29 << 1;
  assign t_r17_c30_2 = p_17_30 << 2;
  assign t_r17_c30_3 = p_17_31 << 1;
  assign t_r17_c30_4 = p_18_30 << 1;
  assign t_r17_c30_5 = t_r17_c30_0 + p_16_29;
  assign t_r17_c30_6 = t_r17_c30_1 + p_16_31;
  assign t_r17_c30_7 = t_r17_c30_2 + t_r17_c30_3;
  assign t_r17_c30_8 = t_r17_c30_4 + p_18_29;
  assign t_r17_c30_9 = t_r17_c30_5 + t_r17_c30_6;
  assign t_r17_c30_10 = t_r17_c30_7 + t_r17_c30_8;
  assign t_r17_c30_11 = t_r17_c30_9 + t_r17_c30_10;
  assign t_r17_c30_12 = t_r17_c30_11 + p_18_31;
  assign out_17_30 = t_r17_c30_12 >> 4;

  assign t_r17_c31_0 = p_16_31 << 1;
  assign t_r17_c31_1 = p_17_30 << 1;
  assign t_r17_c31_2 = p_17_31 << 2;
  assign t_r17_c31_3 = p_17_32 << 1;
  assign t_r17_c31_4 = p_18_31 << 1;
  assign t_r17_c31_5 = t_r17_c31_0 + p_16_30;
  assign t_r17_c31_6 = t_r17_c31_1 + p_16_32;
  assign t_r17_c31_7 = t_r17_c31_2 + t_r17_c31_3;
  assign t_r17_c31_8 = t_r17_c31_4 + p_18_30;
  assign t_r17_c31_9 = t_r17_c31_5 + t_r17_c31_6;
  assign t_r17_c31_10 = t_r17_c31_7 + t_r17_c31_8;
  assign t_r17_c31_11 = t_r17_c31_9 + t_r17_c31_10;
  assign t_r17_c31_12 = t_r17_c31_11 + p_18_32;
  assign out_17_31 = t_r17_c31_12 >> 4;

  assign t_r17_c32_0 = p_16_32 << 1;
  assign t_r17_c32_1 = p_17_31 << 1;
  assign t_r17_c32_2 = p_17_32 << 2;
  assign t_r17_c32_3 = p_17_33 << 1;
  assign t_r17_c32_4 = p_18_32 << 1;
  assign t_r17_c32_5 = t_r17_c32_0 + p_16_31;
  assign t_r17_c32_6 = t_r17_c32_1 + p_16_33;
  assign t_r17_c32_7 = t_r17_c32_2 + t_r17_c32_3;
  assign t_r17_c32_8 = t_r17_c32_4 + p_18_31;
  assign t_r17_c32_9 = t_r17_c32_5 + t_r17_c32_6;
  assign t_r17_c32_10 = t_r17_c32_7 + t_r17_c32_8;
  assign t_r17_c32_11 = t_r17_c32_9 + t_r17_c32_10;
  assign t_r17_c32_12 = t_r17_c32_11 + p_18_33;
  assign out_17_32 = t_r17_c32_12 >> 4;

  assign t_r17_c33_0 = p_16_33 << 1;
  assign t_r17_c33_1 = p_17_32 << 1;
  assign t_r17_c33_2 = p_17_33 << 2;
  assign t_r17_c33_3 = p_17_34 << 1;
  assign t_r17_c33_4 = p_18_33 << 1;
  assign t_r17_c33_5 = t_r17_c33_0 + p_16_32;
  assign t_r17_c33_6 = t_r17_c33_1 + p_16_34;
  assign t_r17_c33_7 = t_r17_c33_2 + t_r17_c33_3;
  assign t_r17_c33_8 = t_r17_c33_4 + p_18_32;
  assign t_r17_c33_9 = t_r17_c33_5 + t_r17_c33_6;
  assign t_r17_c33_10 = t_r17_c33_7 + t_r17_c33_8;
  assign t_r17_c33_11 = t_r17_c33_9 + t_r17_c33_10;
  assign t_r17_c33_12 = t_r17_c33_11 + p_18_34;
  assign out_17_33 = t_r17_c33_12 >> 4;

  assign t_r17_c34_0 = p_16_34 << 1;
  assign t_r17_c34_1 = p_17_33 << 1;
  assign t_r17_c34_2 = p_17_34 << 2;
  assign t_r17_c34_3 = p_17_35 << 1;
  assign t_r17_c34_4 = p_18_34 << 1;
  assign t_r17_c34_5 = t_r17_c34_0 + p_16_33;
  assign t_r17_c34_6 = t_r17_c34_1 + p_16_35;
  assign t_r17_c34_7 = t_r17_c34_2 + t_r17_c34_3;
  assign t_r17_c34_8 = t_r17_c34_4 + p_18_33;
  assign t_r17_c34_9 = t_r17_c34_5 + t_r17_c34_6;
  assign t_r17_c34_10 = t_r17_c34_7 + t_r17_c34_8;
  assign t_r17_c34_11 = t_r17_c34_9 + t_r17_c34_10;
  assign t_r17_c34_12 = t_r17_c34_11 + p_18_35;
  assign out_17_34 = t_r17_c34_12 >> 4;

  assign t_r17_c35_0 = p_16_35 << 1;
  assign t_r17_c35_1 = p_17_34 << 1;
  assign t_r17_c35_2 = p_17_35 << 2;
  assign t_r17_c35_3 = p_17_36 << 1;
  assign t_r17_c35_4 = p_18_35 << 1;
  assign t_r17_c35_5 = t_r17_c35_0 + p_16_34;
  assign t_r17_c35_6 = t_r17_c35_1 + p_16_36;
  assign t_r17_c35_7 = t_r17_c35_2 + t_r17_c35_3;
  assign t_r17_c35_8 = t_r17_c35_4 + p_18_34;
  assign t_r17_c35_9 = t_r17_c35_5 + t_r17_c35_6;
  assign t_r17_c35_10 = t_r17_c35_7 + t_r17_c35_8;
  assign t_r17_c35_11 = t_r17_c35_9 + t_r17_c35_10;
  assign t_r17_c35_12 = t_r17_c35_11 + p_18_36;
  assign out_17_35 = t_r17_c35_12 >> 4;

  assign t_r17_c36_0 = p_16_36 << 1;
  assign t_r17_c36_1 = p_17_35 << 1;
  assign t_r17_c36_2 = p_17_36 << 2;
  assign t_r17_c36_3 = p_17_37 << 1;
  assign t_r17_c36_4 = p_18_36 << 1;
  assign t_r17_c36_5 = t_r17_c36_0 + p_16_35;
  assign t_r17_c36_6 = t_r17_c36_1 + p_16_37;
  assign t_r17_c36_7 = t_r17_c36_2 + t_r17_c36_3;
  assign t_r17_c36_8 = t_r17_c36_4 + p_18_35;
  assign t_r17_c36_9 = t_r17_c36_5 + t_r17_c36_6;
  assign t_r17_c36_10 = t_r17_c36_7 + t_r17_c36_8;
  assign t_r17_c36_11 = t_r17_c36_9 + t_r17_c36_10;
  assign t_r17_c36_12 = t_r17_c36_11 + p_18_37;
  assign out_17_36 = t_r17_c36_12 >> 4;

  assign t_r17_c37_0 = p_16_37 << 1;
  assign t_r17_c37_1 = p_17_36 << 1;
  assign t_r17_c37_2 = p_17_37 << 2;
  assign t_r17_c37_3 = p_17_38 << 1;
  assign t_r17_c37_4 = p_18_37 << 1;
  assign t_r17_c37_5 = t_r17_c37_0 + p_16_36;
  assign t_r17_c37_6 = t_r17_c37_1 + p_16_38;
  assign t_r17_c37_7 = t_r17_c37_2 + t_r17_c37_3;
  assign t_r17_c37_8 = t_r17_c37_4 + p_18_36;
  assign t_r17_c37_9 = t_r17_c37_5 + t_r17_c37_6;
  assign t_r17_c37_10 = t_r17_c37_7 + t_r17_c37_8;
  assign t_r17_c37_11 = t_r17_c37_9 + t_r17_c37_10;
  assign t_r17_c37_12 = t_r17_c37_11 + p_18_38;
  assign out_17_37 = t_r17_c37_12 >> 4;

  assign t_r17_c38_0 = p_16_38 << 1;
  assign t_r17_c38_1 = p_17_37 << 1;
  assign t_r17_c38_2 = p_17_38 << 2;
  assign t_r17_c38_3 = p_17_39 << 1;
  assign t_r17_c38_4 = p_18_38 << 1;
  assign t_r17_c38_5 = t_r17_c38_0 + p_16_37;
  assign t_r17_c38_6 = t_r17_c38_1 + p_16_39;
  assign t_r17_c38_7 = t_r17_c38_2 + t_r17_c38_3;
  assign t_r17_c38_8 = t_r17_c38_4 + p_18_37;
  assign t_r17_c38_9 = t_r17_c38_5 + t_r17_c38_6;
  assign t_r17_c38_10 = t_r17_c38_7 + t_r17_c38_8;
  assign t_r17_c38_11 = t_r17_c38_9 + t_r17_c38_10;
  assign t_r17_c38_12 = t_r17_c38_11 + p_18_39;
  assign out_17_38 = t_r17_c38_12 >> 4;

  assign t_r17_c39_0 = p_16_39 << 1;
  assign t_r17_c39_1 = p_17_38 << 1;
  assign t_r17_c39_2 = p_17_39 << 2;
  assign t_r17_c39_3 = p_17_40 << 1;
  assign t_r17_c39_4 = p_18_39 << 1;
  assign t_r17_c39_5 = t_r17_c39_0 + p_16_38;
  assign t_r17_c39_6 = t_r17_c39_1 + p_16_40;
  assign t_r17_c39_7 = t_r17_c39_2 + t_r17_c39_3;
  assign t_r17_c39_8 = t_r17_c39_4 + p_18_38;
  assign t_r17_c39_9 = t_r17_c39_5 + t_r17_c39_6;
  assign t_r17_c39_10 = t_r17_c39_7 + t_r17_c39_8;
  assign t_r17_c39_11 = t_r17_c39_9 + t_r17_c39_10;
  assign t_r17_c39_12 = t_r17_c39_11 + p_18_40;
  assign out_17_39 = t_r17_c39_12 >> 4;

  assign t_r17_c40_0 = p_16_40 << 1;
  assign t_r17_c40_1 = p_17_39 << 1;
  assign t_r17_c40_2 = p_17_40 << 2;
  assign t_r17_c40_3 = p_17_41 << 1;
  assign t_r17_c40_4 = p_18_40 << 1;
  assign t_r17_c40_5 = t_r17_c40_0 + p_16_39;
  assign t_r17_c40_6 = t_r17_c40_1 + p_16_41;
  assign t_r17_c40_7 = t_r17_c40_2 + t_r17_c40_3;
  assign t_r17_c40_8 = t_r17_c40_4 + p_18_39;
  assign t_r17_c40_9 = t_r17_c40_5 + t_r17_c40_6;
  assign t_r17_c40_10 = t_r17_c40_7 + t_r17_c40_8;
  assign t_r17_c40_11 = t_r17_c40_9 + t_r17_c40_10;
  assign t_r17_c40_12 = t_r17_c40_11 + p_18_41;
  assign out_17_40 = t_r17_c40_12 >> 4;

  assign t_r17_c41_0 = p_16_41 << 1;
  assign t_r17_c41_1 = p_17_40 << 1;
  assign t_r17_c41_2 = p_17_41 << 2;
  assign t_r17_c41_3 = p_17_42 << 1;
  assign t_r17_c41_4 = p_18_41 << 1;
  assign t_r17_c41_5 = t_r17_c41_0 + p_16_40;
  assign t_r17_c41_6 = t_r17_c41_1 + p_16_42;
  assign t_r17_c41_7 = t_r17_c41_2 + t_r17_c41_3;
  assign t_r17_c41_8 = t_r17_c41_4 + p_18_40;
  assign t_r17_c41_9 = t_r17_c41_5 + t_r17_c41_6;
  assign t_r17_c41_10 = t_r17_c41_7 + t_r17_c41_8;
  assign t_r17_c41_11 = t_r17_c41_9 + t_r17_c41_10;
  assign t_r17_c41_12 = t_r17_c41_11 + p_18_42;
  assign out_17_41 = t_r17_c41_12 >> 4;

  assign t_r17_c42_0 = p_16_42 << 1;
  assign t_r17_c42_1 = p_17_41 << 1;
  assign t_r17_c42_2 = p_17_42 << 2;
  assign t_r17_c42_3 = p_17_43 << 1;
  assign t_r17_c42_4 = p_18_42 << 1;
  assign t_r17_c42_5 = t_r17_c42_0 + p_16_41;
  assign t_r17_c42_6 = t_r17_c42_1 + p_16_43;
  assign t_r17_c42_7 = t_r17_c42_2 + t_r17_c42_3;
  assign t_r17_c42_8 = t_r17_c42_4 + p_18_41;
  assign t_r17_c42_9 = t_r17_c42_5 + t_r17_c42_6;
  assign t_r17_c42_10 = t_r17_c42_7 + t_r17_c42_8;
  assign t_r17_c42_11 = t_r17_c42_9 + t_r17_c42_10;
  assign t_r17_c42_12 = t_r17_c42_11 + p_18_43;
  assign out_17_42 = t_r17_c42_12 >> 4;

  assign t_r17_c43_0 = p_16_43 << 1;
  assign t_r17_c43_1 = p_17_42 << 1;
  assign t_r17_c43_2 = p_17_43 << 2;
  assign t_r17_c43_3 = p_17_44 << 1;
  assign t_r17_c43_4 = p_18_43 << 1;
  assign t_r17_c43_5 = t_r17_c43_0 + p_16_42;
  assign t_r17_c43_6 = t_r17_c43_1 + p_16_44;
  assign t_r17_c43_7 = t_r17_c43_2 + t_r17_c43_3;
  assign t_r17_c43_8 = t_r17_c43_4 + p_18_42;
  assign t_r17_c43_9 = t_r17_c43_5 + t_r17_c43_6;
  assign t_r17_c43_10 = t_r17_c43_7 + t_r17_c43_8;
  assign t_r17_c43_11 = t_r17_c43_9 + t_r17_c43_10;
  assign t_r17_c43_12 = t_r17_c43_11 + p_18_44;
  assign out_17_43 = t_r17_c43_12 >> 4;

  assign t_r17_c44_0 = p_16_44 << 1;
  assign t_r17_c44_1 = p_17_43 << 1;
  assign t_r17_c44_2 = p_17_44 << 2;
  assign t_r17_c44_3 = p_17_45 << 1;
  assign t_r17_c44_4 = p_18_44 << 1;
  assign t_r17_c44_5 = t_r17_c44_0 + p_16_43;
  assign t_r17_c44_6 = t_r17_c44_1 + p_16_45;
  assign t_r17_c44_7 = t_r17_c44_2 + t_r17_c44_3;
  assign t_r17_c44_8 = t_r17_c44_4 + p_18_43;
  assign t_r17_c44_9 = t_r17_c44_5 + t_r17_c44_6;
  assign t_r17_c44_10 = t_r17_c44_7 + t_r17_c44_8;
  assign t_r17_c44_11 = t_r17_c44_9 + t_r17_c44_10;
  assign t_r17_c44_12 = t_r17_c44_11 + p_18_45;
  assign out_17_44 = t_r17_c44_12 >> 4;

  assign t_r17_c45_0 = p_16_45 << 1;
  assign t_r17_c45_1 = p_17_44 << 1;
  assign t_r17_c45_2 = p_17_45 << 2;
  assign t_r17_c45_3 = p_17_46 << 1;
  assign t_r17_c45_4 = p_18_45 << 1;
  assign t_r17_c45_5 = t_r17_c45_0 + p_16_44;
  assign t_r17_c45_6 = t_r17_c45_1 + p_16_46;
  assign t_r17_c45_7 = t_r17_c45_2 + t_r17_c45_3;
  assign t_r17_c45_8 = t_r17_c45_4 + p_18_44;
  assign t_r17_c45_9 = t_r17_c45_5 + t_r17_c45_6;
  assign t_r17_c45_10 = t_r17_c45_7 + t_r17_c45_8;
  assign t_r17_c45_11 = t_r17_c45_9 + t_r17_c45_10;
  assign t_r17_c45_12 = t_r17_c45_11 + p_18_46;
  assign out_17_45 = t_r17_c45_12 >> 4;

  assign t_r17_c46_0 = p_16_46 << 1;
  assign t_r17_c46_1 = p_17_45 << 1;
  assign t_r17_c46_2 = p_17_46 << 2;
  assign t_r17_c46_3 = p_17_47 << 1;
  assign t_r17_c46_4 = p_18_46 << 1;
  assign t_r17_c46_5 = t_r17_c46_0 + p_16_45;
  assign t_r17_c46_6 = t_r17_c46_1 + p_16_47;
  assign t_r17_c46_7 = t_r17_c46_2 + t_r17_c46_3;
  assign t_r17_c46_8 = t_r17_c46_4 + p_18_45;
  assign t_r17_c46_9 = t_r17_c46_5 + t_r17_c46_6;
  assign t_r17_c46_10 = t_r17_c46_7 + t_r17_c46_8;
  assign t_r17_c46_11 = t_r17_c46_9 + t_r17_c46_10;
  assign t_r17_c46_12 = t_r17_c46_11 + p_18_47;
  assign out_17_46 = t_r17_c46_12 >> 4;

  assign t_r17_c47_0 = p_16_47 << 1;
  assign t_r17_c47_1 = p_17_46 << 1;
  assign t_r17_c47_2 = p_17_47 << 2;
  assign t_r17_c47_3 = p_17_48 << 1;
  assign t_r17_c47_4 = p_18_47 << 1;
  assign t_r17_c47_5 = t_r17_c47_0 + p_16_46;
  assign t_r17_c47_6 = t_r17_c47_1 + p_16_48;
  assign t_r17_c47_7 = t_r17_c47_2 + t_r17_c47_3;
  assign t_r17_c47_8 = t_r17_c47_4 + p_18_46;
  assign t_r17_c47_9 = t_r17_c47_5 + t_r17_c47_6;
  assign t_r17_c47_10 = t_r17_c47_7 + t_r17_c47_8;
  assign t_r17_c47_11 = t_r17_c47_9 + t_r17_c47_10;
  assign t_r17_c47_12 = t_r17_c47_11 + p_18_48;
  assign out_17_47 = t_r17_c47_12 >> 4;

  assign t_r17_c48_0 = p_16_48 << 1;
  assign t_r17_c48_1 = p_17_47 << 1;
  assign t_r17_c48_2 = p_17_48 << 2;
  assign t_r17_c48_3 = p_17_49 << 1;
  assign t_r17_c48_4 = p_18_48 << 1;
  assign t_r17_c48_5 = t_r17_c48_0 + p_16_47;
  assign t_r17_c48_6 = t_r17_c48_1 + p_16_49;
  assign t_r17_c48_7 = t_r17_c48_2 + t_r17_c48_3;
  assign t_r17_c48_8 = t_r17_c48_4 + p_18_47;
  assign t_r17_c48_9 = t_r17_c48_5 + t_r17_c48_6;
  assign t_r17_c48_10 = t_r17_c48_7 + t_r17_c48_8;
  assign t_r17_c48_11 = t_r17_c48_9 + t_r17_c48_10;
  assign t_r17_c48_12 = t_r17_c48_11 + p_18_49;
  assign out_17_48 = t_r17_c48_12 >> 4;

  assign t_r17_c49_0 = p_16_49 << 1;
  assign t_r17_c49_1 = p_17_48 << 1;
  assign t_r17_c49_2 = p_17_49 << 2;
  assign t_r17_c49_3 = p_17_50 << 1;
  assign t_r17_c49_4 = p_18_49 << 1;
  assign t_r17_c49_5 = t_r17_c49_0 + p_16_48;
  assign t_r17_c49_6 = t_r17_c49_1 + p_16_50;
  assign t_r17_c49_7 = t_r17_c49_2 + t_r17_c49_3;
  assign t_r17_c49_8 = t_r17_c49_4 + p_18_48;
  assign t_r17_c49_9 = t_r17_c49_5 + t_r17_c49_6;
  assign t_r17_c49_10 = t_r17_c49_7 + t_r17_c49_8;
  assign t_r17_c49_11 = t_r17_c49_9 + t_r17_c49_10;
  assign t_r17_c49_12 = t_r17_c49_11 + p_18_50;
  assign out_17_49 = t_r17_c49_12 >> 4;

  assign t_r17_c50_0 = p_16_50 << 1;
  assign t_r17_c50_1 = p_17_49 << 1;
  assign t_r17_c50_2 = p_17_50 << 2;
  assign t_r17_c50_3 = p_17_51 << 1;
  assign t_r17_c50_4 = p_18_50 << 1;
  assign t_r17_c50_5 = t_r17_c50_0 + p_16_49;
  assign t_r17_c50_6 = t_r17_c50_1 + p_16_51;
  assign t_r17_c50_7 = t_r17_c50_2 + t_r17_c50_3;
  assign t_r17_c50_8 = t_r17_c50_4 + p_18_49;
  assign t_r17_c50_9 = t_r17_c50_5 + t_r17_c50_6;
  assign t_r17_c50_10 = t_r17_c50_7 + t_r17_c50_8;
  assign t_r17_c50_11 = t_r17_c50_9 + t_r17_c50_10;
  assign t_r17_c50_12 = t_r17_c50_11 + p_18_51;
  assign out_17_50 = t_r17_c50_12 >> 4;

  assign t_r17_c51_0 = p_16_51 << 1;
  assign t_r17_c51_1 = p_17_50 << 1;
  assign t_r17_c51_2 = p_17_51 << 2;
  assign t_r17_c51_3 = p_17_52 << 1;
  assign t_r17_c51_4 = p_18_51 << 1;
  assign t_r17_c51_5 = t_r17_c51_0 + p_16_50;
  assign t_r17_c51_6 = t_r17_c51_1 + p_16_52;
  assign t_r17_c51_7 = t_r17_c51_2 + t_r17_c51_3;
  assign t_r17_c51_8 = t_r17_c51_4 + p_18_50;
  assign t_r17_c51_9 = t_r17_c51_5 + t_r17_c51_6;
  assign t_r17_c51_10 = t_r17_c51_7 + t_r17_c51_8;
  assign t_r17_c51_11 = t_r17_c51_9 + t_r17_c51_10;
  assign t_r17_c51_12 = t_r17_c51_11 + p_18_52;
  assign out_17_51 = t_r17_c51_12 >> 4;

  assign t_r17_c52_0 = p_16_52 << 1;
  assign t_r17_c52_1 = p_17_51 << 1;
  assign t_r17_c52_2 = p_17_52 << 2;
  assign t_r17_c52_3 = p_17_53 << 1;
  assign t_r17_c52_4 = p_18_52 << 1;
  assign t_r17_c52_5 = t_r17_c52_0 + p_16_51;
  assign t_r17_c52_6 = t_r17_c52_1 + p_16_53;
  assign t_r17_c52_7 = t_r17_c52_2 + t_r17_c52_3;
  assign t_r17_c52_8 = t_r17_c52_4 + p_18_51;
  assign t_r17_c52_9 = t_r17_c52_5 + t_r17_c52_6;
  assign t_r17_c52_10 = t_r17_c52_7 + t_r17_c52_8;
  assign t_r17_c52_11 = t_r17_c52_9 + t_r17_c52_10;
  assign t_r17_c52_12 = t_r17_c52_11 + p_18_53;
  assign out_17_52 = t_r17_c52_12 >> 4;

  assign t_r17_c53_0 = p_16_53 << 1;
  assign t_r17_c53_1 = p_17_52 << 1;
  assign t_r17_c53_2 = p_17_53 << 2;
  assign t_r17_c53_3 = p_17_54 << 1;
  assign t_r17_c53_4 = p_18_53 << 1;
  assign t_r17_c53_5 = t_r17_c53_0 + p_16_52;
  assign t_r17_c53_6 = t_r17_c53_1 + p_16_54;
  assign t_r17_c53_7 = t_r17_c53_2 + t_r17_c53_3;
  assign t_r17_c53_8 = t_r17_c53_4 + p_18_52;
  assign t_r17_c53_9 = t_r17_c53_5 + t_r17_c53_6;
  assign t_r17_c53_10 = t_r17_c53_7 + t_r17_c53_8;
  assign t_r17_c53_11 = t_r17_c53_9 + t_r17_c53_10;
  assign t_r17_c53_12 = t_r17_c53_11 + p_18_54;
  assign out_17_53 = t_r17_c53_12 >> 4;

  assign t_r17_c54_0 = p_16_54 << 1;
  assign t_r17_c54_1 = p_17_53 << 1;
  assign t_r17_c54_2 = p_17_54 << 2;
  assign t_r17_c54_3 = p_17_55 << 1;
  assign t_r17_c54_4 = p_18_54 << 1;
  assign t_r17_c54_5 = t_r17_c54_0 + p_16_53;
  assign t_r17_c54_6 = t_r17_c54_1 + p_16_55;
  assign t_r17_c54_7 = t_r17_c54_2 + t_r17_c54_3;
  assign t_r17_c54_8 = t_r17_c54_4 + p_18_53;
  assign t_r17_c54_9 = t_r17_c54_5 + t_r17_c54_6;
  assign t_r17_c54_10 = t_r17_c54_7 + t_r17_c54_8;
  assign t_r17_c54_11 = t_r17_c54_9 + t_r17_c54_10;
  assign t_r17_c54_12 = t_r17_c54_11 + p_18_55;
  assign out_17_54 = t_r17_c54_12 >> 4;

  assign t_r17_c55_0 = p_16_55 << 1;
  assign t_r17_c55_1 = p_17_54 << 1;
  assign t_r17_c55_2 = p_17_55 << 2;
  assign t_r17_c55_3 = p_17_56 << 1;
  assign t_r17_c55_4 = p_18_55 << 1;
  assign t_r17_c55_5 = t_r17_c55_0 + p_16_54;
  assign t_r17_c55_6 = t_r17_c55_1 + p_16_56;
  assign t_r17_c55_7 = t_r17_c55_2 + t_r17_c55_3;
  assign t_r17_c55_8 = t_r17_c55_4 + p_18_54;
  assign t_r17_c55_9 = t_r17_c55_5 + t_r17_c55_6;
  assign t_r17_c55_10 = t_r17_c55_7 + t_r17_c55_8;
  assign t_r17_c55_11 = t_r17_c55_9 + t_r17_c55_10;
  assign t_r17_c55_12 = t_r17_c55_11 + p_18_56;
  assign out_17_55 = t_r17_c55_12 >> 4;

  assign t_r17_c56_0 = p_16_56 << 1;
  assign t_r17_c56_1 = p_17_55 << 1;
  assign t_r17_c56_2 = p_17_56 << 2;
  assign t_r17_c56_3 = p_17_57 << 1;
  assign t_r17_c56_4 = p_18_56 << 1;
  assign t_r17_c56_5 = t_r17_c56_0 + p_16_55;
  assign t_r17_c56_6 = t_r17_c56_1 + p_16_57;
  assign t_r17_c56_7 = t_r17_c56_2 + t_r17_c56_3;
  assign t_r17_c56_8 = t_r17_c56_4 + p_18_55;
  assign t_r17_c56_9 = t_r17_c56_5 + t_r17_c56_6;
  assign t_r17_c56_10 = t_r17_c56_7 + t_r17_c56_8;
  assign t_r17_c56_11 = t_r17_c56_9 + t_r17_c56_10;
  assign t_r17_c56_12 = t_r17_c56_11 + p_18_57;
  assign out_17_56 = t_r17_c56_12 >> 4;

  assign t_r17_c57_0 = p_16_57 << 1;
  assign t_r17_c57_1 = p_17_56 << 1;
  assign t_r17_c57_2 = p_17_57 << 2;
  assign t_r17_c57_3 = p_17_58 << 1;
  assign t_r17_c57_4 = p_18_57 << 1;
  assign t_r17_c57_5 = t_r17_c57_0 + p_16_56;
  assign t_r17_c57_6 = t_r17_c57_1 + p_16_58;
  assign t_r17_c57_7 = t_r17_c57_2 + t_r17_c57_3;
  assign t_r17_c57_8 = t_r17_c57_4 + p_18_56;
  assign t_r17_c57_9 = t_r17_c57_5 + t_r17_c57_6;
  assign t_r17_c57_10 = t_r17_c57_7 + t_r17_c57_8;
  assign t_r17_c57_11 = t_r17_c57_9 + t_r17_c57_10;
  assign t_r17_c57_12 = t_r17_c57_11 + p_18_58;
  assign out_17_57 = t_r17_c57_12 >> 4;

  assign t_r17_c58_0 = p_16_58 << 1;
  assign t_r17_c58_1 = p_17_57 << 1;
  assign t_r17_c58_2 = p_17_58 << 2;
  assign t_r17_c58_3 = p_17_59 << 1;
  assign t_r17_c58_4 = p_18_58 << 1;
  assign t_r17_c58_5 = t_r17_c58_0 + p_16_57;
  assign t_r17_c58_6 = t_r17_c58_1 + p_16_59;
  assign t_r17_c58_7 = t_r17_c58_2 + t_r17_c58_3;
  assign t_r17_c58_8 = t_r17_c58_4 + p_18_57;
  assign t_r17_c58_9 = t_r17_c58_5 + t_r17_c58_6;
  assign t_r17_c58_10 = t_r17_c58_7 + t_r17_c58_8;
  assign t_r17_c58_11 = t_r17_c58_9 + t_r17_c58_10;
  assign t_r17_c58_12 = t_r17_c58_11 + p_18_59;
  assign out_17_58 = t_r17_c58_12 >> 4;

  assign t_r17_c59_0 = p_16_59 << 1;
  assign t_r17_c59_1 = p_17_58 << 1;
  assign t_r17_c59_2 = p_17_59 << 2;
  assign t_r17_c59_3 = p_17_60 << 1;
  assign t_r17_c59_4 = p_18_59 << 1;
  assign t_r17_c59_5 = t_r17_c59_0 + p_16_58;
  assign t_r17_c59_6 = t_r17_c59_1 + p_16_60;
  assign t_r17_c59_7 = t_r17_c59_2 + t_r17_c59_3;
  assign t_r17_c59_8 = t_r17_c59_4 + p_18_58;
  assign t_r17_c59_9 = t_r17_c59_5 + t_r17_c59_6;
  assign t_r17_c59_10 = t_r17_c59_7 + t_r17_c59_8;
  assign t_r17_c59_11 = t_r17_c59_9 + t_r17_c59_10;
  assign t_r17_c59_12 = t_r17_c59_11 + p_18_60;
  assign out_17_59 = t_r17_c59_12 >> 4;

  assign t_r17_c60_0 = p_16_60 << 1;
  assign t_r17_c60_1 = p_17_59 << 1;
  assign t_r17_c60_2 = p_17_60 << 2;
  assign t_r17_c60_3 = p_17_61 << 1;
  assign t_r17_c60_4 = p_18_60 << 1;
  assign t_r17_c60_5 = t_r17_c60_0 + p_16_59;
  assign t_r17_c60_6 = t_r17_c60_1 + p_16_61;
  assign t_r17_c60_7 = t_r17_c60_2 + t_r17_c60_3;
  assign t_r17_c60_8 = t_r17_c60_4 + p_18_59;
  assign t_r17_c60_9 = t_r17_c60_5 + t_r17_c60_6;
  assign t_r17_c60_10 = t_r17_c60_7 + t_r17_c60_8;
  assign t_r17_c60_11 = t_r17_c60_9 + t_r17_c60_10;
  assign t_r17_c60_12 = t_r17_c60_11 + p_18_61;
  assign out_17_60 = t_r17_c60_12 >> 4;

  assign t_r17_c61_0 = p_16_61 << 1;
  assign t_r17_c61_1 = p_17_60 << 1;
  assign t_r17_c61_2 = p_17_61 << 2;
  assign t_r17_c61_3 = p_17_62 << 1;
  assign t_r17_c61_4 = p_18_61 << 1;
  assign t_r17_c61_5 = t_r17_c61_0 + p_16_60;
  assign t_r17_c61_6 = t_r17_c61_1 + p_16_62;
  assign t_r17_c61_7 = t_r17_c61_2 + t_r17_c61_3;
  assign t_r17_c61_8 = t_r17_c61_4 + p_18_60;
  assign t_r17_c61_9 = t_r17_c61_5 + t_r17_c61_6;
  assign t_r17_c61_10 = t_r17_c61_7 + t_r17_c61_8;
  assign t_r17_c61_11 = t_r17_c61_9 + t_r17_c61_10;
  assign t_r17_c61_12 = t_r17_c61_11 + p_18_62;
  assign out_17_61 = t_r17_c61_12 >> 4;

  assign t_r17_c62_0 = p_16_62 << 1;
  assign t_r17_c62_1 = p_17_61 << 1;
  assign t_r17_c62_2 = p_17_62 << 2;
  assign t_r17_c62_3 = p_17_63 << 1;
  assign t_r17_c62_4 = p_18_62 << 1;
  assign t_r17_c62_5 = t_r17_c62_0 + p_16_61;
  assign t_r17_c62_6 = t_r17_c62_1 + p_16_63;
  assign t_r17_c62_7 = t_r17_c62_2 + t_r17_c62_3;
  assign t_r17_c62_8 = t_r17_c62_4 + p_18_61;
  assign t_r17_c62_9 = t_r17_c62_5 + t_r17_c62_6;
  assign t_r17_c62_10 = t_r17_c62_7 + t_r17_c62_8;
  assign t_r17_c62_11 = t_r17_c62_9 + t_r17_c62_10;
  assign t_r17_c62_12 = t_r17_c62_11 + p_18_63;
  assign out_17_62 = t_r17_c62_12 >> 4;

  assign t_r17_c63_0 = p_16_63 << 1;
  assign t_r17_c63_1 = p_17_62 << 1;
  assign t_r17_c63_2 = p_17_63 << 2;
  assign t_r17_c63_3 = p_17_64 << 1;
  assign t_r17_c63_4 = p_18_63 << 1;
  assign t_r17_c63_5 = t_r17_c63_0 + p_16_62;
  assign t_r17_c63_6 = t_r17_c63_1 + p_16_64;
  assign t_r17_c63_7 = t_r17_c63_2 + t_r17_c63_3;
  assign t_r17_c63_8 = t_r17_c63_4 + p_18_62;
  assign t_r17_c63_9 = t_r17_c63_5 + t_r17_c63_6;
  assign t_r17_c63_10 = t_r17_c63_7 + t_r17_c63_8;
  assign t_r17_c63_11 = t_r17_c63_9 + t_r17_c63_10;
  assign t_r17_c63_12 = t_r17_c63_11 + p_18_64;
  assign out_17_63 = t_r17_c63_12 >> 4;

  assign t_r17_c64_0 = p_16_64 << 1;
  assign t_r17_c64_1 = p_17_63 << 1;
  assign t_r17_c64_2 = p_17_64 << 2;
  assign t_r17_c64_3 = p_17_65 << 1;
  assign t_r17_c64_4 = p_18_64 << 1;
  assign t_r17_c64_5 = t_r17_c64_0 + p_16_63;
  assign t_r17_c64_6 = t_r17_c64_1 + p_16_65;
  assign t_r17_c64_7 = t_r17_c64_2 + t_r17_c64_3;
  assign t_r17_c64_8 = t_r17_c64_4 + p_18_63;
  assign t_r17_c64_9 = t_r17_c64_5 + t_r17_c64_6;
  assign t_r17_c64_10 = t_r17_c64_7 + t_r17_c64_8;
  assign t_r17_c64_11 = t_r17_c64_9 + t_r17_c64_10;
  assign t_r17_c64_12 = t_r17_c64_11 + p_18_65;
  assign out_17_64 = t_r17_c64_12 >> 4;

  assign t_r18_c1_0 = p_17_1 << 1;
  assign t_r18_c1_1 = p_18_0 << 1;
  assign t_r18_c1_2 = p_18_1 << 2;
  assign t_r18_c1_3 = p_18_2 << 1;
  assign t_r18_c1_4 = p_19_1 << 1;
  assign t_r18_c1_5 = t_r18_c1_0 + p_17_0;
  assign t_r18_c1_6 = t_r18_c1_1 + p_17_2;
  assign t_r18_c1_7 = t_r18_c1_2 + t_r18_c1_3;
  assign t_r18_c1_8 = t_r18_c1_4 + p_19_0;
  assign t_r18_c1_9 = t_r18_c1_5 + t_r18_c1_6;
  assign t_r18_c1_10 = t_r18_c1_7 + t_r18_c1_8;
  assign t_r18_c1_11 = t_r18_c1_9 + t_r18_c1_10;
  assign t_r18_c1_12 = t_r18_c1_11 + p_19_2;
  assign out_18_1 = t_r18_c1_12 >> 4;

  assign t_r18_c2_0 = p_17_2 << 1;
  assign t_r18_c2_1 = p_18_1 << 1;
  assign t_r18_c2_2 = p_18_2 << 2;
  assign t_r18_c2_3 = p_18_3 << 1;
  assign t_r18_c2_4 = p_19_2 << 1;
  assign t_r18_c2_5 = t_r18_c2_0 + p_17_1;
  assign t_r18_c2_6 = t_r18_c2_1 + p_17_3;
  assign t_r18_c2_7 = t_r18_c2_2 + t_r18_c2_3;
  assign t_r18_c2_8 = t_r18_c2_4 + p_19_1;
  assign t_r18_c2_9 = t_r18_c2_5 + t_r18_c2_6;
  assign t_r18_c2_10 = t_r18_c2_7 + t_r18_c2_8;
  assign t_r18_c2_11 = t_r18_c2_9 + t_r18_c2_10;
  assign t_r18_c2_12 = t_r18_c2_11 + p_19_3;
  assign out_18_2 = t_r18_c2_12 >> 4;

  assign t_r18_c3_0 = p_17_3 << 1;
  assign t_r18_c3_1 = p_18_2 << 1;
  assign t_r18_c3_2 = p_18_3 << 2;
  assign t_r18_c3_3 = p_18_4 << 1;
  assign t_r18_c3_4 = p_19_3 << 1;
  assign t_r18_c3_5 = t_r18_c3_0 + p_17_2;
  assign t_r18_c3_6 = t_r18_c3_1 + p_17_4;
  assign t_r18_c3_7 = t_r18_c3_2 + t_r18_c3_3;
  assign t_r18_c3_8 = t_r18_c3_4 + p_19_2;
  assign t_r18_c3_9 = t_r18_c3_5 + t_r18_c3_6;
  assign t_r18_c3_10 = t_r18_c3_7 + t_r18_c3_8;
  assign t_r18_c3_11 = t_r18_c3_9 + t_r18_c3_10;
  assign t_r18_c3_12 = t_r18_c3_11 + p_19_4;
  assign out_18_3 = t_r18_c3_12 >> 4;

  assign t_r18_c4_0 = p_17_4 << 1;
  assign t_r18_c4_1 = p_18_3 << 1;
  assign t_r18_c4_2 = p_18_4 << 2;
  assign t_r18_c4_3 = p_18_5 << 1;
  assign t_r18_c4_4 = p_19_4 << 1;
  assign t_r18_c4_5 = t_r18_c4_0 + p_17_3;
  assign t_r18_c4_6 = t_r18_c4_1 + p_17_5;
  assign t_r18_c4_7 = t_r18_c4_2 + t_r18_c4_3;
  assign t_r18_c4_8 = t_r18_c4_4 + p_19_3;
  assign t_r18_c4_9 = t_r18_c4_5 + t_r18_c4_6;
  assign t_r18_c4_10 = t_r18_c4_7 + t_r18_c4_8;
  assign t_r18_c4_11 = t_r18_c4_9 + t_r18_c4_10;
  assign t_r18_c4_12 = t_r18_c4_11 + p_19_5;
  assign out_18_4 = t_r18_c4_12 >> 4;

  assign t_r18_c5_0 = p_17_5 << 1;
  assign t_r18_c5_1 = p_18_4 << 1;
  assign t_r18_c5_2 = p_18_5 << 2;
  assign t_r18_c5_3 = p_18_6 << 1;
  assign t_r18_c5_4 = p_19_5 << 1;
  assign t_r18_c5_5 = t_r18_c5_0 + p_17_4;
  assign t_r18_c5_6 = t_r18_c5_1 + p_17_6;
  assign t_r18_c5_7 = t_r18_c5_2 + t_r18_c5_3;
  assign t_r18_c5_8 = t_r18_c5_4 + p_19_4;
  assign t_r18_c5_9 = t_r18_c5_5 + t_r18_c5_6;
  assign t_r18_c5_10 = t_r18_c5_7 + t_r18_c5_8;
  assign t_r18_c5_11 = t_r18_c5_9 + t_r18_c5_10;
  assign t_r18_c5_12 = t_r18_c5_11 + p_19_6;
  assign out_18_5 = t_r18_c5_12 >> 4;

  assign t_r18_c6_0 = p_17_6 << 1;
  assign t_r18_c6_1 = p_18_5 << 1;
  assign t_r18_c6_2 = p_18_6 << 2;
  assign t_r18_c6_3 = p_18_7 << 1;
  assign t_r18_c6_4 = p_19_6 << 1;
  assign t_r18_c6_5 = t_r18_c6_0 + p_17_5;
  assign t_r18_c6_6 = t_r18_c6_1 + p_17_7;
  assign t_r18_c6_7 = t_r18_c6_2 + t_r18_c6_3;
  assign t_r18_c6_8 = t_r18_c6_4 + p_19_5;
  assign t_r18_c6_9 = t_r18_c6_5 + t_r18_c6_6;
  assign t_r18_c6_10 = t_r18_c6_7 + t_r18_c6_8;
  assign t_r18_c6_11 = t_r18_c6_9 + t_r18_c6_10;
  assign t_r18_c6_12 = t_r18_c6_11 + p_19_7;
  assign out_18_6 = t_r18_c6_12 >> 4;

  assign t_r18_c7_0 = p_17_7 << 1;
  assign t_r18_c7_1 = p_18_6 << 1;
  assign t_r18_c7_2 = p_18_7 << 2;
  assign t_r18_c7_3 = p_18_8 << 1;
  assign t_r18_c7_4 = p_19_7 << 1;
  assign t_r18_c7_5 = t_r18_c7_0 + p_17_6;
  assign t_r18_c7_6 = t_r18_c7_1 + p_17_8;
  assign t_r18_c7_7 = t_r18_c7_2 + t_r18_c7_3;
  assign t_r18_c7_8 = t_r18_c7_4 + p_19_6;
  assign t_r18_c7_9 = t_r18_c7_5 + t_r18_c7_6;
  assign t_r18_c7_10 = t_r18_c7_7 + t_r18_c7_8;
  assign t_r18_c7_11 = t_r18_c7_9 + t_r18_c7_10;
  assign t_r18_c7_12 = t_r18_c7_11 + p_19_8;
  assign out_18_7 = t_r18_c7_12 >> 4;

  assign t_r18_c8_0 = p_17_8 << 1;
  assign t_r18_c8_1 = p_18_7 << 1;
  assign t_r18_c8_2 = p_18_8 << 2;
  assign t_r18_c8_3 = p_18_9 << 1;
  assign t_r18_c8_4 = p_19_8 << 1;
  assign t_r18_c8_5 = t_r18_c8_0 + p_17_7;
  assign t_r18_c8_6 = t_r18_c8_1 + p_17_9;
  assign t_r18_c8_7 = t_r18_c8_2 + t_r18_c8_3;
  assign t_r18_c8_8 = t_r18_c8_4 + p_19_7;
  assign t_r18_c8_9 = t_r18_c8_5 + t_r18_c8_6;
  assign t_r18_c8_10 = t_r18_c8_7 + t_r18_c8_8;
  assign t_r18_c8_11 = t_r18_c8_9 + t_r18_c8_10;
  assign t_r18_c8_12 = t_r18_c8_11 + p_19_9;
  assign out_18_8 = t_r18_c8_12 >> 4;

  assign t_r18_c9_0 = p_17_9 << 1;
  assign t_r18_c9_1 = p_18_8 << 1;
  assign t_r18_c9_2 = p_18_9 << 2;
  assign t_r18_c9_3 = p_18_10 << 1;
  assign t_r18_c9_4 = p_19_9 << 1;
  assign t_r18_c9_5 = t_r18_c9_0 + p_17_8;
  assign t_r18_c9_6 = t_r18_c9_1 + p_17_10;
  assign t_r18_c9_7 = t_r18_c9_2 + t_r18_c9_3;
  assign t_r18_c9_8 = t_r18_c9_4 + p_19_8;
  assign t_r18_c9_9 = t_r18_c9_5 + t_r18_c9_6;
  assign t_r18_c9_10 = t_r18_c9_7 + t_r18_c9_8;
  assign t_r18_c9_11 = t_r18_c9_9 + t_r18_c9_10;
  assign t_r18_c9_12 = t_r18_c9_11 + p_19_10;
  assign out_18_9 = t_r18_c9_12 >> 4;

  assign t_r18_c10_0 = p_17_10 << 1;
  assign t_r18_c10_1 = p_18_9 << 1;
  assign t_r18_c10_2 = p_18_10 << 2;
  assign t_r18_c10_3 = p_18_11 << 1;
  assign t_r18_c10_4 = p_19_10 << 1;
  assign t_r18_c10_5 = t_r18_c10_0 + p_17_9;
  assign t_r18_c10_6 = t_r18_c10_1 + p_17_11;
  assign t_r18_c10_7 = t_r18_c10_2 + t_r18_c10_3;
  assign t_r18_c10_8 = t_r18_c10_4 + p_19_9;
  assign t_r18_c10_9 = t_r18_c10_5 + t_r18_c10_6;
  assign t_r18_c10_10 = t_r18_c10_7 + t_r18_c10_8;
  assign t_r18_c10_11 = t_r18_c10_9 + t_r18_c10_10;
  assign t_r18_c10_12 = t_r18_c10_11 + p_19_11;
  assign out_18_10 = t_r18_c10_12 >> 4;

  assign t_r18_c11_0 = p_17_11 << 1;
  assign t_r18_c11_1 = p_18_10 << 1;
  assign t_r18_c11_2 = p_18_11 << 2;
  assign t_r18_c11_3 = p_18_12 << 1;
  assign t_r18_c11_4 = p_19_11 << 1;
  assign t_r18_c11_5 = t_r18_c11_0 + p_17_10;
  assign t_r18_c11_6 = t_r18_c11_1 + p_17_12;
  assign t_r18_c11_7 = t_r18_c11_2 + t_r18_c11_3;
  assign t_r18_c11_8 = t_r18_c11_4 + p_19_10;
  assign t_r18_c11_9 = t_r18_c11_5 + t_r18_c11_6;
  assign t_r18_c11_10 = t_r18_c11_7 + t_r18_c11_8;
  assign t_r18_c11_11 = t_r18_c11_9 + t_r18_c11_10;
  assign t_r18_c11_12 = t_r18_c11_11 + p_19_12;
  assign out_18_11 = t_r18_c11_12 >> 4;

  assign t_r18_c12_0 = p_17_12 << 1;
  assign t_r18_c12_1 = p_18_11 << 1;
  assign t_r18_c12_2 = p_18_12 << 2;
  assign t_r18_c12_3 = p_18_13 << 1;
  assign t_r18_c12_4 = p_19_12 << 1;
  assign t_r18_c12_5 = t_r18_c12_0 + p_17_11;
  assign t_r18_c12_6 = t_r18_c12_1 + p_17_13;
  assign t_r18_c12_7 = t_r18_c12_2 + t_r18_c12_3;
  assign t_r18_c12_8 = t_r18_c12_4 + p_19_11;
  assign t_r18_c12_9 = t_r18_c12_5 + t_r18_c12_6;
  assign t_r18_c12_10 = t_r18_c12_7 + t_r18_c12_8;
  assign t_r18_c12_11 = t_r18_c12_9 + t_r18_c12_10;
  assign t_r18_c12_12 = t_r18_c12_11 + p_19_13;
  assign out_18_12 = t_r18_c12_12 >> 4;

  assign t_r18_c13_0 = p_17_13 << 1;
  assign t_r18_c13_1 = p_18_12 << 1;
  assign t_r18_c13_2 = p_18_13 << 2;
  assign t_r18_c13_3 = p_18_14 << 1;
  assign t_r18_c13_4 = p_19_13 << 1;
  assign t_r18_c13_5 = t_r18_c13_0 + p_17_12;
  assign t_r18_c13_6 = t_r18_c13_1 + p_17_14;
  assign t_r18_c13_7 = t_r18_c13_2 + t_r18_c13_3;
  assign t_r18_c13_8 = t_r18_c13_4 + p_19_12;
  assign t_r18_c13_9 = t_r18_c13_5 + t_r18_c13_6;
  assign t_r18_c13_10 = t_r18_c13_7 + t_r18_c13_8;
  assign t_r18_c13_11 = t_r18_c13_9 + t_r18_c13_10;
  assign t_r18_c13_12 = t_r18_c13_11 + p_19_14;
  assign out_18_13 = t_r18_c13_12 >> 4;

  assign t_r18_c14_0 = p_17_14 << 1;
  assign t_r18_c14_1 = p_18_13 << 1;
  assign t_r18_c14_2 = p_18_14 << 2;
  assign t_r18_c14_3 = p_18_15 << 1;
  assign t_r18_c14_4 = p_19_14 << 1;
  assign t_r18_c14_5 = t_r18_c14_0 + p_17_13;
  assign t_r18_c14_6 = t_r18_c14_1 + p_17_15;
  assign t_r18_c14_7 = t_r18_c14_2 + t_r18_c14_3;
  assign t_r18_c14_8 = t_r18_c14_4 + p_19_13;
  assign t_r18_c14_9 = t_r18_c14_5 + t_r18_c14_6;
  assign t_r18_c14_10 = t_r18_c14_7 + t_r18_c14_8;
  assign t_r18_c14_11 = t_r18_c14_9 + t_r18_c14_10;
  assign t_r18_c14_12 = t_r18_c14_11 + p_19_15;
  assign out_18_14 = t_r18_c14_12 >> 4;

  assign t_r18_c15_0 = p_17_15 << 1;
  assign t_r18_c15_1 = p_18_14 << 1;
  assign t_r18_c15_2 = p_18_15 << 2;
  assign t_r18_c15_3 = p_18_16 << 1;
  assign t_r18_c15_4 = p_19_15 << 1;
  assign t_r18_c15_5 = t_r18_c15_0 + p_17_14;
  assign t_r18_c15_6 = t_r18_c15_1 + p_17_16;
  assign t_r18_c15_7 = t_r18_c15_2 + t_r18_c15_3;
  assign t_r18_c15_8 = t_r18_c15_4 + p_19_14;
  assign t_r18_c15_9 = t_r18_c15_5 + t_r18_c15_6;
  assign t_r18_c15_10 = t_r18_c15_7 + t_r18_c15_8;
  assign t_r18_c15_11 = t_r18_c15_9 + t_r18_c15_10;
  assign t_r18_c15_12 = t_r18_c15_11 + p_19_16;
  assign out_18_15 = t_r18_c15_12 >> 4;

  assign t_r18_c16_0 = p_17_16 << 1;
  assign t_r18_c16_1 = p_18_15 << 1;
  assign t_r18_c16_2 = p_18_16 << 2;
  assign t_r18_c16_3 = p_18_17 << 1;
  assign t_r18_c16_4 = p_19_16 << 1;
  assign t_r18_c16_5 = t_r18_c16_0 + p_17_15;
  assign t_r18_c16_6 = t_r18_c16_1 + p_17_17;
  assign t_r18_c16_7 = t_r18_c16_2 + t_r18_c16_3;
  assign t_r18_c16_8 = t_r18_c16_4 + p_19_15;
  assign t_r18_c16_9 = t_r18_c16_5 + t_r18_c16_6;
  assign t_r18_c16_10 = t_r18_c16_7 + t_r18_c16_8;
  assign t_r18_c16_11 = t_r18_c16_9 + t_r18_c16_10;
  assign t_r18_c16_12 = t_r18_c16_11 + p_19_17;
  assign out_18_16 = t_r18_c16_12 >> 4;

  assign t_r18_c17_0 = p_17_17 << 1;
  assign t_r18_c17_1 = p_18_16 << 1;
  assign t_r18_c17_2 = p_18_17 << 2;
  assign t_r18_c17_3 = p_18_18 << 1;
  assign t_r18_c17_4 = p_19_17 << 1;
  assign t_r18_c17_5 = t_r18_c17_0 + p_17_16;
  assign t_r18_c17_6 = t_r18_c17_1 + p_17_18;
  assign t_r18_c17_7 = t_r18_c17_2 + t_r18_c17_3;
  assign t_r18_c17_8 = t_r18_c17_4 + p_19_16;
  assign t_r18_c17_9 = t_r18_c17_5 + t_r18_c17_6;
  assign t_r18_c17_10 = t_r18_c17_7 + t_r18_c17_8;
  assign t_r18_c17_11 = t_r18_c17_9 + t_r18_c17_10;
  assign t_r18_c17_12 = t_r18_c17_11 + p_19_18;
  assign out_18_17 = t_r18_c17_12 >> 4;

  assign t_r18_c18_0 = p_17_18 << 1;
  assign t_r18_c18_1 = p_18_17 << 1;
  assign t_r18_c18_2 = p_18_18 << 2;
  assign t_r18_c18_3 = p_18_19 << 1;
  assign t_r18_c18_4 = p_19_18 << 1;
  assign t_r18_c18_5 = t_r18_c18_0 + p_17_17;
  assign t_r18_c18_6 = t_r18_c18_1 + p_17_19;
  assign t_r18_c18_7 = t_r18_c18_2 + t_r18_c18_3;
  assign t_r18_c18_8 = t_r18_c18_4 + p_19_17;
  assign t_r18_c18_9 = t_r18_c18_5 + t_r18_c18_6;
  assign t_r18_c18_10 = t_r18_c18_7 + t_r18_c18_8;
  assign t_r18_c18_11 = t_r18_c18_9 + t_r18_c18_10;
  assign t_r18_c18_12 = t_r18_c18_11 + p_19_19;
  assign out_18_18 = t_r18_c18_12 >> 4;

  assign t_r18_c19_0 = p_17_19 << 1;
  assign t_r18_c19_1 = p_18_18 << 1;
  assign t_r18_c19_2 = p_18_19 << 2;
  assign t_r18_c19_3 = p_18_20 << 1;
  assign t_r18_c19_4 = p_19_19 << 1;
  assign t_r18_c19_5 = t_r18_c19_0 + p_17_18;
  assign t_r18_c19_6 = t_r18_c19_1 + p_17_20;
  assign t_r18_c19_7 = t_r18_c19_2 + t_r18_c19_3;
  assign t_r18_c19_8 = t_r18_c19_4 + p_19_18;
  assign t_r18_c19_9 = t_r18_c19_5 + t_r18_c19_6;
  assign t_r18_c19_10 = t_r18_c19_7 + t_r18_c19_8;
  assign t_r18_c19_11 = t_r18_c19_9 + t_r18_c19_10;
  assign t_r18_c19_12 = t_r18_c19_11 + p_19_20;
  assign out_18_19 = t_r18_c19_12 >> 4;

  assign t_r18_c20_0 = p_17_20 << 1;
  assign t_r18_c20_1 = p_18_19 << 1;
  assign t_r18_c20_2 = p_18_20 << 2;
  assign t_r18_c20_3 = p_18_21 << 1;
  assign t_r18_c20_4 = p_19_20 << 1;
  assign t_r18_c20_5 = t_r18_c20_0 + p_17_19;
  assign t_r18_c20_6 = t_r18_c20_1 + p_17_21;
  assign t_r18_c20_7 = t_r18_c20_2 + t_r18_c20_3;
  assign t_r18_c20_8 = t_r18_c20_4 + p_19_19;
  assign t_r18_c20_9 = t_r18_c20_5 + t_r18_c20_6;
  assign t_r18_c20_10 = t_r18_c20_7 + t_r18_c20_8;
  assign t_r18_c20_11 = t_r18_c20_9 + t_r18_c20_10;
  assign t_r18_c20_12 = t_r18_c20_11 + p_19_21;
  assign out_18_20 = t_r18_c20_12 >> 4;

  assign t_r18_c21_0 = p_17_21 << 1;
  assign t_r18_c21_1 = p_18_20 << 1;
  assign t_r18_c21_2 = p_18_21 << 2;
  assign t_r18_c21_3 = p_18_22 << 1;
  assign t_r18_c21_4 = p_19_21 << 1;
  assign t_r18_c21_5 = t_r18_c21_0 + p_17_20;
  assign t_r18_c21_6 = t_r18_c21_1 + p_17_22;
  assign t_r18_c21_7 = t_r18_c21_2 + t_r18_c21_3;
  assign t_r18_c21_8 = t_r18_c21_4 + p_19_20;
  assign t_r18_c21_9 = t_r18_c21_5 + t_r18_c21_6;
  assign t_r18_c21_10 = t_r18_c21_7 + t_r18_c21_8;
  assign t_r18_c21_11 = t_r18_c21_9 + t_r18_c21_10;
  assign t_r18_c21_12 = t_r18_c21_11 + p_19_22;
  assign out_18_21 = t_r18_c21_12 >> 4;

  assign t_r18_c22_0 = p_17_22 << 1;
  assign t_r18_c22_1 = p_18_21 << 1;
  assign t_r18_c22_2 = p_18_22 << 2;
  assign t_r18_c22_3 = p_18_23 << 1;
  assign t_r18_c22_4 = p_19_22 << 1;
  assign t_r18_c22_5 = t_r18_c22_0 + p_17_21;
  assign t_r18_c22_6 = t_r18_c22_1 + p_17_23;
  assign t_r18_c22_7 = t_r18_c22_2 + t_r18_c22_3;
  assign t_r18_c22_8 = t_r18_c22_4 + p_19_21;
  assign t_r18_c22_9 = t_r18_c22_5 + t_r18_c22_6;
  assign t_r18_c22_10 = t_r18_c22_7 + t_r18_c22_8;
  assign t_r18_c22_11 = t_r18_c22_9 + t_r18_c22_10;
  assign t_r18_c22_12 = t_r18_c22_11 + p_19_23;
  assign out_18_22 = t_r18_c22_12 >> 4;

  assign t_r18_c23_0 = p_17_23 << 1;
  assign t_r18_c23_1 = p_18_22 << 1;
  assign t_r18_c23_2 = p_18_23 << 2;
  assign t_r18_c23_3 = p_18_24 << 1;
  assign t_r18_c23_4 = p_19_23 << 1;
  assign t_r18_c23_5 = t_r18_c23_0 + p_17_22;
  assign t_r18_c23_6 = t_r18_c23_1 + p_17_24;
  assign t_r18_c23_7 = t_r18_c23_2 + t_r18_c23_3;
  assign t_r18_c23_8 = t_r18_c23_4 + p_19_22;
  assign t_r18_c23_9 = t_r18_c23_5 + t_r18_c23_6;
  assign t_r18_c23_10 = t_r18_c23_7 + t_r18_c23_8;
  assign t_r18_c23_11 = t_r18_c23_9 + t_r18_c23_10;
  assign t_r18_c23_12 = t_r18_c23_11 + p_19_24;
  assign out_18_23 = t_r18_c23_12 >> 4;

  assign t_r18_c24_0 = p_17_24 << 1;
  assign t_r18_c24_1 = p_18_23 << 1;
  assign t_r18_c24_2 = p_18_24 << 2;
  assign t_r18_c24_3 = p_18_25 << 1;
  assign t_r18_c24_4 = p_19_24 << 1;
  assign t_r18_c24_5 = t_r18_c24_0 + p_17_23;
  assign t_r18_c24_6 = t_r18_c24_1 + p_17_25;
  assign t_r18_c24_7 = t_r18_c24_2 + t_r18_c24_3;
  assign t_r18_c24_8 = t_r18_c24_4 + p_19_23;
  assign t_r18_c24_9 = t_r18_c24_5 + t_r18_c24_6;
  assign t_r18_c24_10 = t_r18_c24_7 + t_r18_c24_8;
  assign t_r18_c24_11 = t_r18_c24_9 + t_r18_c24_10;
  assign t_r18_c24_12 = t_r18_c24_11 + p_19_25;
  assign out_18_24 = t_r18_c24_12 >> 4;

  assign t_r18_c25_0 = p_17_25 << 1;
  assign t_r18_c25_1 = p_18_24 << 1;
  assign t_r18_c25_2 = p_18_25 << 2;
  assign t_r18_c25_3 = p_18_26 << 1;
  assign t_r18_c25_4 = p_19_25 << 1;
  assign t_r18_c25_5 = t_r18_c25_0 + p_17_24;
  assign t_r18_c25_6 = t_r18_c25_1 + p_17_26;
  assign t_r18_c25_7 = t_r18_c25_2 + t_r18_c25_3;
  assign t_r18_c25_8 = t_r18_c25_4 + p_19_24;
  assign t_r18_c25_9 = t_r18_c25_5 + t_r18_c25_6;
  assign t_r18_c25_10 = t_r18_c25_7 + t_r18_c25_8;
  assign t_r18_c25_11 = t_r18_c25_9 + t_r18_c25_10;
  assign t_r18_c25_12 = t_r18_c25_11 + p_19_26;
  assign out_18_25 = t_r18_c25_12 >> 4;

  assign t_r18_c26_0 = p_17_26 << 1;
  assign t_r18_c26_1 = p_18_25 << 1;
  assign t_r18_c26_2 = p_18_26 << 2;
  assign t_r18_c26_3 = p_18_27 << 1;
  assign t_r18_c26_4 = p_19_26 << 1;
  assign t_r18_c26_5 = t_r18_c26_0 + p_17_25;
  assign t_r18_c26_6 = t_r18_c26_1 + p_17_27;
  assign t_r18_c26_7 = t_r18_c26_2 + t_r18_c26_3;
  assign t_r18_c26_8 = t_r18_c26_4 + p_19_25;
  assign t_r18_c26_9 = t_r18_c26_5 + t_r18_c26_6;
  assign t_r18_c26_10 = t_r18_c26_7 + t_r18_c26_8;
  assign t_r18_c26_11 = t_r18_c26_9 + t_r18_c26_10;
  assign t_r18_c26_12 = t_r18_c26_11 + p_19_27;
  assign out_18_26 = t_r18_c26_12 >> 4;

  assign t_r18_c27_0 = p_17_27 << 1;
  assign t_r18_c27_1 = p_18_26 << 1;
  assign t_r18_c27_2 = p_18_27 << 2;
  assign t_r18_c27_3 = p_18_28 << 1;
  assign t_r18_c27_4 = p_19_27 << 1;
  assign t_r18_c27_5 = t_r18_c27_0 + p_17_26;
  assign t_r18_c27_6 = t_r18_c27_1 + p_17_28;
  assign t_r18_c27_7 = t_r18_c27_2 + t_r18_c27_3;
  assign t_r18_c27_8 = t_r18_c27_4 + p_19_26;
  assign t_r18_c27_9 = t_r18_c27_5 + t_r18_c27_6;
  assign t_r18_c27_10 = t_r18_c27_7 + t_r18_c27_8;
  assign t_r18_c27_11 = t_r18_c27_9 + t_r18_c27_10;
  assign t_r18_c27_12 = t_r18_c27_11 + p_19_28;
  assign out_18_27 = t_r18_c27_12 >> 4;

  assign t_r18_c28_0 = p_17_28 << 1;
  assign t_r18_c28_1 = p_18_27 << 1;
  assign t_r18_c28_2 = p_18_28 << 2;
  assign t_r18_c28_3 = p_18_29 << 1;
  assign t_r18_c28_4 = p_19_28 << 1;
  assign t_r18_c28_5 = t_r18_c28_0 + p_17_27;
  assign t_r18_c28_6 = t_r18_c28_1 + p_17_29;
  assign t_r18_c28_7 = t_r18_c28_2 + t_r18_c28_3;
  assign t_r18_c28_8 = t_r18_c28_4 + p_19_27;
  assign t_r18_c28_9 = t_r18_c28_5 + t_r18_c28_6;
  assign t_r18_c28_10 = t_r18_c28_7 + t_r18_c28_8;
  assign t_r18_c28_11 = t_r18_c28_9 + t_r18_c28_10;
  assign t_r18_c28_12 = t_r18_c28_11 + p_19_29;
  assign out_18_28 = t_r18_c28_12 >> 4;

  assign t_r18_c29_0 = p_17_29 << 1;
  assign t_r18_c29_1 = p_18_28 << 1;
  assign t_r18_c29_2 = p_18_29 << 2;
  assign t_r18_c29_3 = p_18_30 << 1;
  assign t_r18_c29_4 = p_19_29 << 1;
  assign t_r18_c29_5 = t_r18_c29_0 + p_17_28;
  assign t_r18_c29_6 = t_r18_c29_1 + p_17_30;
  assign t_r18_c29_7 = t_r18_c29_2 + t_r18_c29_3;
  assign t_r18_c29_8 = t_r18_c29_4 + p_19_28;
  assign t_r18_c29_9 = t_r18_c29_5 + t_r18_c29_6;
  assign t_r18_c29_10 = t_r18_c29_7 + t_r18_c29_8;
  assign t_r18_c29_11 = t_r18_c29_9 + t_r18_c29_10;
  assign t_r18_c29_12 = t_r18_c29_11 + p_19_30;
  assign out_18_29 = t_r18_c29_12 >> 4;

  assign t_r18_c30_0 = p_17_30 << 1;
  assign t_r18_c30_1 = p_18_29 << 1;
  assign t_r18_c30_2 = p_18_30 << 2;
  assign t_r18_c30_3 = p_18_31 << 1;
  assign t_r18_c30_4 = p_19_30 << 1;
  assign t_r18_c30_5 = t_r18_c30_0 + p_17_29;
  assign t_r18_c30_6 = t_r18_c30_1 + p_17_31;
  assign t_r18_c30_7 = t_r18_c30_2 + t_r18_c30_3;
  assign t_r18_c30_8 = t_r18_c30_4 + p_19_29;
  assign t_r18_c30_9 = t_r18_c30_5 + t_r18_c30_6;
  assign t_r18_c30_10 = t_r18_c30_7 + t_r18_c30_8;
  assign t_r18_c30_11 = t_r18_c30_9 + t_r18_c30_10;
  assign t_r18_c30_12 = t_r18_c30_11 + p_19_31;
  assign out_18_30 = t_r18_c30_12 >> 4;

  assign t_r18_c31_0 = p_17_31 << 1;
  assign t_r18_c31_1 = p_18_30 << 1;
  assign t_r18_c31_2 = p_18_31 << 2;
  assign t_r18_c31_3 = p_18_32 << 1;
  assign t_r18_c31_4 = p_19_31 << 1;
  assign t_r18_c31_5 = t_r18_c31_0 + p_17_30;
  assign t_r18_c31_6 = t_r18_c31_1 + p_17_32;
  assign t_r18_c31_7 = t_r18_c31_2 + t_r18_c31_3;
  assign t_r18_c31_8 = t_r18_c31_4 + p_19_30;
  assign t_r18_c31_9 = t_r18_c31_5 + t_r18_c31_6;
  assign t_r18_c31_10 = t_r18_c31_7 + t_r18_c31_8;
  assign t_r18_c31_11 = t_r18_c31_9 + t_r18_c31_10;
  assign t_r18_c31_12 = t_r18_c31_11 + p_19_32;
  assign out_18_31 = t_r18_c31_12 >> 4;

  assign t_r18_c32_0 = p_17_32 << 1;
  assign t_r18_c32_1 = p_18_31 << 1;
  assign t_r18_c32_2 = p_18_32 << 2;
  assign t_r18_c32_3 = p_18_33 << 1;
  assign t_r18_c32_4 = p_19_32 << 1;
  assign t_r18_c32_5 = t_r18_c32_0 + p_17_31;
  assign t_r18_c32_6 = t_r18_c32_1 + p_17_33;
  assign t_r18_c32_7 = t_r18_c32_2 + t_r18_c32_3;
  assign t_r18_c32_8 = t_r18_c32_4 + p_19_31;
  assign t_r18_c32_9 = t_r18_c32_5 + t_r18_c32_6;
  assign t_r18_c32_10 = t_r18_c32_7 + t_r18_c32_8;
  assign t_r18_c32_11 = t_r18_c32_9 + t_r18_c32_10;
  assign t_r18_c32_12 = t_r18_c32_11 + p_19_33;
  assign out_18_32 = t_r18_c32_12 >> 4;

  assign t_r18_c33_0 = p_17_33 << 1;
  assign t_r18_c33_1 = p_18_32 << 1;
  assign t_r18_c33_2 = p_18_33 << 2;
  assign t_r18_c33_3 = p_18_34 << 1;
  assign t_r18_c33_4 = p_19_33 << 1;
  assign t_r18_c33_5 = t_r18_c33_0 + p_17_32;
  assign t_r18_c33_6 = t_r18_c33_1 + p_17_34;
  assign t_r18_c33_7 = t_r18_c33_2 + t_r18_c33_3;
  assign t_r18_c33_8 = t_r18_c33_4 + p_19_32;
  assign t_r18_c33_9 = t_r18_c33_5 + t_r18_c33_6;
  assign t_r18_c33_10 = t_r18_c33_7 + t_r18_c33_8;
  assign t_r18_c33_11 = t_r18_c33_9 + t_r18_c33_10;
  assign t_r18_c33_12 = t_r18_c33_11 + p_19_34;
  assign out_18_33 = t_r18_c33_12 >> 4;

  assign t_r18_c34_0 = p_17_34 << 1;
  assign t_r18_c34_1 = p_18_33 << 1;
  assign t_r18_c34_2 = p_18_34 << 2;
  assign t_r18_c34_3 = p_18_35 << 1;
  assign t_r18_c34_4 = p_19_34 << 1;
  assign t_r18_c34_5 = t_r18_c34_0 + p_17_33;
  assign t_r18_c34_6 = t_r18_c34_1 + p_17_35;
  assign t_r18_c34_7 = t_r18_c34_2 + t_r18_c34_3;
  assign t_r18_c34_8 = t_r18_c34_4 + p_19_33;
  assign t_r18_c34_9 = t_r18_c34_5 + t_r18_c34_6;
  assign t_r18_c34_10 = t_r18_c34_7 + t_r18_c34_8;
  assign t_r18_c34_11 = t_r18_c34_9 + t_r18_c34_10;
  assign t_r18_c34_12 = t_r18_c34_11 + p_19_35;
  assign out_18_34 = t_r18_c34_12 >> 4;

  assign t_r18_c35_0 = p_17_35 << 1;
  assign t_r18_c35_1 = p_18_34 << 1;
  assign t_r18_c35_2 = p_18_35 << 2;
  assign t_r18_c35_3 = p_18_36 << 1;
  assign t_r18_c35_4 = p_19_35 << 1;
  assign t_r18_c35_5 = t_r18_c35_0 + p_17_34;
  assign t_r18_c35_6 = t_r18_c35_1 + p_17_36;
  assign t_r18_c35_7 = t_r18_c35_2 + t_r18_c35_3;
  assign t_r18_c35_8 = t_r18_c35_4 + p_19_34;
  assign t_r18_c35_9 = t_r18_c35_5 + t_r18_c35_6;
  assign t_r18_c35_10 = t_r18_c35_7 + t_r18_c35_8;
  assign t_r18_c35_11 = t_r18_c35_9 + t_r18_c35_10;
  assign t_r18_c35_12 = t_r18_c35_11 + p_19_36;
  assign out_18_35 = t_r18_c35_12 >> 4;

  assign t_r18_c36_0 = p_17_36 << 1;
  assign t_r18_c36_1 = p_18_35 << 1;
  assign t_r18_c36_2 = p_18_36 << 2;
  assign t_r18_c36_3 = p_18_37 << 1;
  assign t_r18_c36_4 = p_19_36 << 1;
  assign t_r18_c36_5 = t_r18_c36_0 + p_17_35;
  assign t_r18_c36_6 = t_r18_c36_1 + p_17_37;
  assign t_r18_c36_7 = t_r18_c36_2 + t_r18_c36_3;
  assign t_r18_c36_8 = t_r18_c36_4 + p_19_35;
  assign t_r18_c36_9 = t_r18_c36_5 + t_r18_c36_6;
  assign t_r18_c36_10 = t_r18_c36_7 + t_r18_c36_8;
  assign t_r18_c36_11 = t_r18_c36_9 + t_r18_c36_10;
  assign t_r18_c36_12 = t_r18_c36_11 + p_19_37;
  assign out_18_36 = t_r18_c36_12 >> 4;

  assign t_r18_c37_0 = p_17_37 << 1;
  assign t_r18_c37_1 = p_18_36 << 1;
  assign t_r18_c37_2 = p_18_37 << 2;
  assign t_r18_c37_3 = p_18_38 << 1;
  assign t_r18_c37_4 = p_19_37 << 1;
  assign t_r18_c37_5 = t_r18_c37_0 + p_17_36;
  assign t_r18_c37_6 = t_r18_c37_1 + p_17_38;
  assign t_r18_c37_7 = t_r18_c37_2 + t_r18_c37_3;
  assign t_r18_c37_8 = t_r18_c37_4 + p_19_36;
  assign t_r18_c37_9 = t_r18_c37_5 + t_r18_c37_6;
  assign t_r18_c37_10 = t_r18_c37_7 + t_r18_c37_8;
  assign t_r18_c37_11 = t_r18_c37_9 + t_r18_c37_10;
  assign t_r18_c37_12 = t_r18_c37_11 + p_19_38;
  assign out_18_37 = t_r18_c37_12 >> 4;

  assign t_r18_c38_0 = p_17_38 << 1;
  assign t_r18_c38_1 = p_18_37 << 1;
  assign t_r18_c38_2 = p_18_38 << 2;
  assign t_r18_c38_3 = p_18_39 << 1;
  assign t_r18_c38_4 = p_19_38 << 1;
  assign t_r18_c38_5 = t_r18_c38_0 + p_17_37;
  assign t_r18_c38_6 = t_r18_c38_1 + p_17_39;
  assign t_r18_c38_7 = t_r18_c38_2 + t_r18_c38_3;
  assign t_r18_c38_8 = t_r18_c38_4 + p_19_37;
  assign t_r18_c38_9 = t_r18_c38_5 + t_r18_c38_6;
  assign t_r18_c38_10 = t_r18_c38_7 + t_r18_c38_8;
  assign t_r18_c38_11 = t_r18_c38_9 + t_r18_c38_10;
  assign t_r18_c38_12 = t_r18_c38_11 + p_19_39;
  assign out_18_38 = t_r18_c38_12 >> 4;

  assign t_r18_c39_0 = p_17_39 << 1;
  assign t_r18_c39_1 = p_18_38 << 1;
  assign t_r18_c39_2 = p_18_39 << 2;
  assign t_r18_c39_3 = p_18_40 << 1;
  assign t_r18_c39_4 = p_19_39 << 1;
  assign t_r18_c39_5 = t_r18_c39_0 + p_17_38;
  assign t_r18_c39_6 = t_r18_c39_1 + p_17_40;
  assign t_r18_c39_7 = t_r18_c39_2 + t_r18_c39_3;
  assign t_r18_c39_8 = t_r18_c39_4 + p_19_38;
  assign t_r18_c39_9 = t_r18_c39_5 + t_r18_c39_6;
  assign t_r18_c39_10 = t_r18_c39_7 + t_r18_c39_8;
  assign t_r18_c39_11 = t_r18_c39_9 + t_r18_c39_10;
  assign t_r18_c39_12 = t_r18_c39_11 + p_19_40;
  assign out_18_39 = t_r18_c39_12 >> 4;

  assign t_r18_c40_0 = p_17_40 << 1;
  assign t_r18_c40_1 = p_18_39 << 1;
  assign t_r18_c40_2 = p_18_40 << 2;
  assign t_r18_c40_3 = p_18_41 << 1;
  assign t_r18_c40_4 = p_19_40 << 1;
  assign t_r18_c40_5 = t_r18_c40_0 + p_17_39;
  assign t_r18_c40_6 = t_r18_c40_1 + p_17_41;
  assign t_r18_c40_7 = t_r18_c40_2 + t_r18_c40_3;
  assign t_r18_c40_8 = t_r18_c40_4 + p_19_39;
  assign t_r18_c40_9 = t_r18_c40_5 + t_r18_c40_6;
  assign t_r18_c40_10 = t_r18_c40_7 + t_r18_c40_8;
  assign t_r18_c40_11 = t_r18_c40_9 + t_r18_c40_10;
  assign t_r18_c40_12 = t_r18_c40_11 + p_19_41;
  assign out_18_40 = t_r18_c40_12 >> 4;

  assign t_r18_c41_0 = p_17_41 << 1;
  assign t_r18_c41_1 = p_18_40 << 1;
  assign t_r18_c41_2 = p_18_41 << 2;
  assign t_r18_c41_3 = p_18_42 << 1;
  assign t_r18_c41_4 = p_19_41 << 1;
  assign t_r18_c41_5 = t_r18_c41_0 + p_17_40;
  assign t_r18_c41_6 = t_r18_c41_1 + p_17_42;
  assign t_r18_c41_7 = t_r18_c41_2 + t_r18_c41_3;
  assign t_r18_c41_8 = t_r18_c41_4 + p_19_40;
  assign t_r18_c41_9 = t_r18_c41_5 + t_r18_c41_6;
  assign t_r18_c41_10 = t_r18_c41_7 + t_r18_c41_8;
  assign t_r18_c41_11 = t_r18_c41_9 + t_r18_c41_10;
  assign t_r18_c41_12 = t_r18_c41_11 + p_19_42;
  assign out_18_41 = t_r18_c41_12 >> 4;

  assign t_r18_c42_0 = p_17_42 << 1;
  assign t_r18_c42_1 = p_18_41 << 1;
  assign t_r18_c42_2 = p_18_42 << 2;
  assign t_r18_c42_3 = p_18_43 << 1;
  assign t_r18_c42_4 = p_19_42 << 1;
  assign t_r18_c42_5 = t_r18_c42_0 + p_17_41;
  assign t_r18_c42_6 = t_r18_c42_1 + p_17_43;
  assign t_r18_c42_7 = t_r18_c42_2 + t_r18_c42_3;
  assign t_r18_c42_8 = t_r18_c42_4 + p_19_41;
  assign t_r18_c42_9 = t_r18_c42_5 + t_r18_c42_6;
  assign t_r18_c42_10 = t_r18_c42_7 + t_r18_c42_8;
  assign t_r18_c42_11 = t_r18_c42_9 + t_r18_c42_10;
  assign t_r18_c42_12 = t_r18_c42_11 + p_19_43;
  assign out_18_42 = t_r18_c42_12 >> 4;

  assign t_r18_c43_0 = p_17_43 << 1;
  assign t_r18_c43_1 = p_18_42 << 1;
  assign t_r18_c43_2 = p_18_43 << 2;
  assign t_r18_c43_3 = p_18_44 << 1;
  assign t_r18_c43_4 = p_19_43 << 1;
  assign t_r18_c43_5 = t_r18_c43_0 + p_17_42;
  assign t_r18_c43_6 = t_r18_c43_1 + p_17_44;
  assign t_r18_c43_7 = t_r18_c43_2 + t_r18_c43_3;
  assign t_r18_c43_8 = t_r18_c43_4 + p_19_42;
  assign t_r18_c43_9 = t_r18_c43_5 + t_r18_c43_6;
  assign t_r18_c43_10 = t_r18_c43_7 + t_r18_c43_8;
  assign t_r18_c43_11 = t_r18_c43_9 + t_r18_c43_10;
  assign t_r18_c43_12 = t_r18_c43_11 + p_19_44;
  assign out_18_43 = t_r18_c43_12 >> 4;

  assign t_r18_c44_0 = p_17_44 << 1;
  assign t_r18_c44_1 = p_18_43 << 1;
  assign t_r18_c44_2 = p_18_44 << 2;
  assign t_r18_c44_3 = p_18_45 << 1;
  assign t_r18_c44_4 = p_19_44 << 1;
  assign t_r18_c44_5 = t_r18_c44_0 + p_17_43;
  assign t_r18_c44_6 = t_r18_c44_1 + p_17_45;
  assign t_r18_c44_7 = t_r18_c44_2 + t_r18_c44_3;
  assign t_r18_c44_8 = t_r18_c44_4 + p_19_43;
  assign t_r18_c44_9 = t_r18_c44_5 + t_r18_c44_6;
  assign t_r18_c44_10 = t_r18_c44_7 + t_r18_c44_8;
  assign t_r18_c44_11 = t_r18_c44_9 + t_r18_c44_10;
  assign t_r18_c44_12 = t_r18_c44_11 + p_19_45;
  assign out_18_44 = t_r18_c44_12 >> 4;

  assign t_r18_c45_0 = p_17_45 << 1;
  assign t_r18_c45_1 = p_18_44 << 1;
  assign t_r18_c45_2 = p_18_45 << 2;
  assign t_r18_c45_3 = p_18_46 << 1;
  assign t_r18_c45_4 = p_19_45 << 1;
  assign t_r18_c45_5 = t_r18_c45_0 + p_17_44;
  assign t_r18_c45_6 = t_r18_c45_1 + p_17_46;
  assign t_r18_c45_7 = t_r18_c45_2 + t_r18_c45_3;
  assign t_r18_c45_8 = t_r18_c45_4 + p_19_44;
  assign t_r18_c45_9 = t_r18_c45_5 + t_r18_c45_6;
  assign t_r18_c45_10 = t_r18_c45_7 + t_r18_c45_8;
  assign t_r18_c45_11 = t_r18_c45_9 + t_r18_c45_10;
  assign t_r18_c45_12 = t_r18_c45_11 + p_19_46;
  assign out_18_45 = t_r18_c45_12 >> 4;

  assign t_r18_c46_0 = p_17_46 << 1;
  assign t_r18_c46_1 = p_18_45 << 1;
  assign t_r18_c46_2 = p_18_46 << 2;
  assign t_r18_c46_3 = p_18_47 << 1;
  assign t_r18_c46_4 = p_19_46 << 1;
  assign t_r18_c46_5 = t_r18_c46_0 + p_17_45;
  assign t_r18_c46_6 = t_r18_c46_1 + p_17_47;
  assign t_r18_c46_7 = t_r18_c46_2 + t_r18_c46_3;
  assign t_r18_c46_8 = t_r18_c46_4 + p_19_45;
  assign t_r18_c46_9 = t_r18_c46_5 + t_r18_c46_6;
  assign t_r18_c46_10 = t_r18_c46_7 + t_r18_c46_8;
  assign t_r18_c46_11 = t_r18_c46_9 + t_r18_c46_10;
  assign t_r18_c46_12 = t_r18_c46_11 + p_19_47;
  assign out_18_46 = t_r18_c46_12 >> 4;

  assign t_r18_c47_0 = p_17_47 << 1;
  assign t_r18_c47_1 = p_18_46 << 1;
  assign t_r18_c47_2 = p_18_47 << 2;
  assign t_r18_c47_3 = p_18_48 << 1;
  assign t_r18_c47_4 = p_19_47 << 1;
  assign t_r18_c47_5 = t_r18_c47_0 + p_17_46;
  assign t_r18_c47_6 = t_r18_c47_1 + p_17_48;
  assign t_r18_c47_7 = t_r18_c47_2 + t_r18_c47_3;
  assign t_r18_c47_8 = t_r18_c47_4 + p_19_46;
  assign t_r18_c47_9 = t_r18_c47_5 + t_r18_c47_6;
  assign t_r18_c47_10 = t_r18_c47_7 + t_r18_c47_8;
  assign t_r18_c47_11 = t_r18_c47_9 + t_r18_c47_10;
  assign t_r18_c47_12 = t_r18_c47_11 + p_19_48;
  assign out_18_47 = t_r18_c47_12 >> 4;

  assign t_r18_c48_0 = p_17_48 << 1;
  assign t_r18_c48_1 = p_18_47 << 1;
  assign t_r18_c48_2 = p_18_48 << 2;
  assign t_r18_c48_3 = p_18_49 << 1;
  assign t_r18_c48_4 = p_19_48 << 1;
  assign t_r18_c48_5 = t_r18_c48_0 + p_17_47;
  assign t_r18_c48_6 = t_r18_c48_1 + p_17_49;
  assign t_r18_c48_7 = t_r18_c48_2 + t_r18_c48_3;
  assign t_r18_c48_8 = t_r18_c48_4 + p_19_47;
  assign t_r18_c48_9 = t_r18_c48_5 + t_r18_c48_6;
  assign t_r18_c48_10 = t_r18_c48_7 + t_r18_c48_8;
  assign t_r18_c48_11 = t_r18_c48_9 + t_r18_c48_10;
  assign t_r18_c48_12 = t_r18_c48_11 + p_19_49;
  assign out_18_48 = t_r18_c48_12 >> 4;

  assign t_r18_c49_0 = p_17_49 << 1;
  assign t_r18_c49_1 = p_18_48 << 1;
  assign t_r18_c49_2 = p_18_49 << 2;
  assign t_r18_c49_3 = p_18_50 << 1;
  assign t_r18_c49_4 = p_19_49 << 1;
  assign t_r18_c49_5 = t_r18_c49_0 + p_17_48;
  assign t_r18_c49_6 = t_r18_c49_1 + p_17_50;
  assign t_r18_c49_7 = t_r18_c49_2 + t_r18_c49_3;
  assign t_r18_c49_8 = t_r18_c49_4 + p_19_48;
  assign t_r18_c49_9 = t_r18_c49_5 + t_r18_c49_6;
  assign t_r18_c49_10 = t_r18_c49_7 + t_r18_c49_8;
  assign t_r18_c49_11 = t_r18_c49_9 + t_r18_c49_10;
  assign t_r18_c49_12 = t_r18_c49_11 + p_19_50;
  assign out_18_49 = t_r18_c49_12 >> 4;

  assign t_r18_c50_0 = p_17_50 << 1;
  assign t_r18_c50_1 = p_18_49 << 1;
  assign t_r18_c50_2 = p_18_50 << 2;
  assign t_r18_c50_3 = p_18_51 << 1;
  assign t_r18_c50_4 = p_19_50 << 1;
  assign t_r18_c50_5 = t_r18_c50_0 + p_17_49;
  assign t_r18_c50_6 = t_r18_c50_1 + p_17_51;
  assign t_r18_c50_7 = t_r18_c50_2 + t_r18_c50_3;
  assign t_r18_c50_8 = t_r18_c50_4 + p_19_49;
  assign t_r18_c50_9 = t_r18_c50_5 + t_r18_c50_6;
  assign t_r18_c50_10 = t_r18_c50_7 + t_r18_c50_8;
  assign t_r18_c50_11 = t_r18_c50_9 + t_r18_c50_10;
  assign t_r18_c50_12 = t_r18_c50_11 + p_19_51;
  assign out_18_50 = t_r18_c50_12 >> 4;

  assign t_r18_c51_0 = p_17_51 << 1;
  assign t_r18_c51_1 = p_18_50 << 1;
  assign t_r18_c51_2 = p_18_51 << 2;
  assign t_r18_c51_3 = p_18_52 << 1;
  assign t_r18_c51_4 = p_19_51 << 1;
  assign t_r18_c51_5 = t_r18_c51_0 + p_17_50;
  assign t_r18_c51_6 = t_r18_c51_1 + p_17_52;
  assign t_r18_c51_7 = t_r18_c51_2 + t_r18_c51_3;
  assign t_r18_c51_8 = t_r18_c51_4 + p_19_50;
  assign t_r18_c51_9 = t_r18_c51_5 + t_r18_c51_6;
  assign t_r18_c51_10 = t_r18_c51_7 + t_r18_c51_8;
  assign t_r18_c51_11 = t_r18_c51_9 + t_r18_c51_10;
  assign t_r18_c51_12 = t_r18_c51_11 + p_19_52;
  assign out_18_51 = t_r18_c51_12 >> 4;

  assign t_r18_c52_0 = p_17_52 << 1;
  assign t_r18_c52_1 = p_18_51 << 1;
  assign t_r18_c52_2 = p_18_52 << 2;
  assign t_r18_c52_3 = p_18_53 << 1;
  assign t_r18_c52_4 = p_19_52 << 1;
  assign t_r18_c52_5 = t_r18_c52_0 + p_17_51;
  assign t_r18_c52_6 = t_r18_c52_1 + p_17_53;
  assign t_r18_c52_7 = t_r18_c52_2 + t_r18_c52_3;
  assign t_r18_c52_8 = t_r18_c52_4 + p_19_51;
  assign t_r18_c52_9 = t_r18_c52_5 + t_r18_c52_6;
  assign t_r18_c52_10 = t_r18_c52_7 + t_r18_c52_8;
  assign t_r18_c52_11 = t_r18_c52_9 + t_r18_c52_10;
  assign t_r18_c52_12 = t_r18_c52_11 + p_19_53;
  assign out_18_52 = t_r18_c52_12 >> 4;

  assign t_r18_c53_0 = p_17_53 << 1;
  assign t_r18_c53_1 = p_18_52 << 1;
  assign t_r18_c53_2 = p_18_53 << 2;
  assign t_r18_c53_3 = p_18_54 << 1;
  assign t_r18_c53_4 = p_19_53 << 1;
  assign t_r18_c53_5 = t_r18_c53_0 + p_17_52;
  assign t_r18_c53_6 = t_r18_c53_1 + p_17_54;
  assign t_r18_c53_7 = t_r18_c53_2 + t_r18_c53_3;
  assign t_r18_c53_8 = t_r18_c53_4 + p_19_52;
  assign t_r18_c53_9 = t_r18_c53_5 + t_r18_c53_6;
  assign t_r18_c53_10 = t_r18_c53_7 + t_r18_c53_8;
  assign t_r18_c53_11 = t_r18_c53_9 + t_r18_c53_10;
  assign t_r18_c53_12 = t_r18_c53_11 + p_19_54;
  assign out_18_53 = t_r18_c53_12 >> 4;

  assign t_r18_c54_0 = p_17_54 << 1;
  assign t_r18_c54_1 = p_18_53 << 1;
  assign t_r18_c54_2 = p_18_54 << 2;
  assign t_r18_c54_3 = p_18_55 << 1;
  assign t_r18_c54_4 = p_19_54 << 1;
  assign t_r18_c54_5 = t_r18_c54_0 + p_17_53;
  assign t_r18_c54_6 = t_r18_c54_1 + p_17_55;
  assign t_r18_c54_7 = t_r18_c54_2 + t_r18_c54_3;
  assign t_r18_c54_8 = t_r18_c54_4 + p_19_53;
  assign t_r18_c54_9 = t_r18_c54_5 + t_r18_c54_6;
  assign t_r18_c54_10 = t_r18_c54_7 + t_r18_c54_8;
  assign t_r18_c54_11 = t_r18_c54_9 + t_r18_c54_10;
  assign t_r18_c54_12 = t_r18_c54_11 + p_19_55;
  assign out_18_54 = t_r18_c54_12 >> 4;

  assign t_r18_c55_0 = p_17_55 << 1;
  assign t_r18_c55_1 = p_18_54 << 1;
  assign t_r18_c55_2 = p_18_55 << 2;
  assign t_r18_c55_3 = p_18_56 << 1;
  assign t_r18_c55_4 = p_19_55 << 1;
  assign t_r18_c55_5 = t_r18_c55_0 + p_17_54;
  assign t_r18_c55_6 = t_r18_c55_1 + p_17_56;
  assign t_r18_c55_7 = t_r18_c55_2 + t_r18_c55_3;
  assign t_r18_c55_8 = t_r18_c55_4 + p_19_54;
  assign t_r18_c55_9 = t_r18_c55_5 + t_r18_c55_6;
  assign t_r18_c55_10 = t_r18_c55_7 + t_r18_c55_8;
  assign t_r18_c55_11 = t_r18_c55_9 + t_r18_c55_10;
  assign t_r18_c55_12 = t_r18_c55_11 + p_19_56;
  assign out_18_55 = t_r18_c55_12 >> 4;

  assign t_r18_c56_0 = p_17_56 << 1;
  assign t_r18_c56_1 = p_18_55 << 1;
  assign t_r18_c56_2 = p_18_56 << 2;
  assign t_r18_c56_3 = p_18_57 << 1;
  assign t_r18_c56_4 = p_19_56 << 1;
  assign t_r18_c56_5 = t_r18_c56_0 + p_17_55;
  assign t_r18_c56_6 = t_r18_c56_1 + p_17_57;
  assign t_r18_c56_7 = t_r18_c56_2 + t_r18_c56_3;
  assign t_r18_c56_8 = t_r18_c56_4 + p_19_55;
  assign t_r18_c56_9 = t_r18_c56_5 + t_r18_c56_6;
  assign t_r18_c56_10 = t_r18_c56_7 + t_r18_c56_8;
  assign t_r18_c56_11 = t_r18_c56_9 + t_r18_c56_10;
  assign t_r18_c56_12 = t_r18_c56_11 + p_19_57;
  assign out_18_56 = t_r18_c56_12 >> 4;

  assign t_r18_c57_0 = p_17_57 << 1;
  assign t_r18_c57_1 = p_18_56 << 1;
  assign t_r18_c57_2 = p_18_57 << 2;
  assign t_r18_c57_3 = p_18_58 << 1;
  assign t_r18_c57_4 = p_19_57 << 1;
  assign t_r18_c57_5 = t_r18_c57_0 + p_17_56;
  assign t_r18_c57_6 = t_r18_c57_1 + p_17_58;
  assign t_r18_c57_7 = t_r18_c57_2 + t_r18_c57_3;
  assign t_r18_c57_8 = t_r18_c57_4 + p_19_56;
  assign t_r18_c57_9 = t_r18_c57_5 + t_r18_c57_6;
  assign t_r18_c57_10 = t_r18_c57_7 + t_r18_c57_8;
  assign t_r18_c57_11 = t_r18_c57_9 + t_r18_c57_10;
  assign t_r18_c57_12 = t_r18_c57_11 + p_19_58;
  assign out_18_57 = t_r18_c57_12 >> 4;

  assign t_r18_c58_0 = p_17_58 << 1;
  assign t_r18_c58_1 = p_18_57 << 1;
  assign t_r18_c58_2 = p_18_58 << 2;
  assign t_r18_c58_3 = p_18_59 << 1;
  assign t_r18_c58_4 = p_19_58 << 1;
  assign t_r18_c58_5 = t_r18_c58_0 + p_17_57;
  assign t_r18_c58_6 = t_r18_c58_1 + p_17_59;
  assign t_r18_c58_7 = t_r18_c58_2 + t_r18_c58_3;
  assign t_r18_c58_8 = t_r18_c58_4 + p_19_57;
  assign t_r18_c58_9 = t_r18_c58_5 + t_r18_c58_6;
  assign t_r18_c58_10 = t_r18_c58_7 + t_r18_c58_8;
  assign t_r18_c58_11 = t_r18_c58_9 + t_r18_c58_10;
  assign t_r18_c58_12 = t_r18_c58_11 + p_19_59;
  assign out_18_58 = t_r18_c58_12 >> 4;

  assign t_r18_c59_0 = p_17_59 << 1;
  assign t_r18_c59_1 = p_18_58 << 1;
  assign t_r18_c59_2 = p_18_59 << 2;
  assign t_r18_c59_3 = p_18_60 << 1;
  assign t_r18_c59_4 = p_19_59 << 1;
  assign t_r18_c59_5 = t_r18_c59_0 + p_17_58;
  assign t_r18_c59_6 = t_r18_c59_1 + p_17_60;
  assign t_r18_c59_7 = t_r18_c59_2 + t_r18_c59_3;
  assign t_r18_c59_8 = t_r18_c59_4 + p_19_58;
  assign t_r18_c59_9 = t_r18_c59_5 + t_r18_c59_6;
  assign t_r18_c59_10 = t_r18_c59_7 + t_r18_c59_8;
  assign t_r18_c59_11 = t_r18_c59_9 + t_r18_c59_10;
  assign t_r18_c59_12 = t_r18_c59_11 + p_19_60;
  assign out_18_59 = t_r18_c59_12 >> 4;

  assign t_r18_c60_0 = p_17_60 << 1;
  assign t_r18_c60_1 = p_18_59 << 1;
  assign t_r18_c60_2 = p_18_60 << 2;
  assign t_r18_c60_3 = p_18_61 << 1;
  assign t_r18_c60_4 = p_19_60 << 1;
  assign t_r18_c60_5 = t_r18_c60_0 + p_17_59;
  assign t_r18_c60_6 = t_r18_c60_1 + p_17_61;
  assign t_r18_c60_7 = t_r18_c60_2 + t_r18_c60_3;
  assign t_r18_c60_8 = t_r18_c60_4 + p_19_59;
  assign t_r18_c60_9 = t_r18_c60_5 + t_r18_c60_6;
  assign t_r18_c60_10 = t_r18_c60_7 + t_r18_c60_8;
  assign t_r18_c60_11 = t_r18_c60_9 + t_r18_c60_10;
  assign t_r18_c60_12 = t_r18_c60_11 + p_19_61;
  assign out_18_60 = t_r18_c60_12 >> 4;

  assign t_r18_c61_0 = p_17_61 << 1;
  assign t_r18_c61_1 = p_18_60 << 1;
  assign t_r18_c61_2 = p_18_61 << 2;
  assign t_r18_c61_3 = p_18_62 << 1;
  assign t_r18_c61_4 = p_19_61 << 1;
  assign t_r18_c61_5 = t_r18_c61_0 + p_17_60;
  assign t_r18_c61_6 = t_r18_c61_1 + p_17_62;
  assign t_r18_c61_7 = t_r18_c61_2 + t_r18_c61_3;
  assign t_r18_c61_8 = t_r18_c61_4 + p_19_60;
  assign t_r18_c61_9 = t_r18_c61_5 + t_r18_c61_6;
  assign t_r18_c61_10 = t_r18_c61_7 + t_r18_c61_8;
  assign t_r18_c61_11 = t_r18_c61_9 + t_r18_c61_10;
  assign t_r18_c61_12 = t_r18_c61_11 + p_19_62;
  assign out_18_61 = t_r18_c61_12 >> 4;

  assign t_r18_c62_0 = p_17_62 << 1;
  assign t_r18_c62_1 = p_18_61 << 1;
  assign t_r18_c62_2 = p_18_62 << 2;
  assign t_r18_c62_3 = p_18_63 << 1;
  assign t_r18_c62_4 = p_19_62 << 1;
  assign t_r18_c62_5 = t_r18_c62_0 + p_17_61;
  assign t_r18_c62_6 = t_r18_c62_1 + p_17_63;
  assign t_r18_c62_7 = t_r18_c62_2 + t_r18_c62_3;
  assign t_r18_c62_8 = t_r18_c62_4 + p_19_61;
  assign t_r18_c62_9 = t_r18_c62_5 + t_r18_c62_6;
  assign t_r18_c62_10 = t_r18_c62_7 + t_r18_c62_8;
  assign t_r18_c62_11 = t_r18_c62_9 + t_r18_c62_10;
  assign t_r18_c62_12 = t_r18_c62_11 + p_19_63;
  assign out_18_62 = t_r18_c62_12 >> 4;

  assign t_r18_c63_0 = p_17_63 << 1;
  assign t_r18_c63_1 = p_18_62 << 1;
  assign t_r18_c63_2 = p_18_63 << 2;
  assign t_r18_c63_3 = p_18_64 << 1;
  assign t_r18_c63_4 = p_19_63 << 1;
  assign t_r18_c63_5 = t_r18_c63_0 + p_17_62;
  assign t_r18_c63_6 = t_r18_c63_1 + p_17_64;
  assign t_r18_c63_7 = t_r18_c63_2 + t_r18_c63_3;
  assign t_r18_c63_8 = t_r18_c63_4 + p_19_62;
  assign t_r18_c63_9 = t_r18_c63_5 + t_r18_c63_6;
  assign t_r18_c63_10 = t_r18_c63_7 + t_r18_c63_8;
  assign t_r18_c63_11 = t_r18_c63_9 + t_r18_c63_10;
  assign t_r18_c63_12 = t_r18_c63_11 + p_19_64;
  assign out_18_63 = t_r18_c63_12 >> 4;

  assign t_r18_c64_0 = p_17_64 << 1;
  assign t_r18_c64_1 = p_18_63 << 1;
  assign t_r18_c64_2 = p_18_64 << 2;
  assign t_r18_c64_3 = p_18_65 << 1;
  assign t_r18_c64_4 = p_19_64 << 1;
  assign t_r18_c64_5 = t_r18_c64_0 + p_17_63;
  assign t_r18_c64_6 = t_r18_c64_1 + p_17_65;
  assign t_r18_c64_7 = t_r18_c64_2 + t_r18_c64_3;
  assign t_r18_c64_8 = t_r18_c64_4 + p_19_63;
  assign t_r18_c64_9 = t_r18_c64_5 + t_r18_c64_6;
  assign t_r18_c64_10 = t_r18_c64_7 + t_r18_c64_8;
  assign t_r18_c64_11 = t_r18_c64_9 + t_r18_c64_10;
  assign t_r18_c64_12 = t_r18_c64_11 + p_19_65;
  assign out_18_64 = t_r18_c64_12 >> 4;

  assign t_r19_c1_0 = p_18_1 << 1;
  assign t_r19_c1_1 = p_19_0 << 1;
  assign t_r19_c1_2 = p_19_1 << 2;
  assign t_r19_c1_3 = p_19_2 << 1;
  assign t_r19_c1_4 = p_20_1 << 1;
  assign t_r19_c1_5 = t_r19_c1_0 + p_18_0;
  assign t_r19_c1_6 = t_r19_c1_1 + p_18_2;
  assign t_r19_c1_7 = t_r19_c1_2 + t_r19_c1_3;
  assign t_r19_c1_8 = t_r19_c1_4 + p_20_0;
  assign t_r19_c1_9 = t_r19_c1_5 + t_r19_c1_6;
  assign t_r19_c1_10 = t_r19_c1_7 + t_r19_c1_8;
  assign t_r19_c1_11 = t_r19_c1_9 + t_r19_c1_10;
  assign t_r19_c1_12 = t_r19_c1_11 + p_20_2;
  assign out_19_1 = t_r19_c1_12 >> 4;

  assign t_r19_c2_0 = p_18_2 << 1;
  assign t_r19_c2_1 = p_19_1 << 1;
  assign t_r19_c2_2 = p_19_2 << 2;
  assign t_r19_c2_3 = p_19_3 << 1;
  assign t_r19_c2_4 = p_20_2 << 1;
  assign t_r19_c2_5 = t_r19_c2_0 + p_18_1;
  assign t_r19_c2_6 = t_r19_c2_1 + p_18_3;
  assign t_r19_c2_7 = t_r19_c2_2 + t_r19_c2_3;
  assign t_r19_c2_8 = t_r19_c2_4 + p_20_1;
  assign t_r19_c2_9 = t_r19_c2_5 + t_r19_c2_6;
  assign t_r19_c2_10 = t_r19_c2_7 + t_r19_c2_8;
  assign t_r19_c2_11 = t_r19_c2_9 + t_r19_c2_10;
  assign t_r19_c2_12 = t_r19_c2_11 + p_20_3;
  assign out_19_2 = t_r19_c2_12 >> 4;

  assign t_r19_c3_0 = p_18_3 << 1;
  assign t_r19_c3_1 = p_19_2 << 1;
  assign t_r19_c3_2 = p_19_3 << 2;
  assign t_r19_c3_3 = p_19_4 << 1;
  assign t_r19_c3_4 = p_20_3 << 1;
  assign t_r19_c3_5 = t_r19_c3_0 + p_18_2;
  assign t_r19_c3_6 = t_r19_c3_1 + p_18_4;
  assign t_r19_c3_7 = t_r19_c3_2 + t_r19_c3_3;
  assign t_r19_c3_8 = t_r19_c3_4 + p_20_2;
  assign t_r19_c3_9 = t_r19_c3_5 + t_r19_c3_6;
  assign t_r19_c3_10 = t_r19_c3_7 + t_r19_c3_8;
  assign t_r19_c3_11 = t_r19_c3_9 + t_r19_c3_10;
  assign t_r19_c3_12 = t_r19_c3_11 + p_20_4;
  assign out_19_3 = t_r19_c3_12 >> 4;

  assign t_r19_c4_0 = p_18_4 << 1;
  assign t_r19_c4_1 = p_19_3 << 1;
  assign t_r19_c4_2 = p_19_4 << 2;
  assign t_r19_c4_3 = p_19_5 << 1;
  assign t_r19_c4_4 = p_20_4 << 1;
  assign t_r19_c4_5 = t_r19_c4_0 + p_18_3;
  assign t_r19_c4_6 = t_r19_c4_1 + p_18_5;
  assign t_r19_c4_7 = t_r19_c4_2 + t_r19_c4_3;
  assign t_r19_c4_8 = t_r19_c4_4 + p_20_3;
  assign t_r19_c4_9 = t_r19_c4_5 + t_r19_c4_6;
  assign t_r19_c4_10 = t_r19_c4_7 + t_r19_c4_8;
  assign t_r19_c4_11 = t_r19_c4_9 + t_r19_c4_10;
  assign t_r19_c4_12 = t_r19_c4_11 + p_20_5;
  assign out_19_4 = t_r19_c4_12 >> 4;

  assign t_r19_c5_0 = p_18_5 << 1;
  assign t_r19_c5_1 = p_19_4 << 1;
  assign t_r19_c5_2 = p_19_5 << 2;
  assign t_r19_c5_3 = p_19_6 << 1;
  assign t_r19_c5_4 = p_20_5 << 1;
  assign t_r19_c5_5 = t_r19_c5_0 + p_18_4;
  assign t_r19_c5_6 = t_r19_c5_1 + p_18_6;
  assign t_r19_c5_7 = t_r19_c5_2 + t_r19_c5_3;
  assign t_r19_c5_8 = t_r19_c5_4 + p_20_4;
  assign t_r19_c5_9 = t_r19_c5_5 + t_r19_c5_6;
  assign t_r19_c5_10 = t_r19_c5_7 + t_r19_c5_8;
  assign t_r19_c5_11 = t_r19_c5_9 + t_r19_c5_10;
  assign t_r19_c5_12 = t_r19_c5_11 + p_20_6;
  assign out_19_5 = t_r19_c5_12 >> 4;

  assign t_r19_c6_0 = p_18_6 << 1;
  assign t_r19_c6_1 = p_19_5 << 1;
  assign t_r19_c6_2 = p_19_6 << 2;
  assign t_r19_c6_3 = p_19_7 << 1;
  assign t_r19_c6_4 = p_20_6 << 1;
  assign t_r19_c6_5 = t_r19_c6_0 + p_18_5;
  assign t_r19_c6_6 = t_r19_c6_1 + p_18_7;
  assign t_r19_c6_7 = t_r19_c6_2 + t_r19_c6_3;
  assign t_r19_c6_8 = t_r19_c6_4 + p_20_5;
  assign t_r19_c6_9 = t_r19_c6_5 + t_r19_c6_6;
  assign t_r19_c6_10 = t_r19_c6_7 + t_r19_c6_8;
  assign t_r19_c6_11 = t_r19_c6_9 + t_r19_c6_10;
  assign t_r19_c6_12 = t_r19_c6_11 + p_20_7;
  assign out_19_6 = t_r19_c6_12 >> 4;

  assign t_r19_c7_0 = p_18_7 << 1;
  assign t_r19_c7_1 = p_19_6 << 1;
  assign t_r19_c7_2 = p_19_7 << 2;
  assign t_r19_c7_3 = p_19_8 << 1;
  assign t_r19_c7_4 = p_20_7 << 1;
  assign t_r19_c7_5 = t_r19_c7_0 + p_18_6;
  assign t_r19_c7_6 = t_r19_c7_1 + p_18_8;
  assign t_r19_c7_7 = t_r19_c7_2 + t_r19_c7_3;
  assign t_r19_c7_8 = t_r19_c7_4 + p_20_6;
  assign t_r19_c7_9 = t_r19_c7_5 + t_r19_c7_6;
  assign t_r19_c7_10 = t_r19_c7_7 + t_r19_c7_8;
  assign t_r19_c7_11 = t_r19_c7_9 + t_r19_c7_10;
  assign t_r19_c7_12 = t_r19_c7_11 + p_20_8;
  assign out_19_7 = t_r19_c7_12 >> 4;

  assign t_r19_c8_0 = p_18_8 << 1;
  assign t_r19_c8_1 = p_19_7 << 1;
  assign t_r19_c8_2 = p_19_8 << 2;
  assign t_r19_c8_3 = p_19_9 << 1;
  assign t_r19_c8_4 = p_20_8 << 1;
  assign t_r19_c8_5 = t_r19_c8_0 + p_18_7;
  assign t_r19_c8_6 = t_r19_c8_1 + p_18_9;
  assign t_r19_c8_7 = t_r19_c8_2 + t_r19_c8_3;
  assign t_r19_c8_8 = t_r19_c8_4 + p_20_7;
  assign t_r19_c8_9 = t_r19_c8_5 + t_r19_c8_6;
  assign t_r19_c8_10 = t_r19_c8_7 + t_r19_c8_8;
  assign t_r19_c8_11 = t_r19_c8_9 + t_r19_c8_10;
  assign t_r19_c8_12 = t_r19_c8_11 + p_20_9;
  assign out_19_8 = t_r19_c8_12 >> 4;

  assign t_r19_c9_0 = p_18_9 << 1;
  assign t_r19_c9_1 = p_19_8 << 1;
  assign t_r19_c9_2 = p_19_9 << 2;
  assign t_r19_c9_3 = p_19_10 << 1;
  assign t_r19_c9_4 = p_20_9 << 1;
  assign t_r19_c9_5 = t_r19_c9_0 + p_18_8;
  assign t_r19_c9_6 = t_r19_c9_1 + p_18_10;
  assign t_r19_c9_7 = t_r19_c9_2 + t_r19_c9_3;
  assign t_r19_c9_8 = t_r19_c9_4 + p_20_8;
  assign t_r19_c9_9 = t_r19_c9_5 + t_r19_c9_6;
  assign t_r19_c9_10 = t_r19_c9_7 + t_r19_c9_8;
  assign t_r19_c9_11 = t_r19_c9_9 + t_r19_c9_10;
  assign t_r19_c9_12 = t_r19_c9_11 + p_20_10;
  assign out_19_9 = t_r19_c9_12 >> 4;

  assign t_r19_c10_0 = p_18_10 << 1;
  assign t_r19_c10_1 = p_19_9 << 1;
  assign t_r19_c10_2 = p_19_10 << 2;
  assign t_r19_c10_3 = p_19_11 << 1;
  assign t_r19_c10_4 = p_20_10 << 1;
  assign t_r19_c10_5 = t_r19_c10_0 + p_18_9;
  assign t_r19_c10_6 = t_r19_c10_1 + p_18_11;
  assign t_r19_c10_7 = t_r19_c10_2 + t_r19_c10_3;
  assign t_r19_c10_8 = t_r19_c10_4 + p_20_9;
  assign t_r19_c10_9 = t_r19_c10_5 + t_r19_c10_6;
  assign t_r19_c10_10 = t_r19_c10_7 + t_r19_c10_8;
  assign t_r19_c10_11 = t_r19_c10_9 + t_r19_c10_10;
  assign t_r19_c10_12 = t_r19_c10_11 + p_20_11;
  assign out_19_10 = t_r19_c10_12 >> 4;

  assign t_r19_c11_0 = p_18_11 << 1;
  assign t_r19_c11_1 = p_19_10 << 1;
  assign t_r19_c11_2 = p_19_11 << 2;
  assign t_r19_c11_3 = p_19_12 << 1;
  assign t_r19_c11_4 = p_20_11 << 1;
  assign t_r19_c11_5 = t_r19_c11_0 + p_18_10;
  assign t_r19_c11_6 = t_r19_c11_1 + p_18_12;
  assign t_r19_c11_7 = t_r19_c11_2 + t_r19_c11_3;
  assign t_r19_c11_8 = t_r19_c11_4 + p_20_10;
  assign t_r19_c11_9 = t_r19_c11_5 + t_r19_c11_6;
  assign t_r19_c11_10 = t_r19_c11_7 + t_r19_c11_8;
  assign t_r19_c11_11 = t_r19_c11_9 + t_r19_c11_10;
  assign t_r19_c11_12 = t_r19_c11_11 + p_20_12;
  assign out_19_11 = t_r19_c11_12 >> 4;

  assign t_r19_c12_0 = p_18_12 << 1;
  assign t_r19_c12_1 = p_19_11 << 1;
  assign t_r19_c12_2 = p_19_12 << 2;
  assign t_r19_c12_3 = p_19_13 << 1;
  assign t_r19_c12_4 = p_20_12 << 1;
  assign t_r19_c12_5 = t_r19_c12_0 + p_18_11;
  assign t_r19_c12_6 = t_r19_c12_1 + p_18_13;
  assign t_r19_c12_7 = t_r19_c12_2 + t_r19_c12_3;
  assign t_r19_c12_8 = t_r19_c12_4 + p_20_11;
  assign t_r19_c12_9 = t_r19_c12_5 + t_r19_c12_6;
  assign t_r19_c12_10 = t_r19_c12_7 + t_r19_c12_8;
  assign t_r19_c12_11 = t_r19_c12_9 + t_r19_c12_10;
  assign t_r19_c12_12 = t_r19_c12_11 + p_20_13;
  assign out_19_12 = t_r19_c12_12 >> 4;

  assign t_r19_c13_0 = p_18_13 << 1;
  assign t_r19_c13_1 = p_19_12 << 1;
  assign t_r19_c13_2 = p_19_13 << 2;
  assign t_r19_c13_3 = p_19_14 << 1;
  assign t_r19_c13_4 = p_20_13 << 1;
  assign t_r19_c13_5 = t_r19_c13_0 + p_18_12;
  assign t_r19_c13_6 = t_r19_c13_1 + p_18_14;
  assign t_r19_c13_7 = t_r19_c13_2 + t_r19_c13_3;
  assign t_r19_c13_8 = t_r19_c13_4 + p_20_12;
  assign t_r19_c13_9 = t_r19_c13_5 + t_r19_c13_6;
  assign t_r19_c13_10 = t_r19_c13_7 + t_r19_c13_8;
  assign t_r19_c13_11 = t_r19_c13_9 + t_r19_c13_10;
  assign t_r19_c13_12 = t_r19_c13_11 + p_20_14;
  assign out_19_13 = t_r19_c13_12 >> 4;

  assign t_r19_c14_0 = p_18_14 << 1;
  assign t_r19_c14_1 = p_19_13 << 1;
  assign t_r19_c14_2 = p_19_14 << 2;
  assign t_r19_c14_3 = p_19_15 << 1;
  assign t_r19_c14_4 = p_20_14 << 1;
  assign t_r19_c14_5 = t_r19_c14_0 + p_18_13;
  assign t_r19_c14_6 = t_r19_c14_1 + p_18_15;
  assign t_r19_c14_7 = t_r19_c14_2 + t_r19_c14_3;
  assign t_r19_c14_8 = t_r19_c14_4 + p_20_13;
  assign t_r19_c14_9 = t_r19_c14_5 + t_r19_c14_6;
  assign t_r19_c14_10 = t_r19_c14_7 + t_r19_c14_8;
  assign t_r19_c14_11 = t_r19_c14_9 + t_r19_c14_10;
  assign t_r19_c14_12 = t_r19_c14_11 + p_20_15;
  assign out_19_14 = t_r19_c14_12 >> 4;

  assign t_r19_c15_0 = p_18_15 << 1;
  assign t_r19_c15_1 = p_19_14 << 1;
  assign t_r19_c15_2 = p_19_15 << 2;
  assign t_r19_c15_3 = p_19_16 << 1;
  assign t_r19_c15_4 = p_20_15 << 1;
  assign t_r19_c15_5 = t_r19_c15_0 + p_18_14;
  assign t_r19_c15_6 = t_r19_c15_1 + p_18_16;
  assign t_r19_c15_7 = t_r19_c15_2 + t_r19_c15_3;
  assign t_r19_c15_8 = t_r19_c15_4 + p_20_14;
  assign t_r19_c15_9 = t_r19_c15_5 + t_r19_c15_6;
  assign t_r19_c15_10 = t_r19_c15_7 + t_r19_c15_8;
  assign t_r19_c15_11 = t_r19_c15_9 + t_r19_c15_10;
  assign t_r19_c15_12 = t_r19_c15_11 + p_20_16;
  assign out_19_15 = t_r19_c15_12 >> 4;

  assign t_r19_c16_0 = p_18_16 << 1;
  assign t_r19_c16_1 = p_19_15 << 1;
  assign t_r19_c16_2 = p_19_16 << 2;
  assign t_r19_c16_3 = p_19_17 << 1;
  assign t_r19_c16_4 = p_20_16 << 1;
  assign t_r19_c16_5 = t_r19_c16_0 + p_18_15;
  assign t_r19_c16_6 = t_r19_c16_1 + p_18_17;
  assign t_r19_c16_7 = t_r19_c16_2 + t_r19_c16_3;
  assign t_r19_c16_8 = t_r19_c16_4 + p_20_15;
  assign t_r19_c16_9 = t_r19_c16_5 + t_r19_c16_6;
  assign t_r19_c16_10 = t_r19_c16_7 + t_r19_c16_8;
  assign t_r19_c16_11 = t_r19_c16_9 + t_r19_c16_10;
  assign t_r19_c16_12 = t_r19_c16_11 + p_20_17;
  assign out_19_16 = t_r19_c16_12 >> 4;

  assign t_r19_c17_0 = p_18_17 << 1;
  assign t_r19_c17_1 = p_19_16 << 1;
  assign t_r19_c17_2 = p_19_17 << 2;
  assign t_r19_c17_3 = p_19_18 << 1;
  assign t_r19_c17_4 = p_20_17 << 1;
  assign t_r19_c17_5 = t_r19_c17_0 + p_18_16;
  assign t_r19_c17_6 = t_r19_c17_1 + p_18_18;
  assign t_r19_c17_7 = t_r19_c17_2 + t_r19_c17_3;
  assign t_r19_c17_8 = t_r19_c17_4 + p_20_16;
  assign t_r19_c17_9 = t_r19_c17_5 + t_r19_c17_6;
  assign t_r19_c17_10 = t_r19_c17_7 + t_r19_c17_8;
  assign t_r19_c17_11 = t_r19_c17_9 + t_r19_c17_10;
  assign t_r19_c17_12 = t_r19_c17_11 + p_20_18;
  assign out_19_17 = t_r19_c17_12 >> 4;

  assign t_r19_c18_0 = p_18_18 << 1;
  assign t_r19_c18_1 = p_19_17 << 1;
  assign t_r19_c18_2 = p_19_18 << 2;
  assign t_r19_c18_3 = p_19_19 << 1;
  assign t_r19_c18_4 = p_20_18 << 1;
  assign t_r19_c18_5 = t_r19_c18_0 + p_18_17;
  assign t_r19_c18_6 = t_r19_c18_1 + p_18_19;
  assign t_r19_c18_7 = t_r19_c18_2 + t_r19_c18_3;
  assign t_r19_c18_8 = t_r19_c18_4 + p_20_17;
  assign t_r19_c18_9 = t_r19_c18_5 + t_r19_c18_6;
  assign t_r19_c18_10 = t_r19_c18_7 + t_r19_c18_8;
  assign t_r19_c18_11 = t_r19_c18_9 + t_r19_c18_10;
  assign t_r19_c18_12 = t_r19_c18_11 + p_20_19;
  assign out_19_18 = t_r19_c18_12 >> 4;

  assign t_r19_c19_0 = p_18_19 << 1;
  assign t_r19_c19_1 = p_19_18 << 1;
  assign t_r19_c19_2 = p_19_19 << 2;
  assign t_r19_c19_3 = p_19_20 << 1;
  assign t_r19_c19_4 = p_20_19 << 1;
  assign t_r19_c19_5 = t_r19_c19_0 + p_18_18;
  assign t_r19_c19_6 = t_r19_c19_1 + p_18_20;
  assign t_r19_c19_7 = t_r19_c19_2 + t_r19_c19_3;
  assign t_r19_c19_8 = t_r19_c19_4 + p_20_18;
  assign t_r19_c19_9 = t_r19_c19_5 + t_r19_c19_6;
  assign t_r19_c19_10 = t_r19_c19_7 + t_r19_c19_8;
  assign t_r19_c19_11 = t_r19_c19_9 + t_r19_c19_10;
  assign t_r19_c19_12 = t_r19_c19_11 + p_20_20;
  assign out_19_19 = t_r19_c19_12 >> 4;

  assign t_r19_c20_0 = p_18_20 << 1;
  assign t_r19_c20_1 = p_19_19 << 1;
  assign t_r19_c20_2 = p_19_20 << 2;
  assign t_r19_c20_3 = p_19_21 << 1;
  assign t_r19_c20_4 = p_20_20 << 1;
  assign t_r19_c20_5 = t_r19_c20_0 + p_18_19;
  assign t_r19_c20_6 = t_r19_c20_1 + p_18_21;
  assign t_r19_c20_7 = t_r19_c20_2 + t_r19_c20_3;
  assign t_r19_c20_8 = t_r19_c20_4 + p_20_19;
  assign t_r19_c20_9 = t_r19_c20_5 + t_r19_c20_6;
  assign t_r19_c20_10 = t_r19_c20_7 + t_r19_c20_8;
  assign t_r19_c20_11 = t_r19_c20_9 + t_r19_c20_10;
  assign t_r19_c20_12 = t_r19_c20_11 + p_20_21;
  assign out_19_20 = t_r19_c20_12 >> 4;

  assign t_r19_c21_0 = p_18_21 << 1;
  assign t_r19_c21_1 = p_19_20 << 1;
  assign t_r19_c21_2 = p_19_21 << 2;
  assign t_r19_c21_3 = p_19_22 << 1;
  assign t_r19_c21_4 = p_20_21 << 1;
  assign t_r19_c21_5 = t_r19_c21_0 + p_18_20;
  assign t_r19_c21_6 = t_r19_c21_1 + p_18_22;
  assign t_r19_c21_7 = t_r19_c21_2 + t_r19_c21_3;
  assign t_r19_c21_8 = t_r19_c21_4 + p_20_20;
  assign t_r19_c21_9 = t_r19_c21_5 + t_r19_c21_6;
  assign t_r19_c21_10 = t_r19_c21_7 + t_r19_c21_8;
  assign t_r19_c21_11 = t_r19_c21_9 + t_r19_c21_10;
  assign t_r19_c21_12 = t_r19_c21_11 + p_20_22;
  assign out_19_21 = t_r19_c21_12 >> 4;

  assign t_r19_c22_0 = p_18_22 << 1;
  assign t_r19_c22_1 = p_19_21 << 1;
  assign t_r19_c22_2 = p_19_22 << 2;
  assign t_r19_c22_3 = p_19_23 << 1;
  assign t_r19_c22_4 = p_20_22 << 1;
  assign t_r19_c22_5 = t_r19_c22_0 + p_18_21;
  assign t_r19_c22_6 = t_r19_c22_1 + p_18_23;
  assign t_r19_c22_7 = t_r19_c22_2 + t_r19_c22_3;
  assign t_r19_c22_8 = t_r19_c22_4 + p_20_21;
  assign t_r19_c22_9 = t_r19_c22_5 + t_r19_c22_6;
  assign t_r19_c22_10 = t_r19_c22_7 + t_r19_c22_8;
  assign t_r19_c22_11 = t_r19_c22_9 + t_r19_c22_10;
  assign t_r19_c22_12 = t_r19_c22_11 + p_20_23;
  assign out_19_22 = t_r19_c22_12 >> 4;

  assign t_r19_c23_0 = p_18_23 << 1;
  assign t_r19_c23_1 = p_19_22 << 1;
  assign t_r19_c23_2 = p_19_23 << 2;
  assign t_r19_c23_3 = p_19_24 << 1;
  assign t_r19_c23_4 = p_20_23 << 1;
  assign t_r19_c23_5 = t_r19_c23_0 + p_18_22;
  assign t_r19_c23_6 = t_r19_c23_1 + p_18_24;
  assign t_r19_c23_7 = t_r19_c23_2 + t_r19_c23_3;
  assign t_r19_c23_8 = t_r19_c23_4 + p_20_22;
  assign t_r19_c23_9 = t_r19_c23_5 + t_r19_c23_6;
  assign t_r19_c23_10 = t_r19_c23_7 + t_r19_c23_8;
  assign t_r19_c23_11 = t_r19_c23_9 + t_r19_c23_10;
  assign t_r19_c23_12 = t_r19_c23_11 + p_20_24;
  assign out_19_23 = t_r19_c23_12 >> 4;

  assign t_r19_c24_0 = p_18_24 << 1;
  assign t_r19_c24_1 = p_19_23 << 1;
  assign t_r19_c24_2 = p_19_24 << 2;
  assign t_r19_c24_3 = p_19_25 << 1;
  assign t_r19_c24_4 = p_20_24 << 1;
  assign t_r19_c24_5 = t_r19_c24_0 + p_18_23;
  assign t_r19_c24_6 = t_r19_c24_1 + p_18_25;
  assign t_r19_c24_7 = t_r19_c24_2 + t_r19_c24_3;
  assign t_r19_c24_8 = t_r19_c24_4 + p_20_23;
  assign t_r19_c24_9 = t_r19_c24_5 + t_r19_c24_6;
  assign t_r19_c24_10 = t_r19_c24_7 + t_r19_c24_8;
  assign t_r19_c24_11 = t_r19_c24_9 + t_r19_c24_10;
  assign t_r19_c24_12 = t_r19_c24_11 + p_20_25;
  assign out_19_24 = t_r19_c24_12 >> 4;

  assign t_r19_c25_0 = p_18_25 << 1;
  assign t_r19_c25_1 = p_19_24 << 1;
  assign t_r19_c25_2 = p_19_25 << 2;
  assign t_r19_c25_3 = p_19_26 << 1;
  assign t_r19_c25_4 = p_20_25 << 1;
  assign t_r19_c25_5 = t_r19_c25_0 + p_18_24;
  assign t_r19_c25_6 = t_r19_c25_1 + p_18_26;
  assign t_r19_c25_7 = t_r19_c25_2 + t_r19_c25_3;
  assign t_r19_c25_8 = t_r19_c25_4 + p_20_24;
  assign t_r19_c25_9 = t_r19_c25_5 + t_r19_c25_6;
  assign t_r19_c25_10 = t_r19_c25_7 + t_r19_c25_8;
  assign t_r19_c25_11 = t_r19_c25_9 + t_r19_c25_10;
  assign t_r19_c25_12 = t_r19_c25_11 + p_20_26;
  assign out_19_25 = t_r19_c25_12 >> 4;

  assign t_r19_c26_0 = p_18_26 << 1;
  assign t_r19_c26_1 = p_19_25 << 1;
  assign t_r19_c26_2 = p_19_26 << 2;
  assign t_r19_c26_3 = p_19_27 << 1;
  assign t_r19_c26_4 = p_20_26 << 1;
  assign t_r19_c26_5 = t_r19_c26_0 + p_18_25;
  assign t_r19_c26_6 = t_r19_c26_1 + p_18_27;
  assign t_r19_c26_7 = t_r19_c26_2 + t_r19_c26_3;
  assign t_r19_c26_8 = t_r19_c26_4 + p_20_25;
  assign t_r19_c26_9 = t_r19_c26_5 + t_r19_c26_6;
  assign t_r19_c26_10 = t_r19_c26_7 + t_r19_c26_8;
  assign t_r19_c26_11 = t_r19_c26_9 + t_r19_c26_10;
  assign t_r19_c26_12 = t_r19_c26_11 + p_20_27;
  assign out_19_26 = t_r19_c26_12 >> 4;

  assign t_r19_c27_0 = p_18_27 << 1;
  assign t_r19_c27_1 = p_19_26 << 1;
  assign t_r19_c27_2 = p_19_27 << 2;
  assign t_r19_c27_3 = p_19_28 << 1;
  assign t_r19_c27_4 = p_20_27 << 1;
  assign t_r19_c27_5 = t_r19_c27_0 + p_18_26;
  assign t_r19_c27_6 = t_r19_c27_1 + p_18_28;
  assign t_r19_c27_7 = t_r19_c27_2 + t_r19_c27_3;
  assign t_r19_c27_8 = t_r19_c27_4 + p_20_26;
  assign t_r19_c27_9 = t_r19_c27_5 + t_r19_c27_6;
  assign t_r19_c27_10 = t_r19_c27_7 + t_r19_c27_8;
  assign t_r19_c27_11 = t_r19_c27_9 + t_r19_c27_10;
  assign t_r19_c27_12 = t_r19_c27_11 + p_20_28;
  assign out_19_27 = t_r19_c27_12 >> 4;

  assign t_r19_c28_0 = p_18_28 << 1;
  assign t_r19_c28_1 = p_19_27 << 1;
  assign t_r19_c28_2 = p_19_28 << 2;
  assign t_r19_c28_3 = p_19_29 << 1;
  assign t_r19_c28_4 = p_20_28 << 1;
  assign t_r19_c28_5 = t_r19_c28_0 + p_18_27;
  assign t_r19_c28_6 = t_r19_c28_1 + p_18_29;
  assign t_r19_c28_7 = t_r19_c28_2 + t_r19_c28_3;
  assign t_r19_c28_8 = t_r19_c28_4 + p_20_27;
  assign t_r19_c28_9 = t_r19_c28_5 + t_r19_c28_6;
  assign t_r19_c28_10 = t_r19_c28_7 + t_r19_c28_8;
  assign t_r19_c28_11 = t_r19_c28_9 + t_r19_c28_10;
  assign t_r19_c28_12 = t_r19_c28_11 + p_20_29;
  assign out_19_28 = t_r19_c28_12 >> 4;

  assign t_r19_c29_0 = p_18_29 << 1;
  assign t_r19_c29_1 = p_19_28 << 1;
  assign t_r19_c29_2 = p_19_29 << 2;
  assign t_r19_c29_3 = p_19_30 << 1;
  assign t_r19_c29_4 = p_20_29 << 1;
  assign t_r19_c29_5 = t_r19_c29_0 + p_18_28;
  assign t_r19_c29_6 = t_r19_c29_1 + p_18_30;
  assign t_r19_c29_7 = t_r19_c29_2 + t_r19_c29_3;
  assign t_r19_c29_8 = t_r19_c29_4 + p_20_28;
  assign t_r19_c29_9 = t_r19_c29_5 + t_r19_c29_6;
  assign t_r19_c29_10 = t_r19_c29_7 + t_r19_c29_8;
  assign t_r19_c29_11 = t_r19_c29_9 + t_r19_c29_10;
  assign t_r19_c29_12 = t_r19_c29_11 + p_20_30;
  assign out_19_29 = t_r19_c29_12 >> 4;

  assign t_r19_c30_0 = p_18_30 << 1;
  assign t_r19_c30_1 = p_19_29 << 1;
  assign t_r19_c30_2 = p_19_30 << 2;
  assign t_r19_c30_3 = p_19_31 << 1;
  assign t_r19_c30_4 = p_20_30 << 1;
  assign t_r19_c30_5 = t_r19_c30_0 + p_18_29;
  assign t_r19_c30_6 = t_r19_c30_1 + p_18_31;
  assign t_r19_c30_7 = t_r19_c30_2 + t_r19_c30_3;
  assign t_r19_c30_8 = t_r19_c30_4 + p_20_29;
  assign t_r19_c30_9 = t_r19_c30_5 + t_r19_c30_6;
  assign t_r19_c30_10 = t_r19_c30_7 + t_r19_c30_8;
  assign t_r19_c30_11 = t_r19_c30_9 + t_r19_c30_10;
  assign t_r19_c30_12 = t_r19_c30_11 + p_20_31;
  assign out_19_30 = t_r19_c30_12 >> 4;

  assign t_r19_c31_0 = p_18_31 << 1;
  assign t_r19_c31_1 = p_19_30 << 1;
  assign t_r19_c31_2 = p_19_31 << 2;
  assign t_r19_c31_3 = p_19_32 << 1;
  assign t_r19_c31_4 = p_20_31 << 1;
  assign t_r19_c31_5 = t_r19_c31_0 + p_18_30;
  assign t_r19_c31_6 = t_r19_c31_1 + p_18_32;
  assign t_r19_c31_7 = t_r19_c31_2 + t_r19_c31_3;
  assign t_r19_c31_8 = t_r19_c31_4 + p_20_30;
  assign t_r19_c31_9 = t_r19_c31_5 + t_r19_c31_6;
  assign t_r19_c31_10 = t_r19_c31_7 + t_r19_c31_8;
  assign t_r19_c31_11 = t_r19_c31_9 + t_r19_c31_10;
  assign t_r19_c31_12 = t_r19_c31_11 + p_20_32;
  assign out_19_31 = t_r19_c31_12 >> 4;

  assign t_r19_c32_0 = p_18_32 << 1;
  assign t_r19_c32_1 = p_19_31 << 1;
  assign t_r19_c32_2 = p_19_32 << 2;
  assign t_r19_c32_3 = p_19_33 << 1;
  assign t_r19_c32_4 = p_20_32 << 1;
  assign t_r19_c32_5 = t_r19_c32_0 + p_18_31;
  assign t_r19_c32_6 = t_r19_c32_1 + p_18_33;
  assign t_r19_c32_7 = t_r19_c32_2 + t_r19_c32_3;
  assign t_r19_c32_8 = t_r19_c32_4 + p_20_31;
  assign t_r19_c32_9 = t_r19_c32_5 + t_r19_c32_6;
  assign t_r19_c32_10 = t_r19_c32_7 + t_r19_c32_8;
  assign t_r19_c32_11 = t_r19_c32_9 + t_r19_c32_10;
  assign t_r19_c32_12 = t_r19_c32_11 + p_20_33;
  assign out_19_32 = t_r19_c32_12 >> 4;

  assign t_r19_c33_0 = p_18_33 << 1;
  assign t_r19_c33_1 = p_19_32 << 1;
  assign t_r19_c33_2 = p_19_33 << 2;
  assign t_r19_c33_3 = p_19_34 << 1;
  assign t_r19_c33_4 = p_20_33 << 1;
  assign t_r19_c33_5 = t_r19_c33_0 + p_18_32;
  assign t_r19_c33_6 = t_r19_c33_1 + p_18_34;
  assign t_r19_c33_7 = t_r19_c33_2 + t_r19_c33_3;
  assign t_r19_c33_8 = t_r19_c33_4 + p_20_32;
  assign t_r19_c33_9 = t_r19_c33_5 + t_r19_c33_6;
  assign t_r19_c33_10 = t_r19_c33_7 + t_r19_c33_8;
  assign t_r19_c33_11 = t_r19_c33_9 + t_r19_c33_10;
  assign t_r19_c33_12 = t_r19_c33_11 + p_20_34;
  assign out_19_33 = t_r19_c33_12 >> 4;

  assign t_r19_c34_0 = p_18_34 << 1;
  assign t_r19_c34_1 = p_19_33 << 1;
  assign t_r19_c34_2 = p_19_34 << 2;
  assign t_r19_c34_3 = p_19_35 << 1;
  assign t_r19_c34_4 = p_20_34 << 1;
  assign t_r19_c34_5 = t_r19_c34_0 + p_18_33;
  assign t_r19_c34_6 = t_r19_c34_1 + p_18_35;
  assign t_r19_c34_7 = t_r19_c34_2 + t_r19_c34_3;
  assign t_r19_c34_8 = t_r19_c34_4 + p_20_33;
  assign t_r19_c34_9 = t_r19_c34_5 + t_r19_c34_6;
  assign t_r19_c34_10 = t_r19_c34_7 + t_r19_c34_8;
  assign t_r19_c34_11 = t_r19_c34_9 + t_r19_c34_10;
  assign t_r19_c34_12 = t_r19_c34_11 + p_20_35;
  assign out_19_34 = t_r19_c34_12 >> 4;

  assign t_r19_c35_0 = p_18_35 << 1;
  assign t_r19_c35_1 = p_19_34 << 1;
  assign t_r19_c35_2 = p_19_35 << 2;
  assign t_r19_c35_3 = p_19_36 << 1;
  assign t_r19_c35_4 = p_20_35 << 1;
  assign t_r19_c35_5 = t_r19_c35_0 + p_18_34;
  assign t_r19_c35_6 = t_r19_c35_1 + p_18_36;
  assign t_r19_c35_7 = t_r19_c35_2 + t_r19_c35_3;
  assign t_r19_c35_8 = t_r19_c35_4 + p_20_34;
  assign t_r19_c35_9 = t_r19_c35_5 + t_r19_c35_6;
  assign t_r19_c35_10 = t_r19_c35_7 + t_r19_c35_8;
  assign t_r19_c35_11 = t_r19_c35_9 + t_r19_c35_10;
  assign t_r19_c35_12 = t_r19_c35_11 + p_20_36;
  assign out_19_35 = t_r19_c35_12 >> 4;

  assign t_r19_c36_0 = p_18_36 << 1;
  assign t_r19_c36_1 = p_19_35 << 1;
  assign t_r19_c36_2 = p_19_36 << 2;
  assign t_r19_c36_3 = p_19_37 << 1;
  assign t_r19_c36_4 = p_20_36 << 1;
  assign t_r19_c36_5 = t_r19_c36_0 + p_18_35;
  assign t_r19_c36_6 = t_r19_c36_1 + p_18_37;
  assign t_r19_c36_7 = t_r19_c36_2 + t_r19_c36_3;
  assign t_r19_c36_8 = t_r19_c36_4 + p_20_35;
  assign t_r19_c36_9 = t_r19_c36_5 + t_r19_c36_6;
  assign t_r19_c36_10 = t_r19_c36_7 + t_r19_c36_8;
  assign t_r19_c36_11 = t_r19_c36_9 + t_r19_c36_10;
  assign t_r19_c36_12 = t_r19_c36_11 + p_20_37;
  assign out_19_36 = t_r19_c36_12 >> 4;

  assign t_r19_c37_0 = p_18_37 << 1;
  assign t_r19_c37_1 = p_19_36 << 1;
  assign t_r19_c37_2 = p_19_37 << 2;
  assign t_r19_c37_3 = p_19_38 << 1;
  assign t_r19_c37_4 = p_20_37 << 1;
  assign t_r19_c37_5 = t_r19_c37_0 + p_18_36;
  assign t_r19_c37_6 = t_r19_c37_1 + p_18_38;
  assign t_r19_c37_7 = t_r19_c37_2 + t_r19_c37_3;
  assign t_r19_c37_8 = t_r19_c37_4 + p_20_36;
  assign t_r19_c37_9 = t_r19_c37_5 + t_r19_c37_6;
  assign t_r19_c37_10 = t_r19_c37_7 + t_r19_c37_8;
  assign t_r19_c37_11 = t_r19_c37_9 + t_r19_c37_10;
  assign t_r19_c37_12 = t_r19_c37_11 + p_20_38;
  assign out_19_37 = t_r19_c37_12 >> 4;

  assign t_r19_c38_0 = p_18_38 << 1;
  assign t_r19_c38_1 = p_19_37 << 1;
  assign t_r19_c38_2 = p_19_38 << 2;
  assign t_r19_c38_3 = p_19_39 << 1;
  assign t_r19_c38_4 = p_20_38 << 1;
  assign t_r19_c38_5 = t_r19_c38_0 + p_18_37;
  assign t_r19_c38_6 = t_r19_c38_1 + p_18_39;
  assign t_r19_c38_7 = t_r19_c38_2 + t_r19_c38_3;
  assign t_r19_c38_8 = t_r19_c38_4 + p_20_37;
  assign t_r19_c38_9 = t_r19_c38_5 + t_r19_c38_6;
  assign t_r19_c38_10 = t_r19_c38_7 + t_r19_c38_8;
  assign t_r19_c38_11 = t_r19_c38_9 + t_r19_c38_10;
  assign t_r19_c38_12 = t_r19_c38_11 + p_20_39;
  assign out_19_38 = t_r19_c38_12 >> 4;

  assign t_r19_c39_0 = p_18_39 << 1;
  assign t_r19_c39_1 = p_19_38 << 1;
  assign t_r19_c39_2 = p_19_39 << 2;
  assign t_r19_c39_3 = p_19_40 << 1;
  assign t_r19_c39_4 = p_20_39 << 1;
  assign t_r19_c39_5 = t_r19_c39_0 + p_18_38;
  assign t_r19_c39_6 = t_r19_c39_1 + p_18_40;
  assign t_r19_c39_7 = t_r19_c39_2 + t_r19_c39_3;
  assign t_r19_c39_8 = t_r19_c39_4 + p_20_38;
  assign t_r19_c39_9 = t_r19_c39_5 + t_r19_c39_6;
  assign t_r19_c39_10 = t_r19_c39_7 + t_r19_c39_8;
  assign t_r19_c39_11 = t_r19_c39_9 + t_r19_c39_10;
  assign t_r19_c39_12 = t_r19_c39_11 + p_20_40;
  assign out_19_39 = t_r19_c39_12 >> 4;

  assign t_r19_c40_0 = p_18_40 << 1;
  assign t_r19_c40_1 = p_19_39 << 1;
  assign t_r19_c40_2 = p_19_40 << 2;
  assign t_r19_c40_3 = p_19_41 << 1;
  assign t_r19_c40_4 = p_20_40 << 1;
  assign t_r19_c40_5 = t_r19_c40_0 + p_18_39;
  assign t_r19_c40_6 = t_r19_c40_1 + p_18_41;
  assign t_r19_c40_7 = t_r19_c40_2 + t_r19_c40_3;
  assign t_r19_c40_8 = t_r19_c40_4 + p_20_39;
  assign t_r19_c40_9 = t_r19_c40_5 + t_r19_c40_6;
  assign t_r19_c40_10 = t_r19_c40_7 + t_r19_c40_8;
  assign t_r19_c40_11 = t_r19_c40_9 + t_r19_c40_10;
  assign t_r19_c40_12 = t_r19_c40_11 + p_20_41;
  assign out_19_40 = t_r19_c40_12 >> 4;

  assign t_r19_c41_0 = p_18_41 << 1;
  assign t_r19_c41_1 = p_19_40 << 1;
  assign t_r19_c41_2 = p_19_41 << 2;
  assign t_r19_c41_3 = p_19_42 << 1;
  assign t_r19_c41_4 = p_20_41 << 1;
  assign t_r19_c41_5 = t_r19_c41_0 + p_18_40;
  assign t_r19_c41_6 = t_r19_c41_1 + p_18_42;
  assign t_r19_c41_7 = t_r19_c41_2 + t_r19_c41_3;
  assign t_r19_c41_8 = t_r19_c41_4 + p_20_40;
  assign t_r19_c41_9 = t_r19_c41_5 + t_r19_c41_6;
  assign t_r19_c41_10 = t_r19_c41_7 + t_r19_c41_8;
  assign t_r19_c41_11 = t_r19_c41_9 + t_r19_c41_10;
  assign t_r19_c41_12 = t_r19_c41_11 + p_20_42;
  assign out_19_41 = t_r19_c41_12 >> 4;

  assign t_r19_c42_0 = p_18_42 << 1;
  assign t_r19_c42_1 = p_19_41 << 1;
  assign t_r19_c42_2 = p_19_42 << 2;
  assign t_r19_c42_3 = p_19_43 << 1;
  assign t_r19_c42_4 = p_20_42 << 1;
  assign t_r19_c42_5 = t_r19_c42_0 + p_18_41;
  assign t_r19_c42_6 = t_r19_c42_1 + p_18_43;
  assign t_r19_c42_7 = t_r19_c42_2 + t_r19_c42_3;
  assign t_r19_c42_8 = t_r19_c42_4 + p_20_41;
  assign t_r19_c42_9 = t_r19_c42_5 + t_r19_c42_6;
  assign t_r19_c42_10 = t_r19_c42_7 + t_r19_c42_8;
  assign t_r19_c42_11 = t_r19_c42_9 + t_r19_c42_10;
  assign t_r19_c42_12 = t_r19_c42_11 + p_20_43;
  assign out_19_42 = t_r19_c42_12 >> 4;

  assign t_r19_c43_0 = p_18_43 << 1;
  assign t_r19_c43_1 = p_19_42 << 1;
  assign t_r19_c43_2 = p_19_43 << 2;
  assign t_r19_c43_3 = p_19_44 << 1;
  assign t_r19_c43_4 = p_20_43 << 1;
  assign t_r19_c43_5 = t_r19_c43_0 + p_18_42;
  assign t_r19_c43_6 = t_r19_c43_1 + p_18_44;
  assign t_r19_c43_7 = t_r19_c43_2 + t_r19_c43_3;
  assign t_r19_c43_8 = t_r19_c43_4 + p_20_42;
  assign t_r19_c43_9 = t_r19_c43_5 + t_r19_c43_6;
  assign t_r19_c43_10 = t_r19_c43_7 + t_r19_c43_8;
  assign t_r19_c43_11 = t_r19_c43_9 + t_r19_c43_10;
  assign t_r19_c43_12 = t_r19_c43_11 + p_20_44;
  assign out_19_43 = t_r19_c43_12 >> 4;

  assign t_r19_c44_0 = p_18_44 << 1;
  assign t_r19_c44_1 = p_19_43 << 1;
  assign t_r19_c44_2 = p_19_44 << 2;
  assign t_r19_c44_3 = p_19_45 << 1;
  assign t_r19_c44_4 = p_20_44 << 1;
  assign t_r19_c44_5 = t_r19_c44_0 + p_18_43;
  assign t_r19_c44_6 = t_r19_c44_1 + p_18_45;
  assign t_r19_c44_7 = t_r19_c44_2 + t_r19_c44_3;
  assign t_r19_c44_8 = t_r19_c44_4 + p_20_43;
  assign t_r19_c44_9 = t_r19_c44_5 + t_r19_c44_6;
  assign t_r19_c44_10 = t_r19_c44_7 + t_r19_c44_8;
  assign t_r19_c44_11 = t_r19_c44_9 + t_r19_c44_10;
  assign t_r19_c44_12 = t_r19_c44_11 + p_20_45;
  assign out_19_44 = t_r19_c44_12 >> 4;

  assign t_r19_c45_0 = p_18_45 << 1;
  assign t_r19_c45_1 = p_19_44 << 1;
  assign t_r19_c45_2 = p_19_45 << 2;
  assign t_r19_c45_3 = p_19_46 << 1;
  assign t_r19_c45_4 = p_20_45 << 1;
  assign t_r19_c45_5 = t_r19_c45_0 + p_18_44;
  assign t_r19_c45_6 = t_r19_c45_1 + p_18_46;
  assign t_r19_c45_7 = t_r19_c45_2 + t_r19_c45_3;
  assign t_r19_c45_8 = t_r19_c45_4 + p_20_44;
  assign t_r19_c45_9 = t_r19_c45_5 + t_r19_c45_6;
  assign t_r19_c45_10 = t_r19_c45_7 + t_r19_c45_8;
  assign t_r19_c45_11 = t_r19_c45_9 + t_r19_c45_10;
  assign t_r19_c45_12 = t_r19_c45_11 + p_20_46;
  assign out_19_45 = t_r19_c45_12 >> 4;

  assign t_r19_c46_0 = p_18_46 << 1;
  assign t_r19_c46_1 = p_19_45 << 1;
  assign t_r19_c46_2 = p_19_46 << 2;
  assign t_r19_c46_3 = p_19_47 << 1;
  assign t_r19_c46_4 = p_20_46 << 1;
  assign t_r19_c46_5 = t_r19_c46_0 + p_18_45;
  assign t_r19_c46_6 = t_r19_c46_1 + p_18_47;
  assign t_r19_c46_7 = t_r19_c46_2 + t_r19_c46_3;
  assign t_r19_c46_8 = t_r19_c46_4 + p_20_45;
  assign t_r19_c46_9 = t_r19_c46_5 + t_r19_c46_6;
  assign t_r19_c46_10 = t_r19_c46_7 + t_r19_c46_8;
  assign t_r19_c46_11 = t_r19_c46_9 + t_r19_c46_10;
  assign t_r19_c46_12 = t_r19_c46_11 + p_20_47;
  assign out_19_46 = t_r19_c46_12 >> 4;

  assign t_r19_c47_0 = p_18_47 << 1;
  assign t_r19_c47_1 = p_19_46 << 1;
  assign t_r19_c47_2 = p_19_47 << 2;
  assign t_r19_c47_3 = p_19_48 << 1;
  assign t_r19_c47_4 = p_20_47 << 1;
  assign t_r19_c47_5 = t_r19_c47_0 + p_18_46;
  assign t_r19_c47_6 = t_r19_c47_1 + p_18_48;
  assign t_r19_c47_7 = t_r19_c47_2 + t_r19_c47_3;
  assign t_r19_c47_8 = t_r19_c47_4 + p_20_46;
  assign t_r19_c47_9 = t_r19_c47_5 + t_r19_c47_6;
  assign t_r19_c47_10 = t_r19_c47_7 + t_r19_c47_8;
  assign t_r19_c47_11 = t_r19_c47_9 + t_r19_c47_10;
  assign t_r19_c47_12 = t_r19_c47_11 + p_20_48;
  assign out_19_47 = t_r19_c47_12 >> 4;

  assign t_r19_c48_0 = p_18_48 << 1;
  assign t_r19_c48_1 = p_19_47 << 1;
  assign t_r19_c48_2 = p_19_48 << 2;
  assign t_r19_c48_3 = p_19_49 << 1;
  assign t_r19_c48_4 = p_20_48 << 1;
  assign t_r19_c48_5 = t_r19_c48_0 + p_18_47;
  assign t_r19_c48_6 = t_r19_c48_1 + p_18_49;
  assign t_r19_c48_7 = t_r19_c48_2 + t_r19_c48_3;
  assign t_r19_c48_8 = t_r19_c48_4 + p_20_47;
  assign t_r19_c48_9 = t_r19_c48_5 + t_r19_c48_6;
  assign t_r19_c48_10 = t_r19_c48_7 + t_r19_c48_8;
  assign t_r19_c48_11 = t_r19_c48_9 + t_r19_c48_10;
  assign t_r19_c48_12 = t_r19_c48_11 + p_20_49;
  assign out_19_48 = t_r19_c48_12 >> 4;

  assign t_r19_c49_0 = p_18_49 << 1;
  assign t_r19_c49_1 = p_19_48 << 1;
  assign t_r19_c49_2 = p_19_49 << 2;
  assign t_r19_c49_3 = p_19_50 << 1;
  assign t_r19_c49_4 = p_20_49 << 1;
  assign t_r19_c49_5 = t_r19_c49_0 + p_18_48;
  assign t_r19_c49_6 = t_r19_c49_1 + p_18_50;
  assign t_r19_c49_7 = t_r19_c49_2 + t_r19_c49_3;
  assign t_r19_c49_8 = t_r19_c49_4 + p_20_48;
  assign t_r19_c49_9 = t_r19_c49_5 + t_r19_c49_6;
  assign t_r19_c49_10 = t_r19_c49_7 + t_r19_c49_8;
  assign t_r19_c49_11 = t_r19_c49_9 + t_r19_c49_10;
  assign t_r19_c49_12 = t_r19_c49_11 + p_20_50;
  assign out_19_49 = t_r19_c49_12 >> 4;

  assign t_r19_c50_0 = p_18_50 << 1;
  assign t_r19_c50_1 = p_19_49 << 1;
  assign t_r19_c50_2 = p_19_50 << 2;
  assign t_r19_c50_3 = p_19_51 << 1;
  assign t_r19_c50_4 = p_20_50 << 1;
  assign t_r19_c50_5 = t_r19_c50_0 + p_18_49;
  assign t_r19_c50_6 = t_r19_c50_1 + p_18_51;
  assign t_r19_c50_7 = t_r19_c50_2 + t_r19_c50_3;
  assign t_r19_c50_8 = t_r19_c50_4 + p_20_49;
  assign t_r19_c50_9 = t_r19_c50_5 + t_r19_c50_6;
  assign t_r19_c50_10 = t_r19_c50_7 + t_r19_c50_8;
  assign t_r19_c50_11 = t_r19_c50_9 + t_r19_c50_10;
  assign t_r19_c50_12 = t_r19_c50_11 + p_20_51;
  assign out_19_50 = t_r19_c50_12 >> 4;

  assign t_r19_c51_0 = p_18_51 << 1;
  assign t_r19_c51_1 = p_19_50 << 1;
  assign t_r19_c51_2 = p_19_51 << 2;
  assign t_r19_c51_3 = p_19_52 << 1;
  assign t_r19_c51_4 = p_20_51 << 1;
  assign t_r19_c51_5 = t_r19_c51_0 + p_18_50;
  assign t_r19_c51_6 = t_r19_c51_1 + p_18_52;
  assign t_r19_c51_7 = t_r19_c51_2 + t_r19_c51_3;
  assign t_r19_c51_8 = t_r19_c51_4 + p_20_50;
  assign t_r19_c51_9 = t_r19_c51_5 + t_r19_c51_6;
  assign t_r19_c51_10 = t_r19_c51_7 + t_r19_c51_8;
  assign t_r19_c51_11 = t_r19_c51_9 + t_r19_c51_10;
  assign t_r19_c51_12 = t_r19_c51_11 + p_20_52;
  assign out_19_51 = t_r19_c51_12 >> 4;

  assign t_r19_c52_0 = p_18_52 << 1;
  assign t_r19_c52_1 = p_19_51 << 1;
  assign t_r19_c52_2 = p_19_52 << 2;
  assign t_r19_c52_3 = p_19_53 << 1;
  assign t_r19_c52_4 = p_20_52 << 1;
  assign t_r19_c52_5 = t_r19_c52_0 + p_18_51;
  assign t_r19_c52_6 = t_r19_c52_1 + p_18_53;
  assign t_r19_c52_7 = t_r19_c52_2 + t_r19_c52_3;
  assign t_r19_c52_8 = t_r19_c52_4 + p_20_51;
  assign t_r19_c52_9 = t_r19_c52_5 + t_r19_c52_6;
  assign t_r19_c52_10 = t_r19_c52_7 + t_r19_c52_8;
  assign t_r19_c52_11 = t_r19_c52_9 + t_r19_c52_10;
  assign t_r19_c52_12 = t_r19_c52_11 + p_20_53;
  assign out_19_52 = t_r19_c52_12 >> 4;

  assign t_r19_c53_0 = p_18_53 << 1;
  assign t_r19_c53_1 = p_19_52 << 1;
  assign t_r19_c53_2 = p_19_53 << 2;
  assign t_r19_c53_3 = p_19_54 << 1;
  assign t_r19_c53_4 = p_20_53 << 1;
  assign t_r19_c53_5 = t_r19_c53_0 + p_18_52;
  assign t_r19_c53_6 = t_r19_c53_1 + p_18_54;
  assign t_r19_c53_7 = t_r19_c53_2 + t_r19_c53_3;
  assign t_r19_c53_8 = t_r19_c53_4 + p_20_52;
  assign t_r19_c53_9 = t_r19_c53_5 + t_r19_c53_6;
  assign t_r19_c53_10 = t_r19_c53_7 + t_r19_c53_8;
  assign t_r19_c53_11 = t_r19_c53_9 + t_r19_c53_10;
  assign t_r19_c53_12 = t_r19_c53_11 + p_20_54;
  assign out_19_53 = t_r19_c53_12 >> 4;

  assign t_r19_c54_0 = p_18_54 << 1;
  assign t_r19_c54_1 = p_19_53 << 1;
  assign t_r19_c54_2 = p_19_54 << 2;
  assign t_r19_c54_3 = p_19_55 << 1;
  assign t_r19_c54_4 = p_20_54 << 1;
  assign t_r19_c54_5 = t_r19_c54_0 + p_18_53;
  assign t_r19_c54_6 = t_r19_c54_1 + p_18_55;
  assign t_r19_c54_7 = t_r19_c54_2 + t_r19_c54_3;
  assign t_r19_c54_8 = t_r19_c54_4 + p_20_53;
  assign t_r19_c54_9 = t_r19_c54_5 + t_r19_c54_6;
  assign t_r19_c54_10 = t_r19_c54_7 + t_r19_c54_8;
  assign t_r19_c54_11 = t_r19_c54_9 + t_r19_c54_10;
  assign t_r19_c54_12 = t_r19_c54_11 + p_20_55;
  assign out_19_54 = t_r19_c54_12 >> 4;

  assign t_r19_c55_0 = p_18_55 << 1;
  assign t_r19_c55_1 = p_19_54 << 1;
  assign t_r19_c55_2 = p_19_55 << 2;
  assign t_r19_c55_3 = p_19_56 << 1;
  assign t_r19_c55_4 = p_20_55 << 1;
  assign t_r19_c55_5 = t_r19_c55_0 + p_18_54;
  assign t_r19_c55_6 = t_r19_c55_1 + p_18_56;
  assign t_r19_c55_7 = t_r19_c55_2 + t_r19_c55_3;
  assign t_r19_c55_8 = t_r19_c55_4 + p_20_54;
  assign t_r19_c55_9 = t_r19_c55_5 + t_r19_c55_6;
  assign t_r19_c55_10 = t_r19_c55_7 + t_r19_c55_8;
  assign t_r19_c55_11 = t_r19_c55_9 + t_r19_c55_10;
  assign t_r19_c55_12 = t_r19_c55_11 + p_20_56;
  assign out_19_55 = t_r19_c55_12 >> 4;

  assign t_r19_c56_0 = p_18_56 << 1;
  assign t_r19_c56_1 = p_19_55 << 1;
  assign t_r19_c56_2 = p_19_56 << 2;
  assign t_r19_c56_3 = p_19_57 << 1;
  assign t_r19_c56_4 = p_20_56 << 1;
  assign t_r19_c56_5 = t_r19_c56_0 + p_18_55;
  assign t_r19_c56_6 = t_r19_c56_1 + p_18_57;
  assign t_r19_c56_7 = t_r19_c56_2 + t_r19_c56_3;
  assign t_r19_c56_8 = t_r19_c56_4 + p_20_55;
  assign t_r19_c56_9 = t_r19_c56_5 + t_r19_c56_6;
  assign t_r19_c56_10 = t_r19_c56_7 + t_r19_c56_8;
  assign t_r19_c56_11 = t_r19_c56_9 + t_r19_c56_10;
  assign t_r19_c56_12 = t_r19_c56_11 + p_20_57;
  assign out_19_56 = t_r19_c56_12 >> 4;

  assign t_r19_c57_0 = p_18_57 << 1;
  assign t_r19_c57_1 = p_19_56 << 1;
  assign t_r19_c57_2 = p_19_57 << 2;
  assign t_r19_c57_3 = p_19_58 << 1;
  assign t_r19_c57_4 = p_20_57 << 1;
  assign t_r19_c57_5 = t_r19_c57_0 + p_18_56;
  assign t_r19_c57_6 = t_r19_c57_1 + p_18_58;
  assign t_r19_c57_7 = t_r19_c57_2 + t_r19_c57_3;
  assign t_r19_c57_8 = t_r19_c57_4 + p_20_56;
  assign t_r19_c57_9 = t_r19_c57_5 + t_r19_c57_6;
  assign t_r19_c57_10 = t_r19_c57_7 + t_r19_c57_8;
  assign t_r19_c57_11 = t_r19_c57_9 + t_r19_c57_10;
  assign t_r19_c57_12 = t_r19_c57_11 + p_20_58;
  assign out_19_57 = t_r19_c57_12 >> 4;

  assign t_r19_c58_0 = p_18_58 << 1;
  assign t_r19_c58_1 = p_19_57 << 1;
  assign t_r19_c58_2 = p_19_58 << 2;
  assign t_r19_c58_3 = p_19_59 << 1;
  assign t_r19_c58_4 = p_20_58 << 1;
  assign t_r19_c58_5 = t_r19_c58_0 + p_18_57;
  assign t_r19_c58_6 = t_r19_c58_1 + p_18_59;
  assign t_r19_c58_7 = t_r19_c58_2 + t_r19_c58_3;
  assign t_r19_c58_8 = t_r19_c58_4 + p_20_57;
  assign t_r19_c58_9 = t_r19_c58_5 + t_r19_c58_6;
  assign t_r19_c58_10 = t_r19_c58_7 + t_r19_c58_8;
  assign t_r19_c58_11 = t_r19_c58_9 + t_r19_c58_10;
  assign t_r19_c58_12 = t_r19_c58_11 + p_20_59;
  assign out_19_58 = t_r19_c58_12 >> 4;

  assign t_r19_c59_0 = p_18_59 << 1;
  assign t_r19_c59_1 = p_19_58 << 1;
  assign t_r19_c59_2 = p_19_59 << 2;
  assign t_r19_c59_3 = p_19_60 << 1;
  assign t_r19_c59_4 = p_20_59 << 1;
  assign t_r19_c59_5 = t_r19_c59_0 + p_18_58;
  assign t_r19_c59_6 = t_r19_c59_1 + p_18_60;
  assign t_r19_c59_7 = t_r19_c59_2 + t_r19_c59_3;
  assign t_r19_c59_8 = t_r19_c59_4 + p_20_58;
  assign t_r19_c59_9 = t_r19_c59_5 + t_r19_c59_6;
  assign t_r19_c59_10 = t_r19_c59_7 + t_r19_c59_8;
  assign t_r19_c59_11 = t_r19_c59_9 + t_r19_c59_10;
  assign t_r19_c59_12 = t_r19_c59_11 + p_20_60;
  assign out_19_59 = t_r19_c59_12 >> 4;

  assign t_r19_c60_0 = p_18_60 << 1;
  assign t_r19_c60_1 = p_19_59 << 1;
  assign t_r19_c60_2 = p_19_60 << 2;
  assign t_r19_c60_3 = p_19_61 << 1;
  assign t_r19_c60_4 = p_20_60 << 1;
  assign t_r19_c60_5 = t_r19_c60_0 + p_18_59;
  assign t_r19_c60_6 = t_r19_c60_1 + p_18_61;
  assign t_r19_c60_7 = t_r19_c60_2 + t_r19_c60_3;
  assign t_r19_c60_8 = t_r19_c60_4 + p_20_59;
  assign t_r19_c60_9 = t_r19_c60_5 + t_r19_c60_6;
  assign t_r19_c60_10 = t_r19_c60_7 + t_r19_c60_8;
  assign t_r19_c60_11 = t_r19_c60_9 + t_r19_c60_10;
  assign t_r19_c60_12 = t_r19_c60_11 + p_20_61;
  assign out_19_60 = t_r19_c60_12 >> 4;

  assign t_r19_c61_0 = p_18_61 << 1;
  assign t_r19_c61_1 = p_19_60 << 1;
  assign t_r19_c61_2 = p_19_61 << 2;
  assign t_r19_c61_3 = p_19_62 << 1;
  assign t_r19_c61_4 = p_20_61 << 1;
  assign t_r19_c61_5 = t_r19_c61_0 + p_18_60;
  assign t_r19_c61_6 = t_r19_c61_1 + p_18_62;
  assign t_r19_c61_7 = t_r19_c61_2 + t_r19_c61_3;
  assign t_r19_c61_8 = t_r19_c61_4 + p_20_60;
  assign t_r19_c61_9 = t_r19_c61_5 + t_r19_c61_6;
  assign t_r19_c61_10 = t_r19_c61_7 + t_r19_c61_8;
  assign t_r19_c61_11 = t_r19_c61_9 + t_r19_c61_10;
  assign t_r19_c61_12 = t_r19_c61_11 + p_20_62;
  assign out_19_61 = t_r19_c61_12 >> 4;

  assign t_r19_c62_0 = p_18_62 << 1;
  assign t_r19_c62_1 = p_19_61 << 1;
  assign t_r19_c62_2 = p_19_62 << 2;
  assign t_r19_c62_3 = p_19_63 << 1;
  assign t_r19_c62_4 = p_20_62 << 1;
  assign t_r19_c62_5 = t_r19_c62_0 + p_18_61;
  assign t_r19_c62_6 = t_r19_c62_1 + p_18_63;
  assign t_r19_c62_7 = t_r19_c62_2 + t_r19_c62_3;
  assign t_r19_c62_8 = t_r19_c62_4 + p_20_61;
  assign t_r19_c62_9 = t_r19_c62_5 + t_r19_c62_6;
  assign t_r19_c62_10 = t_r19_c62_7 + t_r19_c62_8;
  assign t_r19_c62_11 = t_r19_c62_9 + t_r19_c62_10;
  assign t_r19_c62_12 = t_r19_c62_11 + p_20_63;
  assign out_19_62 = t_r19_c62_12 >> 4;

  assign t_r19_c63_0 = p_18_63 << 1;
  assign t_r19_c63_1 = p_19_62 << 1;
  assign t_r19_c63_2 = p_19_63 << 2;
  assign t_r19_c63_3 = p_19_64 << 1;
  assign t_r19_c63_4 = p_20_63 << 1;
  assign t_r19_c63_5 = t_r19_c63_0 + p_18_62;
  assign t_r19_c63_6 = t_r19_c63_1 + p_18_64;
  assign t_r19_c63_7 = t_r19_c63_2 + t_r19_c63_3;
  assign t_r19_c63_8 = t_r19_c63_4 + p_20_62;
  assign t_r19_c63_9 = t_r19_c63_5 + t_r19_c63_6;
  assign t_r19_c63_10 = t_r19_c63_7 + t_r19_c63_8;
  assign t_r19_c63_11 = t_r19_c63_9 + t_r19_c63_10;
  assign t_r19_c63_12 = t_r19_c63_11 + p_20_64;
  assign out_19_63 = t_r19_c63_12 >> 4;

  assign t_r19_c64_0 = p_18_64 << 1;
  assign t_r19_c64_1 = p_19_63 << 1;
  assign t_r19_c64_2 = p_19_64 << 2;
  assign t_r19_c64_3 = p_19_65 << 1;
  assign t_r19_c64_4 = p_20_64 << 1;
  assign t_r19_c64_5 = t_r19_c64_0 + p_18_63;
  assign t_r19_c64_6 = t_r19_c64_1 + p_18_65;
  assign t_r19_c64_7 = t_r19_c64_2 + t_r19_c64_3;
  assign t_r19_c64_8 = t_r19_c64_4 + p_20_63;
  assign t_r19_c64_9 = t_r19_c64_5 + t_r19_c64_6;
  assign t_r19_c64_10 = t_r19_c64_7 + t_r19_c64_8;
  assign t_r19_c64_11 = t_r19_c64_9 + t_r19_c64_10;
  assign t_r19_c64_12 = t_r19_c64_11 + p_20_65;
  assign out_19_64 = t_r19_c64_12 >> 4;

  assign t_r20_c1_0 = p_19_1 << 1;
  assign t_r20_c1_1 = p_20_0 << 1;
  assign t_r20_c1_2 = p_20_1 << 2;
  assign t_r20_c1_3 = p_20_2 << 1;
  assign t_r20_c1_4 = p_21_1 << 1;
  assign t_r20_c1_5 = t_r20_c1_0 + p_19_0;
  assign t_r20_c1_6 = t_r20_c1_1 + p_19_2;
  assign t_r20_c1_7 = t_r20_c1_2 + t_r20_c1_3;
  assign t_r20_c1_8 = t_r20_c1_4 + p_21_0;
  assign t_r20_c1_9 = t_r20_c1_5 + t_r20_c1_6;
  assign t_r20_c1_10 = t_r20_c1_7 + t_r20_c1_8;
  assign t_r20_c1_11 = t_r20_c1_9 + t_r20_c1_10;
  assign t_r20_c1_12 = t_r20_c1_11 + p_21_2;
  assign out_20_1 = t_r20_c1_12 >> 4;

  assign t_r20_c2_0 = p_19_2 << 1;
  assign t_r20_c2_1 = p_20_1 << 1;
  assign t_r20_c2_2 = p_20_2 << 2;
  assign t_r20_c2_3 = p_20_3 << 1;
  assign t_r20_c2_4 = p_21_2 << 1;
  assign t_r20_c2_5 = t_r20_c2_0 + p_19_1;
  assign t_r20_c2_6 = t_r20_c2_1 + p_19_3;
  assign t_r20_c2_7 = t_r20_c2_2 + t_r20_c2_3;
  assign t_r20_c2_8 = t_r20_c2_4 + p_21_1;
  assign t_r20_c2_9 = t_r20_c2_5 + t_r20_c2_6;
  assign t_r20_c2_10 = t_r20_c2_7 + t_r20_c2_8;
  assign t_r20_c2_11 = t_r20_c2_9 + t_r20_c2_10;
  assign t_r20_c2_12 = t_r20_c2_11 + p_21_3;
  assign out_20_2 = t_r20_c2_12 >> 4;

  assign t_r20_c3_0 = p_19_3 << 1;
  assign t_r20_c3_1 = p_20_2 << 1;
  assign t_r20_c3_2 = p_20_3 << 2;
  assign t_r20_c3_3 = p_20_4 << 1;
  assign t_r20_c3_4 = p_21_3 << 1;
  assign t_r20_c3_5 = t_r20_c3_0 + p_19_2;
  assign t_r20_c3_6 = t_r20_c3_1 + p_19_4;
  assign t_r20_c3_7 = t_r20_c3_2 + t_r20_c3_3;
  assign t_r20_c3_8 = t_r20_c3_4 + p_21_2;
  assign t_r20_c3_9 = t_r20_c3_5 + t_r20_c3_6;
  assign t_r20_c3_10 = t_r20_c3_7 + t_r20_c3_8;
  assign t_r20_c3_11 = t_r20_c3_9 + t_r20_c3_10;
  assign t_r20_c3_12 = t_r20_c3_11 + p_21_4;
  assign out_20_3 = t_r20_c3_12 >> 4;

  assign t_r20_c4_0 = p_19_4 << 1;
  assign t_r20_c4_1 = p_20_3 << 1;
  assign t_r20_c4_2 = p_20_4 << 2;
  assign t_r20_c4_3 = p_20_5 << 1;
  assign t_r20_c4_4 = p_21_4 << 1;
  assign t_r20_c4_5 = t_r20_c4_0 + p_19_3;
  assign t_r20_c4_6 = t_r20_c4_1 + p_19_5;
  assign t_r20_c4_7 = t_r20_c4_2 + t_r20_c4_3;
  assign t_r20_c4_8 = t_r20_c4_4 + p_21_3;
  assign t_r20_c4_9 = t_r20_c4_5 + t_r20_c4_6;
  assign t_r20_c4_10 = t_r20_c4_7 + t_r20_c4_8;
  assign t_r20_c4_11 = t_r20_c4_9 + t_r20_c4_10;
  assign t_r20_c4_12 = t_r20_c4_11 + p_21_5;
  assign out_20_4 = t_r20_c4_12 >> 4;

  assign t_r20_c5_0 = p_19_5 << 1;
  assign t_r20_c5_1 = p_20_4 << 1;
  assign t_r20_c5_2 = p_20_5 << 2;
  assign t_r20_c5_3 = p_20_6 << 1;
  assign t_r20_c5_4 = p_21_5 << 1;
  assign t_r20_c5_5 = t_r20_c5_0 + p_19_4;
  assign t_r20_c5_6 = t_r20_c5_1 + p_19_6;
  assign t_r20_c5_7 = t_r20_c5_2 + t_r20_c5_3;
  assign t_r20_c5_8 = t_r20_c5_4 + p_21_4;
  assign t_r20_c5_9 = t_r20_c5_5 + t_r20_c5_6;
  assign t_r20_c5_10 = t_r20_c5_7 + t_r20_c5_8;
  assign t_r20_c5_11 = t_r20_c5_9 + t_r20_c5_10;
  assign t_r20_c5_12 = t_r20_c5_11 + p_21_6;
  assign out_20_5 = t_r20_c5_12 >> 4;

  assign t_r20_c6_0 = p_19_6 << 1;
  assign t_r20_c6_1 = p_20_5 << 1;
  assign t_r20_c6_2 = p_20_6 << 2;
  assign t_r20_c6_3 = p_20_7 << 1;
  assign t_r20_c6_4 = p_21_6 << 1;
  assign t_r20_c6_5 = t_r20_c6_0 + p_19_5;
  assign t_r20_c6_6 = t_r20_c6_1 + p_19_7;
  assign t_r20_c6_7 = t_r20_c6_2 + t_r20_c6_3;
  assign t_r20_c6_8 = t_r20_c6_4 + p_21_5;
  assign t_r20_c6_9 = t_r20_c6_5 + t_r20_c6_6;
  assign t_r20_c6_10 = t_r20_c6_7 + t_r20_c6_8;
  assign t_r20_c6_11 = t_r20_c6_9 + t_r20_c6_10;
  assign t_r20_c6_12 = t_r20_c6_11 + p_21_7;
  assign out_20_6 = t_r20_c6_12 >> 4;

  assign t_r20_c7_0 = p_19_7 << 1;
  assign t_r20_c7_1 = p_20_6 << 1;
  assign t_r20_c7_2 = p_20_7 << 2;
  assign t_r20_c7_3 = p_20_8 << 1;
  assign t_r20_c7_4 = p_21_7 << 1;
  assign t_r20_c7_5 = t_r20_c7_0 + p_19_6;
  assign t_r20_c7_6 = t_r20_c7_1 + p_19_8;
  assign t_r20_c7_7 = t_r20_c7_2 + t_r20_c7_3;
  assign t_r20_c7_8 = t_r20_c7_4 + p_21_6;
  assign t_r20_c7_9 = t_r20_c7_5 + t_r20_c7_6;
  assign t_r20_c7_10 = t_r20_c7_7 + t_r20_c7_8;
  assign t_r20_c7_11 = t_r20_c7_9 + t_r20_c7_10;
  assign t_r20_c7_12 = t_r20_c7_11 + p_21_8;
  assign out_20_7 = t_r20_c7_12 >> 4;

  assign t_r20_c8_0 = p_19_8 << 1;
  assign t_r20_c8_1 = p_20_7 << 1;
  assign t_r20_c8_2 = p_20_8 << 2;
  assign t_r20_c8_3 = p_20_9 << 1;
  assign t_r20_c8_4 = p_21_8 << 1;
  assign t_r20_c8_5 = t_r20_c8_0 + p_19_7;
  assign t_r20_c8_6 = t_r20_c8_1 + p_19_9;
  assign t_r20_c8_7 = t_r20_c8_2 + t_r20_c8_3;
  assign t_r20_c8_8 = t_r20_c8_4 + p_21_7;
  assign t_r20_c8_9 = t_r20_c8_5 + t_r20_c8_6;
  assign t_r20_c8_10 = t_r20_c8_7 + t_r20_c8_8;
  assign t_r20_c8_11 = t_r20_c8_9 + t_r20_c8_10;
  assign t_r20_c8_12 = t_r20_c8_11 + p_21_9;
  assign out_20_8 = t_r20_c8_12 >> 4;

  assign t_r20_c9_0 = p_19_9 << 1;
  assign t_r20_c9_1 = p_20_8 << 1;
  assign t_r20_c9_2 = p_20_9 << 2;
  assign t_r20_c9_3 = p_20_10 << 1;
  assign t_r20_c9_4 = p_21_9 << 1;
  assign t_r20_c9_5 = t_r20_c9_0 + p_19_8;
  assign t_r20_c9_6 = t_r20_c9_1 + p_19_10;
  assign t_r20_c9_7 = t_r20_c9_2 + t_r20_c9_3;
  assign t_r20_c9_8 = t_r20_c9_4 + p_21_8;
  assign t_r20_c9_9 = t_r20_c9_5 + t_r20_c9_6;
  assign t_r20_c9_10 = t_r20_c9_7 + t_r20_c9_8;
  assign t_r20_c9_11 = t_r20_c9_9 + t_r20_c9_10;
  assign t_r20_c9_12 = t_r20_c9_11 + p_21_10;
  assign out_20_9 = t_r20_c9_12 >> 4;

  assign t_r20_c10_0 = p_19_10 << 1;
  assign t_r20_c10_1 = p_20_9 << 1;
  assign t_r20_c10_2 = p_20_10 << 2;
  assign t_r20_c10_3 = p_20_11 << 1;
  assign t_r20_c10_4 = p_21_10 << 1;
  assign t_r20_c10_5 = t_r20_c10_0 + p_19_9;
  assign t_r20_c10_6 = t_r20_c10_1 + p_19_11;
  assign t_r20_c10_7 = t_r20_c10_2 + t_r20_c10_3;
  assign t_r20_c10_8 = t_r20_c10_4 + p_21_9;
  assign t_r20_c10_9 = t_r20_c10_5 + t_r20_c10_6;
  assign t_r20_c10_10 = t_r20_c10_7 + t_r20_c10_8;
  assign t_r20_c10_11 = t_r20_c10_9 + t_r20_c10_10;
  assign t_r20_c10_12 = t_r20_c10_11 + p_21_11;
  assign out_20_10 = t_r20_c10_12 >> 4;

  assign t_r20_c11_0 = p_19_11 << 1;
  assign t_r20_c11_1 = p_20_10 << 1;
  assign t_r20_c11_2 = p_20_11 << 2;
  assign t_r20_c11_3 = p_20_12 << 1;
  assign t_r20_c11_4 = p_21_11 << 1;
  assign t_r20_c11_5 = t_r20_c11_0 + p_19_10;
  assign t_r20_c11_6 = t_r20_c11_1 + p_19_12;
  assign t_r20_c11_7 = t_r20_c11_2 + t_r20_c11_3;
  assign t_r20_c11_8 = t_r20_c11_4 + p_21_10;
  assign t_r20_c11_9 = t_r20_c11_5 + t_r20_c11_6;
  assign t_r20_c11_10 = t_r20_c11_7 + t_r20_c11_8;
  assign t_r20_c11_11 = t_r20_c11_9 + t_r20_c11_10;
  assign t_r20_c11_12 = t_r20_c11_11 + p_21_12;
  assign out_20_11 = t_r20_c11_12 >> 4;

  assign t_r20_c12_0 = p_19_12 << 1;
  assign t_r20_c12_1 = p_20_11 << 1;
  assign t_r20_c12_2 = p_20_12 << 2;
  assign t_r20_c12_3 = p_20_13 << 1;
  assign t_r20_c12_4 = p_21_12 << 1;
  assign t_r20_c12_5 = t_r20_c12_0 + p_19_11;
  assign t_r20_c12_6 = t_r20_c12_1 + p_19_13;
  assign t_r20_c12_7 = t_r20_c12_2 + t_r20_c12_3;
  assign t_r20_c12_8 = t_r20_c12_4 + p_21_11;
  assign t_r20_c12_9 = t_r20_c12_5 + t_r20_c12_6;
  assign t_r20_c12_10 = t_r20_c12_7 + t_r20_c12_8;
  assign t_r20_c12_11 = t_r20_c12_9 + t_r20_c12_10;
  assign t_r20_c12_12 = t_r20_c12_11 + p_21_13;
  assign out_20_12 = t_r20_c12_12 >> 4;

  assign t_r20_c13_0 = p_19_13 << 1;
  assign t_r20_c13_1 = p_20_12 << 1;
  assign t_r20_c13_2 = p_20_13 << 2;
  assign t_r20_c13_3 = p_20_14 << 1;
  assign t_r20_c13_4 = p_21_13 << 1;
  assign t_r20_c13_5 = t_r20_c13_0 + p_19_12;
  assign t_r20_c13_6 = t_r20_c13_1 + p_19_14;
  assign t_r20_c13_7 = t_r20_c13_2 + t_r20_c13_3;
  assign t_r20_c13_8 = t_r20_c13_4 + p_21_12;
  assign t_r20_c13_9 = t_r20_c13_5 + t_r20_c13_6;
  assign t_r20_c13_10 = t_r20_c13_7 + t_r20_c13_8;
  assign t_r20_c13_11 = t_r20_c13_9 + t_r20_c13_10;
  assign t_r20_c13_12 = t_r20_c13_11 + p_21_14;
  assign out_20_13 = t_r20_c13_12 >> 4;

  assign t_r20_c14_0 = p_19_14 << 1;
  assign t_r20_c14_1 = p_20_13 << 1;
  assign t_r20_c14_2 = p_20_14 << 2;
  assign t_r20_c14_3 = p_20_15 << 1;
  assign t_r20_c14_4 = p_21_14 << 1;
  assign t_r20_c14_5 = t_r20_c14_0 + p_19_13;
  assign t_r20_c14_6 = t_r20_c14_1 + p_19_15;
  assign t_r20_c14_7 = t_r20_c14_2 + t_r20_c14_3;
  assign t_r20_c14_8 = t_r20_c14_4 + p_21_13;
  assign t_r20_c14_9 = t_r20_c14_5 + t_r20_c14_6;
  assign t_r20_c14_10 = t_r20_c14_7 + t_r20_c14_8;
  assign t_r20_c14_11 = t_r20_c14_9 + t_r20_c14_10;
  assign t_r20_c14_12 = t_r20_c14_11 + p_21_15;
  assign out_20_14 = t_r20_c14_12 >> 4;

  assign t_r20_c15_0 = p_19_15 << 1;
  assign t_r20_c15_1 = p_20_14 << 1;
  assign t_r20_c15_2 = p_20_15 << 2;
  assign t_r20_c15_3 = p_20_16 << 1;
  assign t_r20_c15_4 = p_21_15 << 1;
  assign t_r20_c15_5 = t_r20_c15_0 + p_19_14;
  assign t_r20_c15_6 = t_r20_c15_1 + p_19_16;
  assign t_r20_c15_7 = t_r20_c15_2 + t_r20_c15_3;
  assign t_r20_c15_8 = t_r20_c15_4 + p_21_14;
  assign t_r20_c15_9 = t_r20_c15_5 + t_r20_c15_6;
  assign t_r20_c15_10 = t_r20_c15_7 + t_r20_c15_8;
  assign t_r20_c15_11 = t_r20_c15_9 + t_r20_c15_10;
  assign t_r20_c15_12 = t_r20_c15_11 + p_21_16;
  assign out_20_15 = t_r20_c15_12 >> 4;

  assign t_r20_c16_0 = p_19_16 << 1;
  assign t_r20_c16_1 = p_20_15 << 1;
  assign t_r20_c16_2 = p_20_16 << 2;
  assign t_r20_c16_3 = p_20_17 << 1;
  assign t_r20_c16_4 = p_21_16 << 1;
  assign t_r20_c16_5 = t_r20_c16_0 + p_19_15;
  assign t_r20_c16_6 = t_r20_c16_1 + p_19_17;
  assign t_r20_c16_7 = t_r20_c16_2 + t_r20_c16_3;
  assign t_r20_c16_8 = t_r20_c16_4 + p_21_15;
  assign t_r20_c16_9 = t_r20_c16_5 + t_r20_c16_6;
  assign t_r20_c16_10 = t_r20_c16_7 + t_r20_c16_8;
  assign t_r20_c16_11 = t_r20_c16_9 + t_r20_c16_10;
  assign t_r20_c16_12 = t_r20_c16_11 + p_21_17;
  assign out_20_16 = t_r20_c16_12 >> 4;

  assign t_r20_c17_0 = p_19_17 << 1;
  assign t_r20_c17_1 = p_20_16 << 1;
  assign t_r20_c17_2 = p_20_17 << 2;
  assign t_r20_c17_3 = p_20_18 << 1;
  assign t_r20_c17_4 = p_21_17 << 1;
  assign t_r20_c17_5 = t_r20_c17_0 + p_19_16;
  assign t_r20_c17_6 = t_r20_c17_1 + p_19_18;
  assign t_r20_c17_7 = t_r20_c17_2 + t_r20_c17_3;
  assign t_r20_c17_8 = t_r20_c17_4 + p_21_16;
  assign t_r20_c17_9 = t_r20_c17_5 + t_r20_c17_6;
  assign t_r20_c17_10 = t_r20_c17_7 + t_r20_c17_8;
  assign t_r20_c17_11 = t_r20_c17_9 + t_r20_c17_10;
  assign t_r20_c17_12 = t_r20_c17_11 + p_21_18;
  assign out_20_17 = t_r20_c17_12 >> 4;

  assign t_r20_c18_0 = p_19_18 << 1;
  assign t_r20_c18_1 = p_20_17 << 1;
  assign t_r20_c18_2 = p_20_18 << 2;
  assign t_r20_c18_3 = p_20_19 << 1;
  assign t_r20_c18_4 = p_21_18 << 1;
  assign t_r20_c18_5 = t_r20_c18_0 + p_19_17;
  assign t_r20_c18_6 = t_r20_c18_1 + p_19_19;
  assign t_r20_c18_7 = t_r20_c18_2 + t_r20_c18_3;
  assign t_r20_c18_8 = t_r20_c18_4 + p_21_17;
  assign t_r20_c18_9 = t_r20_c18_5 + t_r20_c18_6;
  assign t_r20_c18_10 = t_r20_c18_7 + t_r20_c18_8;
  assign t_r20_c18_11 = t_r20_c18_9 + t_r20_c18_10;
  assign t_r20_c18_12 = t_r20_c18_11 + p_21_19;
  assign out_20_18 = t_r20_c18_12 >> 4;

  assign t_r20_c19_0 = p_19_19 << 1;
  assign t_r20_c19_1 = p_20_18 << 1;
  assign t_r20_c19_2 = p_20_19 << 2;
  assign t_r20_c19_3 = p_20_20 << 1;
  assign t_r20_c19_4 = p_21_19 << 1;
  assign t_r20_c19_5 = t_r20_c19_0 + p_19_18;
  assign t_r20_c19_6 = t_r20_c19_1 + p_19_20;
  assign t_r20_c19_7 = t_r20_c19_2 + t_r20_c19_3;
  assign t_r20_c19_8 = t_r20_c19_4 + p_21_18;
  assign t_r20_c19_9 = t_r20_c19_5 + t_r20_c19_6;
  assign t_r20_c19_10 = t_r20_c19_7 + t_r20_c19_8;
  assign t_r20_c19_11 = t_r20_c19_9 + t_r20_c19_10;
  assign t_r20_c19_12 = t_r20_c19_11 + p_21_20;
  assign out_20_19 = t_r20_c19_12 >> 4;

  assign t_r20_c20_0 = p_19_20 << 1;
  assign t_r20_c20_1 = p_20_19 << 1;
  assign t_r20_c20_2 = p_20_20 << 2;
  assign t_r20_c20_3 = p_20_21 << 1;
  assign t_r20_c20_4 = p_21_20 << 1;
  assign t_r20_c20_5 = t_r20_c20_0 + p_19_19;
  assign t_r20_c20_6 = t_r20_c20_1 + p_19_21;
  assign t_r20_c20_7 = t_r20_c20_2 + t_r20_c20_3;
  assign t_r20_c20_8 = t_r20_c20_4 + p_21_19;
  assign t_r20_c20_9 = t_r20_c20_5 + t_r20_c20_6;
  assign t_r20_c20_10 = t_r20_c20_7 + t_r20_c20_8;
  assign t_r20_c20_11 = t_r20_c20_9 + t_r20_c20_10;
  assign t_r20_c20_12 = t_r20_c20_11 + p_21_21;
  assign out_20_20 = t_r20_c20_12 >> 4;

  assign t_r20_c21_0 = p_19_21 << 1;
  assign t_r20_c21_1 = p_20_20 << 1;
  assign t_r20_c21_2 = p_20_21 << 2;
  assign t_r20_c21_3 = p_20_22 << 1;
  assign t_r20_c21_4 = p_21_21 << 1;
  assign t_r20_c21_5 = t_r20_c21_0 + p_19_20;
  assign t_r20_c21_6 = t_r20_c21_1 + p_19_22;
  assign t_r20_c21_7 = t_r20_c21_2 + t_r20_c21_3;
  assign t_r20_c21_8 = t_r20_c21_4 + p_21_20;
  assign t_r20_c21_9 = t_r20_c21_5 + t_r20_c21_6;
  assign t_r20_c21_10 = t_r20_c21_7 + t_r20_c21_8;
  assign t_r20_c21_11 = t_r20_c21_9 + t_r20_c21_10;
  assign t_r20_c21_12 = t_r20_c21_11 + p_21_22;
  assign out_20_21 = t_r20_c21_12 >> 4;

  assign t_r20_c22_0 = p_19_22 << 1;
  assign t_r20_c22_1 = p_20_21 << 1;
  assign t_r20_c22_2 = p_20_22 << 2;
  assign t_r20_c22_3 = p_20_23 << 1;
  assign t_r20_c22_4 = p_21_22 << 1;
  assign t_r20_c22_5 = t_r20_c22_0 + p_19_21;
  assign t_r20_c22_6 = t_r20_c22_1 + p_19_23;
  assign t_r20_c22_7 = t_r20_c22_2 + t_r20_c22_3;
  assign t_r20_c22_8 = t_r20_c22_4 + p_21_21;
  assign t_r20_c22_9 = t_r20_c22_5 + t_r20_c22_6;
  assign t_r20_c22_10 = t_r20_c22_7 + t_r20_c22_8;
  assign t_r20_c22_11 = t_r20_c22_9 + t_r20_c22_10;
  assign t_r20_c22_12 = t_r20_c22_11 + p_21_23;
  assign out_20_22 = t_r20_c22_12 >> 4;

  assign t_r20_c23_0 = p_19_23 << 1;
  assign t_r20_c23_1 = p_20_22 << 1;
  assign t_r20_c23_2 = p_20_23 << 2;
  assign t_r20_c23_3 = p_20_24 << 1;
  assign t_r20_c23_4 = p_21_23 << 1;
  assign t_r20_c23_5 = t_r20_c23_0 + p_19_22;
  assign t_r20_c23_6 = t_r20_c23_1 + p_19_24;
  assign t_r20_c23_7 = t_r20_c23_2 + t_r20_c23_3;
  assign t_r20_c23_8 = t_r20_c23_4 + p_21_22;
  assign t_r20_c23_9 = t_r20_c23_5 + t_r20_c23_6;
  assign t_r20_c23_10 = t_r20_c23_7 + t_r20_c23_8;
  assign t_r20_c23_11 = t_r20_c23_9 + t_r20_c23_10;
  assign t_r20_c23_12 = t_r20_c23_11 + p_21_24;
  assign out_20_23 = t_r20_c23_12 >> 4;

  assign t_r20_c24_0 = p_19_24 << 1;
  assign t_r20_c24_1 = p_20_23 << 1;
  assign t_r20_c24_2 = p_20_24 << 2;
  assign t_r20_c24_3 = p_20_25 << 1;
  assign t_r20_c24_4 = p_21_24 << 1;
  assign t_r20_c24_5 = t_r20_c24_0 + p_19_23;
  assign t_r20_c24_6 = t_r20_c24_1 + p_19_25;
  assign t_r20_c24_7 = t_r20_c24_2 + t_r20_c24_3;
  assign t_r20_c24_8 = t_r20_c24_4 + p_21_23;
  assign t_r20_c24_9 = t_r20_c24_5 + t_r20_c24_6;
  assign t_r20_c24_10 = t_r20_c24_7 + t_r20_c24_8;
  assign t_r20_c24_11 = t_r20_c24_9 + t_r20_c24_10;
  assign t_r20_c24_12 = t_r20_c24_11 + p_21_25;
  assign out_20_24 = t_r20_c24_12 >> 4;

  assign t_r20_c25_0 = p_19_25 << 1;
  assign t_r20_c25_1 = p_20_24 << 1;
  assign t_r20_c25_2 = p_20_25 << 2;
  assign t_r20_c25_3 = p_20_26 << 1;
  assign t_r20_c25_4 = p_21_25 << 1;
  assign t_r20_c25_5 = t_r20_c25_0 + p_19_24;
  assign t_r20_c25_6 = t_r20_c25_1 + p_19_26;
  assign t_r20_c25_7 = t_r20_c25_2 + t_r20_c25_3;
  assign t_r20_c25_8 = t_r20_c25_4 + p_21_24;
  assign t_r20_c25_9 = t_r20_c25_5 + t_r20_c25_6;
  assign t_r20_c25_10 = t_r20_c25_7 + t_r20_c25_8;
  assign t_r20_c25_11 = t_r20_c25_9 + t_r20_c25_10;
  assign t_r20_c25_12 = t_r20_c25_11 + p_21_26;
  assign out_20_25 = t_r20_c25_12 >> 4;

  assign t_r20_c26_0 = p_19_26 << 1;
  assign t_r20_c26_1 = p_20_25 << 1;
  assign t_r20_c26_2 = p_20_26 << 2;
  assign t_r20_c26_3 = p_20_27 << 1;
  assign t_r20_c26_4 = p_21_26 << 1;
  assign t_r20_c26_5 = t_r20_c26_0 + p_19_25;
  assign t_r20_c26_6 = t_r20_c26_1 + p_19_27;
  assign t_r20_c26_7 = t_r20_c26_2 + t_r20_c26_3;
  assign t_r20_c26_8 = t_r20_c26_4 + p_21_25;
  assign t_r20_c26_9 = t_r20_c26_5 + t_r20_c26_6;
  assign t_r20_c26_10 = t_r20_c26_7 + t_r20_c26_8;
  assign t_r20_c26_11 = t_r20_c26_9 + t_r20_c26_10;
  assign t_r20_c26_12 = t_r20_c26_11 + p_21_27;
  assign out_20_26 = t_r20_c26_12 >> 4;

  assign t_r20_c27_0 = p_19_27 << 1;
  assign t_r20_c27_1 = p_20_26 << 1;
  assign t_r20_c27_2 = p_20_27 << 2;
  assign t_r20_c27_3 = p_20_28 << 1;
  assign t_r20_c27_4 = p_21_27 << 1;
  assign t_r20_c27_5 = t_r20_c27_0 + p_19_26;
  assign t_r20_c27_6 = t_r20_c27_1 + p_19_28;
  assign t_r20_c27_7 = t_r20_c27_2 + t_r20_c27_3;
  assign t_r20_c27_8 = t_r20_c27_4 + p_21_26;
  assign t_r20_c27_9 = t_r20_c27_5 + t_r20_c27_6;
  assign t_r20_c27_10 = t_r20_c27_7 + t_r20_c27_8;
  assign t_r20_c27_11 = t_r20_c27_9 + t_r20_c27_10;
  assign t_r20_c27_12 = t_r20_c27_11 + p_21_28;
  assign out_20_27 = t_r20_c27_12 >> 4;

  assign t_r20_c28_0 = p_19_28 << 1;
  assign t_r20_c28_1 = p_20_27 << 1;
  assign t_r20_c28_2 = p_20_28 << 2;
  assign t_r20_c28_3 = p_20_29 << 1;
  assign t_r20_c28_4 = p_21_28 << 1;
  assign t_r20_c28_5 = t_r20_c28_0 + p_19_27;
  assign t_r20_c28_6 = t_r20_c28_1 + p_19_29;
  assign t_r20_c28_7 = t_r20_c28_2 + t_r20_c28_3;
  assign t_r20_c28_8 = t_r20_c28_4 + p_21_27;
  assign t_r20_c28_9 = t_r20_c28_5 + t_r20_c28_6;
  assign t_r20_c28_10 = t_r20_c28_7 + t_r20_c28_8;
  assign t_r20_c28_11 = t_r20_c28_9 + t_r20_c28_10;
  assign t_r20_c28_12 = t_r20_c28_11 + p_21_29;
  assign out_20_28 = t_r20_c28_12 >> 4;

  assign t_r20_c29_0 = p_19_29 << 1;
  assign t_r20_c29_1 = p_20_28 << 1;
  assign t_r20_c29_2 = p_20_29 << 2;
  assign t_r20_c29_3 = p_20_30 << 1;
  assign t_r20_c29_4 = p_21_29 << 1;
  assign t_r20_c29_5 = t_r20_c29_0 + p_19_28;
  assign t_r20_c29_6 = t_r20_c29_1 + p_19_30;
  assign t_r20_c29_7 = t_r20_c29_2 + t_r20_c29_3;
  assign t_r20_c29_8 = t_r20_c29_4 + p_21_28;
  assign t_r20_c29_9 = t_r20_c29_5 + t_r20_c29_6;
  assign t_r20_c29_10 = t_r20_c29_7 + t_r20_c29_8;
  assign t_r20_c29_11 = t_r20_c29_9 + t_r20_c29_10;
  assign t_r20_c29_12 = t_r20_c29_11 + p_21_30;
  assign out_20_29 = t_r20_c29_12 >> 4;

  assign t_r20_c30_0 = p_19_30 << 1;
  assign t_r20_c30_1 = p_20_29 << 1;
  assign t_r20_c30_2 = p_20_30 << 2;
  assign t_r20_c30_3 = p_20_31 << 1;
  assign t_r20_c30_4 = p_21_30 << 1;
  assign t_r20_c30_5 = t_r20_c30_0 + p_19_29;
  assign t_r20_c30_6 = t_r20_c30_1 + p_19_31;
  assign t_r20_c30_7 = t_r20_c30_2 + t_r20_c30_3;
  assign t_r20_c30_8 = t_r20_c30_4 + p_21_29;
  assign t_r20_c30_9 = t_r20_c30_5 + t_r20_c30_6;
  assign t_r20_c30_10 = t_r20_c30_7 + t_r20_c30_8;
  assign t_r20_c30_11 = t_r20_c30_9 + t_r20_c30_10;
  assign t_r20_c30_12 = t_r20_c30_11 + p_21_31;
  assign out_20_30 = t_r20_c30_12 >> 4;

  assign t_r20_c31_0 = p_19_31 << 1;
  assign t_r20_c31_1 = p_20_30 << 1;
  assign t_r20_c31_2 = p_20_31 << 2;
  assign t_r20_c31_3 = p_20_32 << 1;
  assign t_r20_c31_4 = p_21_31 << 1;
  assign t_r20_c31_5 = t_r20_c31_0 + p_19_30;
  assign t_r20_c31_6 = t_r20_c31_1 + p_19_32;
  assign t_r20_c31_7 = t_r20_c31_2 + t_r20_c31_3;
  assign t_r20_c31_8 = t_r20_c31_4 + p_21_30;
  assign t_r20_c31_9 = t_r20_c31_5 + t_r20_c31_6;
  assign t_r20_c31_10 = t_r20_c31_7 + t_r20_c31_8;
  assign t_r20_c31_11 = t_r20_c31_9 + t_r20_c31_10;
  assign t_r20_c31_12 = t_r20_c31_11 + p_21_32;
  assign out_20_31 = t_r20_c31_12 >> 4;

  assign t_r20_c32_0 = p_19_32 << 1;
  assign t_r20_c32_1 = p_20_31 << 1;
  assign t_r20_c32_2 = p_20_32 << 2;
  assign t_r20_c32_3 = p_20_33 << 1;
  assign t_r20_c32_4 = p_21_32 << 1;
  assign t_r20_c32_5 = t_r20_c32_0 + p_19_31;
  assign t_r20_c32_6 = t_r20_c32_1 + p_19_33;
  assign t_r20_c32_7 = t_r20_c32_2 + t_r20_c32_3;
  assign t_r20_c32_8 = t_r20_c32_4 + p_21_31;
  assign t_r20_c32_9 = t_r20_c32_5 + t_r20_c32_6;
  assign t_r20_c32_10 = t_r20_c32_7 + t_r20_c32_8;
  assign t_r20_c32_11 = t_r20_c32_9 + t_r20_c32_10;
  assign t_r20_c32_12 = t_r20_c32_11 + p_21_33;
  assign out_20_32 = t_r20_c32_12 >> 4;

  assign t_r20_c33_0 = p_19_33 << 1;
  assign t_r20_c33_1 = p_20_32 << 1;
  assign t_r20_c33_2 = p_20_33 << 2;
  assign t_r20_c33_3 = p_20_34 << 1;
  assign t_r20_c33_4 = p_21_33 << 1;
  assign t_r20_c33_5 = t_r20_c33_0 + p_19_32;
  assign t_r20_c33_6 = t_r20_c33_1 + p_19_34;
  assign t_r20_c33_7 = t_r20_c33_2 + t_r20_c33_3;
  assign t_r20_c33_8 = t_r20_c33_4 + p_21_32;
  assign t_r20_c33_9 = t_r20_c33_5 + t_r20_c33_6;
  assign t_r20_c33_10 = t_r20_c33_7 + t_r20_c33_8;
  assign t_r20_c33_11 = t_r20_c33_9 + t_r20_c33_10;
  assign t_r20_c33_12 = t_r20_c33_11 + p_21_34;
  assign out_20_33 = t_r20_c33_12 >> 4;

  assign t_r20_c34_0 = p_19_34 << 1;
  assign t_r20_c34_1 = p_20_33 << 1;
  assign t_r20_c34_2 = p_20_34 << 2;
  assign t_r20_c34_3 = p_20_35 << 1;
  assign t_r20_c34_4 = p_21_34 << 1;
  assign t_r20_c34_5 = t_r20_c34_0 + p_19_33;
  assign t_r20_c34_6 = t_r20_c34_1 + p_19_35;
  assign t_r20_c34_7 = t_r20_c34_2 + t_r20_c34_3;
  assign t_r20_c34_8 = t_r20_c34_4 + p_21_33;
  assign t_r20_c34_9 = t_r20_c34_5 + t_r20_c34_6;
  assign t_r20_c34_10 = t_r20_c34_7 + t_r20_c34_8;
  assign t_r20_c34_11 = t_r20_c34_9 + t_r20_c34_10;
  assign t_r20_c34_12 = t_r20_c34_11 + p_21_35;
  assign out_20_34 = t_r20_c34_12 >> 4;

  assign t_r20_c35_0 = p_19_35 << 1;
  assign t_r20_c35_1 = p_20_34 << 1;
  assign t_r20_c35_2 = p_20_35 << 2;
  assign t_r20_c35_3 = p_20_36 << 1;
  assign t_r20_c35_4 = p_21_35 << 1;
  assign t_r20_c35_5 = t_r20_c35_0 + p_19_34;
  assign t_r20_c35_6 = t_r20_c35_1 + p_19_36;
  assign t_r20_c35_7 = t_r20_c35_2 + t_r20_c35_3;
  assign t_r20_c35_8 = t_r20_c35_4 + p_21_34;
  assign t_r20_c35_9 = t_r20_c35_5 + t_r20_c35_6;
  assign t_r20_c35_10 = t_r20_c35_7 + t_r20_c35_8;
  assign t_r20_c35_11 = t_r20_c35_9 + t_r20_c35_10;
  assign t_r20_c35_12 = t_r20_c35_11 + p_21_36;
  assign out_20_35 = t_r20_c35_12 >> 4;

  assign t_r20_c36_0 = p_19_36 << 1;
  assign t_r20_c36_1 = p_20_35 << 1;
  assign t_r20_c36_2 = p_20_36 << 2;
  assign t_r20_c36_3 = p_20_37 << 1;
  assign t_r20_c36_4 = p_21_36 << 1;
  assign t_r20_c36_5 = t_r20_c36_0 + p_19_35;
  assign t_r20_c36_6 = t_r20_c36_1 + p_19_37;
  assign t_r20_c36_7 = t_r20_c36_2 + t_r20_c36_3;
  assign t_r20_c36_8 = t_r20_c36_4 + p_21_35;
  assign t_r20_c36_9 = t_r20_c36_5 + t_r20_c36_6;
  assign t_r20_c36_10 = t_r20_c36_7 + t_r20_c36_8;
  assign t_r20_c36_11 = t_r20_c36_9 + t_r20_c36_10;
  assign t_r20_c36_12 = t_r20_c36_11 + p_21_37;
  assign out_20_36 = t_r20_c36_12 >> 4;

  assign t_r20_c37_0 = p_19_37 << 1;
  assign t_r20_c37_1 = p_20_36 << 1;
  assign t_r20_c37_2 = p_20_37 << 2;
  assign t_r20_c37_3 = p_20_38 << 1;
  assign t_r20_c37_4 = p_21_37 << 1;
  assign t_r20_c37_5 = t_r20_c37_0 + p_19_36;
  assign t_r20_c37_6 = t_r20_c37_1 + p_19_38;
  assign t_r20_c37_7 = t_r20_c37_2 + t_r20_c37_3;
  assign t_r20_c37_8 = t_r20_c37_4 + p_21_36;
  assign t_r20_c37_9 = t_r20_c37_5 + t_r20_c37_6;
  assign t_r20_c37_10 = t_r20_c37_7 + t_r20_c37_8;
  assign t_r20_c37_11 = t_r20_c37_9 + t_r20_c37_10;
  assign t_r20_c37_12 = t_r20_c37_11 + p_21_38;
  assign out_20_37 = t_r20_c37_12 >> 4;

  assign t_r20_c38_0 = p_19_38 << 1;
  assign t_r20_c38_1 = p_20_37 << 1;
  assign t_r20_c38_2 = p_20_38 << 2;
  assign t_r20_c38_3 = p_20_39 << 1;
  assign t_r20_c38_4 = p_21_38 << 1;
  assign t_r20_c38_5 = t_r20_c38_0 + p_19_37;
  assign t_r20_c38_6 = t_r20_c38_1 + p_19_39;
  assign t_r20_c38_7 = t_r20_c38_2 + t_r20_c38_3;
  assign t_r20_c38_8 = t_r20_c38_4 + p_21_37;
  assign t_r20_c38_9 = t_r20_c38_5 + t_r20_c38_6;
  assign t_r20_c38_10 = t_r20_c38_7 + t_r20_c38_8;
  assign t_r20_c38_11 = t_r20_c38_9 + t_r20_c38_10;
  assign t_r20_c38_12 = t_r20_c38_11 + p_21_39;
  assign out_20_38 = t_r20_c38_12 >> 4;

  assign t_r20_c39_0 = p_19_39 << 1;
  assign t_r20_c39_1 = p_20_38 << 1;
  assign t_r20_c39_2 = p_20_39 << 2;
  assign t_r20_c39_3 = p_20_40 << 1;
  assign t_r20_c39_4 = p_21_39 << 1;
  assign t_r20_c39_5 = t_r20_c39_0 + p_19_38;
  assign t_r20_c39_6 = t_r20_c39_1 + p_19_40;
  assign t_r20_c39_7 = t_r20_c39_2 + t_r20_c39_3;
  assign t_r20_c39_8 = t_r20_c39_4 + p_21_38;
  assign t_r20_c39_9 = t_r20_c39_5 + t_r20_c39_6;
  assign t_r20_c39_10 = t_r20_c39_7 + t_r20_c39_8;
  assign t_r20_c39_11 = t_r20_c39_9 + t_r20_c39_10;
  assign t_r20_c39_12 = t_r20_c39_11 + p_21_40;
  assign out_20_39 = t_r20_c39_12 >> 4;

  assign t_r20_c40_0 = p_19_40 << 1;
  assign t_r20_c40_1 = p_20_39 << 1;
  assign t_r20_c40_2 = p_20_40 << 2;
  assign t_r20_c40_3 = p_20_41 << 1;
  assign t_r20_c40_4 = p_21_40 << 1;
  assign t_r20_c40_5 = t_r20_c40_0 + p_19_39;
  assign t_r20_c40_6 = t_r20_c40_1 + p_19_41;
  assign t_r20_c40_7 = t_r20_c40_2 + t_r20_c40_3;
  assign t_r20_c40_8 = t_r20_c40_4 + p_21_39;
  assign t_r20_c40_9 = t_r20_c40_5 + t_r20_c40_6;
  assign t_r20_c40_10 = t_r20_c40_7 + t_r20_c40_8;
  assign t_r20_c40_11 = t_r20_c40_9 + t_r20_c40_10;
  assign t_r20_c40_12 = t_r20_c40_11 + p_21_41;
  assign out_20_40 = t_r20_c40_12 >> 4;

  assign t_r20_c41_0 = p_19_41 << 1;
  assign t_r20_c41_1 = p_20_40 << 1;
  assign t_r20_c41_2 = p_20_41 << 2;
  assign t_r20_c41_3 = p_20_42 << 1;
  assign t_r20_c41_4 = p_21_41 << 1;
  assign t_r20_c41_5 = t_r20_c41_0 + p_19_40;
  assign t_r20_c41_6 = t_r20_c41_1 + p_19_42;
  assign t_r20_c41_7 = t_r20_c41_2 + t_r20_c41_3;
  assign t_r20_c41_8 = t_r20_c41_4 + p_21_40;
  assign t_r20_c41_9 = t_r20_c41_5 + t_r20_c41_6;
  assign t_r20_c41_10 = t_r20_c41_7 + t_r20_c41_8;
  assign t_r20_c41_11 = t_r20_c41_9 + t_r20_c41_10;
  assign t_r20_c41_12 = t_r20_c41_11 + p_21_42;
  assign out_20_41 = t_r20_c41_12 >> 4;

  assign t_r20_c42_0 = p_19_42 << 1;
  assign t_r20_c42_1 = p_20_41 << 1;
  assign t_r20_c42_2 = p_20_42 << 2;
  assign t_r20_c42_3 = p_20_43 << 1;
  assign t_r20_c42_4 = p_21_42 << 1;
  assign t_r20_c42_5 = t_r20_c42_0 + p_19_41;
  assign t_r20_c42_6 = t_r20_c42_1 + p_19_43;
  assign t_r20_c42_7 = t_r20_c42_2 + t_r20_c42_3;
  assign t_r20_c42_8 = t_r20_c42_4 + p_21_41;
  assign t_r20_c42_9 = t_r20_c42_5 + t_r20_c42_6;
  assign t_r20_c42_10 = t_r20_c42_7 + t_r20_c42_8;
  assign t_r20_c42_11 = t_r20_c42_9 + t_r20_c42_10;
  assign t_r20_c42_12 = t_r20_c42_11 + p_21_43;
  assign out_20_42 = t_r20_c42_12 >> 4;

  assign t_r20_c43_0 = p_19_43 << 1;
  assign t_r20_c43_1 = p_20_42 << 1;
  assign t_r20_c43_2 = p_20_43 << 2;
  assign t_r20_c43_3 = p_20_44 << 1;
  assign t_r20_c43_4 = p_21_43 << 1;
  assign t_r20_c43_5 = t_r20_c43_0 + p_19_42;
  assign t_r20_c43_6 = t_r20_c43_1 + p_19_44;
  assign t_r20_c43_7 = t_r20_c43_2 + t_r20_c43_3;
  assign t_r20_c43_8 = t_r20_c43_4 + p_21_42;
  assign t_r20_c43_9 = t_r20_c43_5 + t_r20_c43_6;
  assign t_r20_c43_10 = t_r20_c43_7 + t_r20_c43_8;
  assign t_r20_c43_11 = t_r20_c43_9 + t_r20_c43_10;
  assign t_r20_c43_12 = t_r20_c43_11 + p_21_44;
  assign out_20_43 = t_r20_c43_12 >> 4;

  assign t_r20_c44_0 = p_19_44 << 1;
  assign t_r20_c44_1 = p_20_43 << 1;
  assign t_r20_c44_2 = p_20_44 << 2;
  assign t_r20_c44_3 = p_20_45 << 1;
  assign t_r20_c44_4 = p_21_44 << 1;
  assign t_r20_c44_5 = t_r20_c44_0 + p_19_43;
  assign t_r20_c44_6 = t_r20_c44_1 + p_19_45;
  assign t_r20_c44_7 = t_r20_c44_2 + t_r20_c44_3;
  assign t_r20_c44_8 = t_r20_c44_4 + p_21_43;
  assign t_r20_c44_9 = t_r20_c44_5 + t_r20_c44_6;
  assign t_r20_c44_10 = t_r20_c44_7 + t_r20_c44_8;
  assign t_r20_c44_11 = t_r20_c44_9 + t_r20_c44_10;
  assign t_r20_c44_12 = t_r20_c44_11 + p_21_45;
  assign out_20_44 = t_r20_c44_12 >> 4;

  assign t_r20_c45_0 = p_19_45 << 1;
  assign t_r20_c45_1 = p_20_44 << 1;
  assign t_r20_c45_2 = p_20_45 << 2;
  assign t_r20_c45_3 = p_20_46 << 1;
  assign t_r20_c45_4 = p_21_45 << 1;
  assign t_r20_c45_5 = t_r20_c45_0 + p_19_44;
  assign t_r20_c45_6 = t_r20_c45_1 + p_19_46;
  assign t_r20_c45_7 = t_r20_c45_2 + t_r20_c45_3;
  assign t_r20_c45_8 = t_r20_c45_4 + p_21_44;
  assign t_r20_c45_9 = t_r20_c45_5 + t_r20_c45_6;
  assign t_r20_c45_10 = t_r20_c45_7 + t_r20_c45_8;
  assign t_r20_c45_11 = t_r20_c45_9 + t_r20_c45_10;
  assign t_r20_c45_12 = t_r20_c45_11 + p_21_46;
  assign out_20_45 = t_r20_c45_12 >> 4;

  assign t_r20_c46_0 = p_19_46 << 1;
  assign t_r20_c46_1 = p_20_45 << 1;
  assign t_r20_c46_2 = p_20_46 << 2;
  assign t_r20_c46_3 = p_20_47 << 1;
  assign t_r20_c46_4 = p_21_46 << 1;
  assign t_r20_c46_5 = t_r20_c46_0 + p_19_45;
  assign t_r20_c46_6 = t_r20_c46_1 + p_19_47;
  assign t_r20_c46_7 = t_r20_c46_2 + t_r20_c46_3;
  assign t_r20_c46_8 = t_r20_c46_4 + p_21_45;
  assign t_r20_c46_9 = t_r20_c46_5 + t_r20_c46_6;
  assign t_r20_c46_10 = t_r20_c46_7 + t_r20_c46_8;
  assign t_r20_c46_11 = t_r20_c46_9 + t_r20_c46_10;
  assign t_r20_c46_12 = t_r20_c46_11 + p_21_47;
  assign out_20_46 = t_r20_c46_12 >> 4;

  assign t_r20_c47_0 = p_19_47 << 1;
  assign t_r20_c47_1 = p_20_46 << 1;
  assign t_r20_c47_2 = p_20_47 << 2;
  assign t_r20_c47_3 = p_20_48 << 1;
  assign t_r20_c47_4 = p_21_47 << 1;
  assign t_r20_c47_5 = t_r20_c47_0 + p_19_46;
  assign t_r20_c47_6 = t_r20_c47_1 + p_19_48;
  assign t_r20_c47_7 = t_r20_c47_2 + t_r20_c47_3;
  assign t_r20_c47_8 = t_r20_c47_4 + p_21_46;
  assign t_r20_c47_9 = t_r20_c47_5 + t_r20_c47_6;
  assign t_r20_c47_10 = t_r20_c47_7 + t_r20_c47_8;
  assign t_r20_c47_11 = t_r20_c47_9 + t_r20_c47_10;
  assign t_r20_c47_12 = t_r20_c47_11 + p_21_48;
  assign out_20_47 = t_r20_c47_12 >> 4;

  assign t_r20_c48_0 = p_19_48 << 1;
  assign t_r20_c48_1 = p_20_47 << 1;
  assign t_r20_c48_2 = p_20_48 << 2;
  assign t_r20_c48_3 = p_20_49 << 1;
  assign t_r20_c48_4 = p_21_48 << 1;
  assign t_r20_c48_5 = t_r20_c48_0 + p_19_47;
  assign t_r20_c48_6 = t_r20_c48_1 + p_19_49;
  assign t_r20_c48_7 = t_r20_c48_2 + t_r20_c48_3;
  assign t_r20_c48_8 = t_r20_c48_4 + p_21_47;
  assign t_r20_c48_9 = t_r20_c48_5 + t_r20_c48_6;
  assign t_r20_c48_10 = t_r20_c48_7 + t_r20_c48_8;
  assign t_r20_c48_11 = t_r20_c48_9 + t_r20_c48_10;
  assign t_r20_c48_12 = t_r20_c48_11 + p_21_49;
  assign out_20_48 = t_r20_c48_12 >> 4;

  assign t_r20_c49_0 = p_19_49 << 1;
  assign t_r20_c49_1 = p_20_48 << 1;
  assign t_r20_c49_2 = p_20_49 << 2;
  assign t_r20_c49_3 = p_20_50 << 1;
  assign t_r20_c49_4 = p_21_49 << 1;
  assign t_r20_c49_5 = t_r20_c49_0 + p_19_48;
  assign t_r20_c49_6 = t_r20_c49_1 + p_19_50;
  assign t_r20_c49_7 = t_r20_c49_2 + t_r20_c49_3;
  assign t_r20_c49_8 = t_r20_c49_4 + p_21_48;
  assign t_r20_c49_9 = t_r20_c49_5 + t_r20_c49_6;
  assign t_r20_c49_10 = t_r20_c49_7 + t_r20_c49_8;
  assign t_r20_c49_11 = t_r20_c49_9 + t_r20_c49_10;
  assign t_r20_c49_12 = t_r20_c49_11 + p_21_50;
  assign out_20_49 = t_r20_c49_12 >> 4;

  assign t_r20_c50_0 = p_19_50 << 1;
  assign t_r20_c50_1 = p_20_49 << 1;
  assign t_r20_c50_2 = p_20_50 << 2;
  assign t_r20_c50_3 = p_20_51 << 1;
  assign t_r20_c50_4 = p_21_50 << 1;
  assign t_r20_c50_5 = t_r20_c50_0 + p_19_49;
  assign t_r20_c50_6 = t_r20_c50_1 + p_19_51;
  assign t_r20_c50_7 = t_r20_c50_2 + t_r20_c50_3;
  assign t_r20_c50_8 = t_r20_c50_4 + p_21_49;
  assign t_r20_c50_9 = t_r20_c50_5 + t_r20_c50_6;
  assign t_r20_c50_10 = t_r20_c50_7 + t_r20_c50_8;
  assign t_r20_c50_11 = t_r20_c50_9 + t_r20_c50_10;
  assign t_r20_c50_12 = t_r20_c50_11 + p_21_51;
  assign out_20_50 = t_r20_c50_12 >> 4;

  assign t_r20_c51_0 = p_19_51 << 1;
  assign t_r20_c51_1 = p_20_50 << 1;
  assign t_r20_c51_2 = p_20_51 << 2;
  assign t_r20_c51_3 = p_20_52 << 1;
  assign t_r20_c51_4 = p_21_51 << 1;
  assign t_r20_c51_5 = t_r20_c51_0 + p_19_50;
  assign t_r20_c51_6 = t_r20_c51_1 + p_19_52;
  assign t_r20_c51_7 = t_r20_c51_2 + t_r20_c51_3;
  assign t_r20_c51_8 = t_r20_c51_4 + p_21_50;
  assign t_r20_c51_9 = t_r20_c51_5 + t_r20_c51_6;
  assign t_r20_c51_10 = t_r20_c51_7 + t_r20_c51_8;
  assign t_r20_c51_11 = t_r20_c51_9 + t_r20_c51_10;
  assign t_r20_c51_12 = t_r20_c51_11 + p_21_52;
  assign out_20_51 = t_r20_c51_12 >> 4;

  assign t_r20_c52_0 = p_19_52 << 1;
  assign t_r20_c52_1 = p_20_51 << 1;
  assign t_r20_c52_2 = p_20_52 << 2;
  assign t_r20_c52_3 = p_20_53 << 1;
  assign t_r20_c52_4 = p_21_52 << 1;
  assign t_r20_c52_5 = t_r20_c52_0 + p_19_51;
  assign t_r20_c52_6 = t_r20_c52_1 + p_19_53;
  assign t_r20_c52_7 = t_r20_c52_2 + t_r20_c52_3;
  assign t_r20_c52_8 = t_r20_c52_4 + p_21_51;
  assign t_r20_c52_9 = t_r20_c52_5 + t_r20_c52_6;
  assign t_r20_c52_10 = t_r20_c52_7 + t_r20_c52_8;
  assign t_r20_c52_11 = t_r20_c52_9 + t_r20_c52_10;
  assign t_r20_c52_12 = t_r20_c52_11 + p_21_53;
  assign out_20_52 = t_r20_c52_12 >> 4;

  assign t_r20_c53_0 = p_19_53 << 1;
  assign t_r20_c53_1 = p_20_52 << 1;
  assign t_r20_c53_2 = p_20_53 << 2;
  assign t_r20_c53_3 = p_20_54 << 1;
  assign t_r20_c53_4 = p_21_53 << 1;
  assign t_r20_c53_5 = t_r20_c53_0 + p_19_52;
  assign t_r20_c53_6 = t_r20_c53_1 + p_19_54;
  assign t_r20_c53_7 = t_r20_c53_2 + t_r20_c53_3;
  assign t_r20_c53_8 = t_r20_c53_4 + p_21_52;
  assign t_r20_c53_9 = t_r20_c53_5 + t_r20_c53_6;
  assign t_r20_c53_10 = t_r20_c53_7 + t_r20_c53_8;
  assign t_r20_c53_11 = t_r20_c53_9 + t_r20_c53_10;
  assign t_r20_c53_12 = t_r20_c53_11 + p_21_54;
  assign out_20_53 = t_r20_c53_12 >> 4;

  assign t_r20_c54_0 = p_19_54 << 1;
  assign t_r20_c54_1 = p_20_53 << 1;
  assign t_r20_c54_2 = p_20_54 << 2;
  assign t_r20_c54_3 = p_20_55 << 1;
  assign t_r20_c54_4 = p_21_54 << 1;
  assign t_r20_c54_5 = t_r20_c54_0 + p_19_53;
  assign t_r20_c54_6 = t_r20_c54_1 + p_19_55;
  assign t_r20_c54_7 = t_r20_c54_2 + t_r20_c54_3;
  assign t_r20_c54_8 = t_r20_c54_4 + p_21_53;
  assign t_r20_c54_9 = t_r20_c54_5 + t_r20_c54_6;
  assign t_r20_c54_10 = t_r20_c54_7 + t_r20_c54_8;
  assign t_r20_c54_11 = t_r20_c54_9 + t_r20_c54_10;
  assign t_r20_c54_12 = t_r20_c54_11 + p_21_55;
  assign out_20_54 = t_r20_c54_12 >> 4;

  assign t_r20_c55_0 = p_19_55 << 1;
  assign t_r20_c55_1 = p_20_54 << 1;
  assign t_r20_c55_2 = p_20_55 << 2;
  assign t_r20_c55_3 = p_20_56 << 1;
  assign t_r20_c55_4 = p_21_55 << 1;
  assign t_r20_c55_5 = t_r20_c55_0 + p_19_54;
  assign t_r20_c55_6 = t_r20_c55_1 + p_19_56;
  assign t_r20_c55_7 = t_r20_c55_2 + t_r20_c55_3;
  assign t_r20_c55_8 = t_r20_c55_4 + p_21_54;
  assign t_r20_c55_9 = t_r20_c55_5 + t_r20_c55_6;
  assign t_r20_c55_10 = t_r20_c55_7 + t_r20_c55_8;
  assign t_r20_c55_11 = t_r20_c55_9 + t_r20_c55_10;
  assign t_r20_c55_12 = t_r20_c55_11 + p_21_56;
  assign out_20_55 = t_r20_c55_12 >> 4;

  assign t_r20_c56_0 = p_19_56 << 1;
  assign t_r20_c56_1 = p_20_55 << 1;
  assign t_r20_c56_2 = p_20_56 << 2;
  assign t_r20_c56_3 = p_20_57 << 1;
  assign t_r20_c56_4 = p_21_56 << 1;
  assign t_r20_c56_5 = t_r20_c56_0 + p_19_55;
  assign t_r20_c56_6 = t_r20_c56_1 + p_19_57;
  assign t_r20_c56_7 = t_r20_c56_2 + t_r20_c56_3;
  assign t_r20_c56_8 = t_r20_c56_4 + p_21_55;
  assign t_r20_c56_9 = t_r20_c56_5 + t_r20_c56_6;
  assign t_r20_c56_10 = t_r20_c56_7 + t_r20_c56_8;
  assign t_r20_c56_11 = t_r20_c56_9 + t_r20_c56_10;
  assign t_r20_c56_12 = t_r20_c56_11 + p_21_57;
  assign out_20_56 = t_r20_c56_12 >> 4;

  assign t_r20_c57_0 = p_19_57 << 1;
  assign t_r20_c57_1 = p_20_56 << 1;
  assign t_r20_c57_2 = p_20_57 << 2;
  assign t_r20_c57_3 = p_20_58 << 1;
  assign t_r20_c57_4 = p_21_57 << 1;
  assign t_r20_c57_5 = t_r20_c57_0 + p_19_56;
  assign t_r20_c57_6 = t_r20_c57_1 + p_19_58;
  assign t_r20_c57_7 = t_r20_c57_2 + t_r20_c57_3;
  assign t_r20_c57_8 = t_r20_c57_4 + p_21_56;
  assign t_r20_c57_9 = t_r20_c57_5 + t_r20_c57_6;
  assign t_r20_c57_10 = t_r20_c57_7 + t_r20_c57_8;
  assign t_r20_c57_11 = t_r20_c57_9 + t_r20_c57_10;
  assign t_r20_c57_12 = t_r20_c57_11 + p_21_58;
  assign out_20_57 = t_r20_c57_12 >> 4;

  assign t_r20_c58_0 = p_19_58 << 1;
  assign t_r20_c58_1 = p_20_57 << 1;
  assign t_r20_c58_2 = p_20_58 << 2;
  assign t_r20_c58_3 = p_20_59 << 1;
  assign t_r20_c58_4 = p_21_58 << 1;
  assign t_r20_c58_5 = t_r20_c58_0 + p_19_57;
  assign t_r20_c58_6 = t_r20_c58_1 + p_19_59;
  assign t_r20_c58_7 = t_r20_c58_2 + t_r20_c58_3;
  assign t_r20_c58_8 = t_r20_c58_4 + p_21_57;
  assign t_r20_c58_9 = t_r20_c58_5 + t_r20_c58_6;
  assign t_r20_c58_10 = t_r20_c58_7 + t_r20_c58_8;
  assign t_r20_c58_11 = t_r20_c58_9 + t_r20_c58_10;
  assign t_r20_c58_12 = t_r20_c58_11 + p_21_59;
  assign out_20_58 = t_r20_c58_12 >> 4;

  assign t_r20_c59_0 = p_19_59 << 1;
  assign t_r20_c59_1 = p_20_58 << 1;
  assign t_r20_c59_2 = p_20_59 << 2;
  assign t_r20_c59_3 = p_20_60 << 1;
  assign t_r20_c59_4 = p_21_59 << 1;
  assign t_r20_c59_5 = t_r20_c59_0 + p_19_58;
  assign t_r20_c59_6 = t_r20_c59_1 + p_19_60;
  assign t_r20_c59_7 = t_r20_c59_2 + t_r20_c59_3;
  assign t_r20_c59_8 = t_r20_c59_4 + p_21_58;
  assign t_r20_c59_9 = t_r20_c59_5 + t_r20_c59_6;
  assign t_r20_c59_10 = t_r20_c59_7 + t_r20_c59_8;
  assign t_r20_c59_11 = t_r20_c59_9 + t_r20_c59_10;
  assign t_r20_c59_12 = t_r20_c59_11 + p_21_60;
  assign out_20_59 = t_r20_c59_12 >> 4;

  assign t_r20_c60_0 = p_19_60 << 1;
  assign t_r20_c60_1 = p_20_59 << 1;
  assign t_r20_c60_2 = p_20_60 << 2;
  assign t_r20_c60_3 = p_20_61 << 1;
  assign t_r20_c60_4 = p_21_60 << 1;
  assign t_r20_c60_5 = t_r20_c60_0 + p_19_59;
  assign t_r20_c60_6 = t_r20_c60_1 + p_19_61;
  assign t_r20_c60_7 = t_r20_c60_2 + t_r20_c60_3;
  assign t_r20_c60_8 = t_r20_c60_4 + p_21_59;
  assign t_r20_c60_9 = t_r20_c60_5 + t_r20_c60_6;
  assign t_r20_c60_10 = t_r20_c60_7 + t_r20_c60_8;
  assign t_r20_c60_11 = t_r20_c60_9 + t_r20_c60_10;
  assign t_r20_c60_12 = t_r20_c60_11 + p_21_61;
  assign out_20_60 = t_r20_c60_12 >> 4;

  assign t_r20_c61_0 = p_19_61 << 1;
  assign t_r20_c61_1 = p_20_60 << 1;
  assign t_r20_c61_2 = p_20_61 << 2;
  assign t_r20_c61_3 = p_20_62 << 1;
  assign t_r20_c61_4 = p_21_61 << 1;
  assign t_r20_c61_5 = t_r20_c61_0 + p_19_60;
  assign t_r20_c61_6 = t_r20_c61_1 + p_19_62;
  assign t_r20_c61_7 = t_r20_c61_2 + t_r20_c61_3;
  assign t_r20_c61_8 = t_r20_c61_4 + p_21_60;
  assign t_r20_c61_9 = t_r20_c61_5 + t_r20_c61_6;
  assign t_r20_c61_10 = t_r20_c61_7 + t_r20_c61_8;
  assign t_r20_c61_11 = t_r20_c61_9 + t_r20_c61_10;
  assign t_r20_c61_12 = t_r20_c61_11 + p_21_62;
  assign out_20_61 = t_r20_c61_12 >> 4;

  assign t_r20_c62_0 = p_19_62 << 1;
  assign t_r20_c62_1 = p_20_61 << 1;
  assign t_r20_c62_2 = p_20_62 << 2;
  assign t_r20_c62_3 = p_20_63 << 1;
  assign t_r20_c62_4 = p_21_62 << 1;
  assign t_r20_c62_5 = t_r20_c62_0 + p_19_61;
  assign t_r20_c62_6 = t_r20_c62_1 + p_19_63;
  assign t_r20_c62_7 = t_r20_c62_2 + t_r20_c62_3;
  assign t_r20_c62_8 = t_r20_c62_4 + p_21_61;
  assign t_r20_c62_9 = t_r20_c62_5 + t_r20_c62_6;
  assign t_r20_c62_10 = t_r20_c62_7 + t_r20_c62_8;
  assign t_r20_c62_11 = t_r20_c62_9 + t_r20_c62_10;
  assign t_r20_c62_12 = t_r20_c62_11 + p_21_63;
  assign out_20_62 = t_r20_c62_12 >> 4;

  assign t_r20_c63_0 = p_19_63 << 1;
  assign t_r20_c63_1 = p_20_62 << 1;
  assign t_r20_c63_2 = p_20_63 << 2;
  assign t_r20_c63_3 = p_20_64 << 1;
  assign t_r20_c63_4 = p_21_63 << 1;
  assign t_r20_c63_5 = t_r20_c63_0 + p_19_62;
  assign t_r20_c63_6 = t_r20_c63_1 + p_19_64;
  assign t_r20_c63_7 = t_r20_c63_2 + t_r20_c63_3;
  assign t_r20_c63_8 = t_r20_c63_4 + p_21_62;
  assign t_r20_c63_9 = t_r20_c63_5 + t_r20_c63_6;
  assign t_r20_c63_10 = t_r20_c63_7 + t_r20_c63_8;
  assign t_r20_c63_11 = t_r20_c63_9 + t_r20_c63_10;
  assign t_r20_c63_12 = t_r20_c63_11 + p_21_64;
  assign out_20_63 = t_r20_c63_12 >> 4;

  assign t_r20_c64_0 = p_19_64 << 1;
  assign t_r20_c64_1 = p_20_63 << 1;
  assign t_r20_c64_2 = p_20_64 << 2;
  assign t_r20_c64_3 = p_20_65 << 1;
  assign t_r20_c64_4 = p_21_64 << 1;
  assign t_r20_c64_5 = t_r20_c64_0 + p_19_63;
  assign t_r20_c64_6 = t_r20_c64_1 + p_19_65;
  assign t_r20_c64_7 = t_r20_c64_2 + t_r20_c64_3;
  assign t_r20_c64_8 = t_r20_c64_4 + p_21_63;
  assign t_r20_c64_9 = t_r20_c64_5 + t_r20_c64_6;
  assign t_r20_c64_10 = t_r20_c64_7 + t_r20_c64_8;
  assign t_r20_c64_11 = t_r20_c64_9 + t_r20_c64_10;
  assign t_r20_c64_12 = t_r20_c64_11 + p_21_65;
  assign out_20_64 = t_r20_c64_12 >> 4;

  assign t_r21_c1_0 = p_20_1 << 1;
  assign t_r21_c1_1 = p_21_0 << 1;
  assign t_r21_c1_2 = p_21_1 << 2;
  assign t_r21_c1_3 = p_21_2 << 1;
  assign t_r21_c1_4 = p_22_1 << 1;
  assign t_r21_c1_5 = t_r21_c1_0 + p_20_0;
  assign t_r21_c1_6 = t_r21_c1_1 + p_20_2;
  assign t_r21_c1_7 = t_r21_c1_2 + t_r21_c1_3;
  assign t_r21_c1_8 = t_r21_c1_4 + p_22_0;
  assign t_r21_c1_9 = t_r21_c1_5 + t_r21_c1_6;
  assign t_r21_c1_10 = t_r21_c1_7 + t_r21_c1_8;
  assign t_r21_c1_11 = t_r21_c1_9 + t_r21_c1_10;
  assign t_r21_c1_12 = t_r21_c1_11 + p_22_2;
  assign out_21_1 = t_r21_c1_12 >> 4;

  assign t_r21_c2_0 = p_20_2 << 1;
  assign t_r21_c2_1 = p_21_1 << 1;
  assign t_r21_c2_2 = p_21_2 << 2;
  assign t_r21_c2_3 = p_21_3 << 1;
  assign t_r21_c2_4 = p_22_2 << 1;
  assign t_r21_c2_5 = t_r21_c2_0 + p_20_1;
  assign t_r21_c2_6 = t_r21_c2_1 + p_20_3;
  assign t_r21_c2_7 = t_r21_c2_2 + t_r21_c2_3;
  assign t_r21_c2_8 = t_r21_c2_4 + p_22_1;
  assign t_r21_c2_9 = t_r21_c2_5 + t_r21_c2_6;
  assign t_r21_c2_10 = t_r21_c2_7 + t_r21_c2_8;
  assign t_r21_c2_11 = t_r21_c2_9 + t_r21_c2_10;
  assign t_r21_c2_12 = t_r21_c2_11 + p_22_3;
  assign out_21_2 = t_r21_c2_12 >> 4;

  assign t_r21_c3_0 = p_20_3 << 1;
  assign t_r21_c3_1 = p_21_2 << 1;
  assign t_r21_c3_2 = p_21_3 << 2;
  assign t_r21_c3_3 = p_21_4 << 1;
  assign t_r21_c3_4 = p_22_3 << 1;
  assign t_r21_c3_5 = t_r21_c3_0 + p_20_2;
  assign t_r21_c3_6 = t_r21_c3_1 + p_20_4;
  assign t_r21_c3_7 = t_r21_c3_2 + t_r21_c3_3;
  assign t_r21_c3_8 = t_r21_c3_4 + p_22_2;
  assign t_r21_c3_9 = t_r21_c3_5 + t_r21_c3_6;
  assign t_r21_c3_10 = t_r21_c3_7 + t_r21_c3_8;
  assign t_r21_c3_11 = t_r21_c3_9 + t_r21_c3_10;
  assign t_r21_c3_12 = t_r21_c3_11 + p_22_4;
  assign out_21_3 = t_r21_c3_12 >> 4;

  assign t_r21_c4_0 = p_20_4 << 1;
  assign t_r21_c4_1 = p_21_3 << 1;
  assign t_r21_c4_2 = p_21_4 << 2;
  assign t_r21_c4_3 = p_21_5 << 1;
  assign t_r21_c4_4 = p_22_4 << 1;
  assign t_r21_c4_5 = t_r21_c4_0 + p_20_3;
  assign t_r21_c4_6 = t_r21_c4_1 + p_20_5;
  assign t_r21_c4_7 = t_r21_c4_2 + t_r21_c4_3;
  assign t_r21_c4_8 = t_r21_c4_4 + p_22_3;
  assign t_r21_c4_9 = t_r21_c4_5 + t_r21_c4_6;
  assign t_r21_c4_10 = t_r21_c4_7 + t_r21_c4_8;
  assign t_r21_c4_11 = t_r21_c4_9 + t_r21_c4_10;
  assign t_r21_c4_12 = t_r21_c4_11 + p_22_5;
  assign out_21_4 = t_r21_c4_12 >> 4;

  assign t_r21_c5_0 = p_20_5 << 1;
  assign t_r21_c5_1 = p_21_4 << 1;
  assign t_r21_c5_2 = p_21_5 << 2;
  assign t_r21_c5_3 = p_21_6 << 1;
  assign t_r21_c5_4 = p_22_5 << 1;
  assign t_r21_c5_5 = t_r21_c5_0 + p_20_4;
  assign t_r21_c5_6 = t_r21_c5_1 + p_20_6;
  assign t_r21_c5_7 = t_r21_c5_2 + t_r21_c5_3;
  assign t_r21_c5_8 = t_r21_c5_4 + p_22_4;
  assign t_r21_c5_9 = t_r21_c5_5 + t_r21_c5_6;
  assign t_r21_c5_10 = t_r21_c5_7 + t_r21_c5_8;
  assign t_r21_c5_11 = t_r21_c5_9 + t_r21_c5_10;
  assign t_r21_c5_12 = t_r21_c5_11 + p_22_6;
  assign out_21_5 = t_r21_c5_12 >> 4;

  assign t_r21_c6_0 = p_20_6 << 1;
  assign t_r21_c6_1 = p_21_5 << 1;
  assign t_r21_c6_2 = p_21_6 << 2;
  assign t_r21_c6_3 = p_21_7 << 1;
  assign t_r21_c6_4 = p_22_6 << 1;
  assign t_r21_c6_5 = t_r21_c6_0 + p_20_5;
  assign t_r21_c6_6 = t_r21_c6_1 + p_20_7;
  assign t_r21_c6_7 = t_r21_c6_2 + t_r21_c6_3;
  assign t_r21_c6_8 = t_r21_c6_4 + p_22_5;
  assign t_r21_c6_9 = t_r21_c6_5 + t_r21_c6_6;
  assign t_r21_c6_10 = t_r21_c6_7 + t_r21_c6_8;
  assign t_r21_c6_11 = t_r21_c6_9 + t_r21_c6_10;
  assign t_r21_c6_12 = t_r21_c6_11 + p_22_7;
  assign out_21_6 = t_r21_c6_12 >> 4;

  assign t_r21_c7_0 = p_20_7 << 1;
  assign t_r21_c7_1 = p_21_6 << 1;
  assign t_r21_c7_2 = p_21_7 << 2;
  assign t_r21_c7_3 = p_21_8 << 1;
  assign t_r21_c7_4 = p_22_7 << 1;
  assign t_r21_c7_5 = t_r21_c7_0 + p_20_6;
  assign t_r21_c7_6 = t_r21_c7_1 + p_20_8;
  assign t_r21_c7_7 = t_r21_c7_2 + t_r21_c7_3;
  assign t_r21_c7_8 = t_r21_c7_4 + p_22_6;
  assign t_r21_c7_9 = t_r21_c7_5 + t_r21_c7_6;
  assign t_r21_c7_10 = t_r21_c7_7 + t_r21_c7_8;
  assign t_r21_c7_11 = t_r21_c7_9 + t_r21_c7_10;
  assign t_r21_c7_12 = t_r21_c7_11 + p_22_8;
  assign out_21_7 = t_r21_c7_12 >> 4;

  assign t_r21_c8_0 = p_20_8 << 1;
  assign t_r21_c8_1 = p_21_7 << 1;
  assign t_r21_c8_2 = p_21_8 << 2;
  assign t_r21_c8_3 = p_21_9 << 1;
  assign t_r21_c8_4 = p_22_8 << 1;
  assign t_r21_c8_5 = t_r21_c8_0 + p_20_7;
  assign t_r21_c8_6 = t_r21_c8_1 + p_20_9;
  assign t_r21_c8_7 = t_r21_c8_2 + t_r21_c8_3;
  assign t_r21_c8_8 = t_r21_c8_4 + p_22_7;
  assign t_r21_c8_9 = t_r21_c8_5 + t_r21_c8_6;
  assign t_r21_c8_10 = t_r21_c8_7 + t_r21_c8_8;
  assign t_r21_c8_11 = t_r21_c8_9 + t_r21_c8_10;
  assign t_r21_c8_12 = t_r21_c8_11 + p_22_9;
  assign out_21_8 = t_r21_c8_12 >> 4;

  assign t_r21_c9_0 = p_20_9 << 1;
  assign t_r21_c9_1 = p_21_8 << 1;
  assign t_r21_c9_2 = p_21_9 << 2;
  assign t_r21_c9_3 = p_21_10 << 1;
  assign t_r21_c9_4 = p_22_9 << 1;
  assign t_r21_c9_5 = t_r21_c9_0 + p_20_8;
  assign t_r21_c9_6 = t_r21_c9_1 + p_20_10;
  assign t_r21_c9_7 = t_r21_c9_2 + t_r21_c9_3;
  assign t_r21_c9_8 = t_r21_c9_4 + p_22_8;
  assign t_r21_c9_9 = t_r21_c9_5 + t_r21_c9_6;
  assign t_r21_c9_10 = t_r21_c9_7 + t_r21_c9_8;
  assign t_r21_c9_11 = t_r21_c9_9 + t_r21_c9_10;
  assign t_r21_c9_12 = t_r21_c9_11 + p_22_10;
  assign out_21_9 = t_r21_c9_12 >> 4;

  assign t_r21_c10_0 = p_20_10 << 1;
  assign t_r21_c10_1 = p_21_9 << 1;
  assign t_r21_c10_2 = p_21_10 << 2;
  assign t_r21_c10_3 = p_21_11 << 1;
  assign t_r21_c10_4 = p_22_10 << 1;
  assign t_r21_c10_5 = t_r21_c10_0 + p_20_9;
  assign t_r21_c10_6 = t_r21_c10_1 + p_20_11;
  assign t_r21_c10_7 = t_r21_c10_2 + t_r21_c10_3;
  assign t_r21_c10_8 = t_r21_c10_4 + p_22_9;
  assign t_r21_c10_9 = t_r21_c10_5 + t_r21_c10_6;
  assign t_r21_c10_10 = t_r21_c10_7 + t_r21_c10_8;
  assign t_r21_c10_11 = t_r21_c10_9 + t_r21_c10_10;
  assign t_r21_c10_12 = t_r21_c10_11 + p_22_11;
  assign out_21_10 = t_r21_c10_12 >> 4;

  assign t_r21_c11_0 = p_20_11 << 1;
  assign t_r21_c11_1 = p_21_10 << 1;
  assign t_r21_c11_2 = p_21_11 << 2;
  assign t_r21_c11_3 = p_21_12 << 1;
  assign t_r21_c11_4 = p_22_11 << 1;
  assign t_r21_c11_5 = t_r21_c11_0 + p_20_10;
  assign t_r21_c11_6 = t_r21_c11_1 + p_20_12;
  assign t_r21_c11_7 = t_r21_c11_2 + t_r21_c11_3;
  assign t_r21_c11_8 = t_r21_c11_4 + p_22_10;
  assign t_r21_c11_9 = t_r21_c11_5 + t_r21_c11_6;
  assign t_r21_c11_10 = t_r21_c11_7 + t_r21_c11_8;
  assign t_r21_c11_11 = t_r21_c11_9 + t_r21_c11_10;
  assign t_r21_c11_12 = t_r21_c11_11 + p_22_12;
  assign out_21_11 = t_r21_c11_12 >> 4;

  assign t_r21_c12_0 = p_20_12 << 1;
  assign t_r21_c12_1 = p_21_11 << 1;
  assign t_r21_c12_2 = p_21_12 << 2;
  assign t_r21_c12_3 = p_21_13 << 1;
  assign t_r21_c12_4 = p_22_12 << 1;
  assign t_r21_c12_5 = t_r21_c12_0 + p_20_11;
  assign t_r21_c12_6 = t_r21_c12_1 + p_20_13;
  assign t_r21_c12_7 = t_r21_c12_2 + t_r21_c12_3;
  assign t_r21_c12_8 = t_r21_c12_4 + p_22_11;
  assign t_r21_c12_9 = t_r21_c12_5 + t_r21_c12_6;
  assign t_r21_c12_10 = t_r21_c12_7 + t_r21_c12_8;
  assign t_r21_c12_11 = t_r21_c12_9 + t_r21_c12_10;
  assign t_r21_c12_12 = t_r21_c12_11 + p_22_13;
  assign out_21_12 = t_r21_c12_12 >> 4;

  assign t_r21_c13_0 = p_20_13 << 1;
  assign t_r21_c13_1 = p_21_12 << 1;
  assign t_r21_c13_2 = p_21_13 << 2;
  assign t_r21_c13_3 = p_21_14 << 1;
  assign t_r21_c13_4 = p_22_13 << 1;
  assign t_r21_c13_5 = t_r21_c13_0 + p_20_12;
  assign t_r21_c13_6 = t_r21_c13_1 + p_20_14;
  assign t_r21_c13_7 = t_r21_c13_2 + t_r21_c13_3;
  assign t_r21_c13_8 = t_r21_c13_4 + p_22_12;
  assign t_r21_c13_9 = t_r21_c13_5 + t_r21_c13_6;
  assign t_r21_c13_10 = t_r21_c13_7 + t_r21_c13_8;
  assign t_r21_c13_11 = t_r21_c13_9 + t_r21_c13_10;
  assign t_r21_c13_12 = t_r21_c13_11 + p_22_14;
  assign out_21_13 = t_r21_c13_12 >> 4;

  assign t_r21_c14_0 = p_20_14 << 1;
  assign t_r21_c14_1 = p_21_13 << 1;
  assign t_r21_c14_2 = p_21_14 << 2;
  assign t_r21_c14_3 = p_21_15 << 1;
  assign t_r21_c14_4 = p_22_14 << 1;
  assign t_r21_c14_5 = t_r21_c14_0 + p_20_13;
  assign t_r21_c14_6 = t_r21_c14_1 + p_20_15;
  assign t_r21_c14_7 = t_r21_c14_2 + t_r21_c14_3;
  assign t_r21_c14_8 = t_r21_c14_4 + p_22_13;
  assign t_r21_c14_9 = t_r21_c14_5 + t_r21_c14_6;
  assign t_r21_c14_10 = t_r21_c14_7 + t_r21_c14_8;
  assign t_r21_c14_11 = t_r21_c14_9 + t_r21_c14_10;
  assign t_r21_c14_12 = t_r21_c14_11 + p_22_15;
  assign out_21_14 = t_r21_c14_12 >> 4;

  assign t_r21_c15_0 = p_20_15 << 1;
  assign t_r21_c15_1 = p_21_14 << 1;
  assign t_r21_c15_2 = p_21_15 << 2;
  assign t_r21_c15_3 = p_21_16 << 1;
  assign t_r21_c15_4 = p_22_15 << 1;
  assign t_r21_c15_5 = t_r21_c15_0 + p_20_14;
  assign t_r21_c15_6 = t_r21_c15_1 + p_20_16;
  assign t_r21_c15_7 = t_r21_c15_2 + t_r21_c15_3;
  assign t_r21_c15_8 = t_r21_c15_4 + p_22_14;
  assign t_r21_c15_9 = t_r21_c15_5 + t_r21_c15_6;
  assign t_r21_c15_10 = t_r21_c15_7 + t_r21_c15_8;
  assign t_r21_c15_11 = t_r21_c15_9 + t_r21_c15_10;
  assign t_r21_c15_12 = t_r21_c15_11 + p_22_16;
  assign out_21_15 = t_r21_c15_12 >> 4;

  assign t_r21_c16_0 = p_20_16 << 1;
  assign t_r21_c16_1 = p_21_15 << 1;
  assign t_r21_c16_2 = p_21_16 << 2;
  assign t_r21_c16_3 = p_21_17 << 1;
  assign t_r21_c16_4 = p_22_16 << 1;
  assign t_r21_c16_5 = t_r21_c16_0 + p_20_15;
  assign t_r21_c16_6 = t_r21_c16_1 + p_20_17;
  assign t_r21_c16_7 = t_r21_c16_2 + t_r21_c16_3;
  assign t_r21_c16_8 = t_r21_c16_4 + p_22_15;
  assign t_r21_c16_9 = t_r21_c16_5 + t_r21_c16_6;
  assign t_r21_c16_10 = t_r21_c16_7 + t_r21_c16_8;
  assign t_r21_c16_11 = t_r21_c16_9 + t_r21_c16_10;
  assign t_r21_c16_12 = t_r21_c16_11 + p_22_17;
  assign out_21_16 = t_r21_c16_12 >> 4;

  assign t_r21_c17_0 = p_20_17 << 1;
  assign t_r21_c17_1 = p_21_16 << 1;
  assign t_r21_c17_2 = p_21_17 << 2;
  assign t_r21_c17_3 = p_21_18 << 1;
  assign t_r21_c17_4 = p_22_17 << 1;
  assign t_r21_c17_5 = t_r21_c17_0 + p_20_16;
  assign t_r21_c17_6 = t_r21_c17_1 + p_20_18;
  assign t_r21_c17_7 = t_r21_c17_2 + t_r21_c17_3;
  assign t_r21_c17_8 = t_r21_c17_4 + p_22_16;
  assign t_r21_c17_9 = t_r21_c17_5 + t_r21_c17_6;
  assign t_r21_c17_10 = t_r21_c17_7 + t_r21_c17_8;
  assign t_r21_c17_11 = t_r21_c17_9 + t_r21_c17_10;
  assign t_r21_c17_12 = t_r21_c17_11 + p_22_18;
  assign out_21_17 = t_r21_c17_12 >> 4;

  assign t_r21_c18_0 = p_20_18 << 1;
  assign t_r21_c18_1 = p_21_17 << 1;
  assign t_r21_c18_2 = p_21_18 << 2;
  assign t_r21_c18_3 = p_21_19 << 1;
  assign t_r21_c18_4 = p_22_18 << 1;
  assign t_r21_c18_5 = t_r21_c18_0 + p_20_17;
  assign t_r21_c18_6 = t_r21_c18_1 + p_20_19;
  assign t_r21_c18_7 = t_r21_c18_2 + t_r21_c18_3;
  assign t_r21_c18_8 = t_r21_c18_4 + p_22_17;
  assign t_r21_c18_9 = t_r21_c18_5 + t_r21_c18_6;
  assign t_r21_c18_10 = t_r21_c18_7 + t_r21_c18_8;
  assign t_r21_c18_11 = t_r21_c18_9 + t_r21_c18_10;
  assign t_r21_c18_12 = t_r21_c18_11 + p_22_19;
  assign out_21_18 = t_r21_c18_12 >> 4;

  assign t_r21_c19_0 = p_20_19 << 1;
  assign t_r21_c19_1 = p_21_18 << 1;
  assign t_r21_c19_2 = p_21_19 << 2;
  assign t_r21_c19_3 = p_21_20 << 1;
  assign t_r21_c19_4 = p_22_19 << 1;
  assign t_r21_c19_5 = t_r21_c19_0 + p_20_18;
  assign t_r21_c19_6 = t_r21_c19_1 + p_20_20;
  assign t_r21_c19_7 = t_r21_c19_2 + t_r21_c19_3;
  assign t_r21_c19_8 = t_r21_c19_4 + p_22_18;
  assign t_r21_c19_9 = t_r21_c19_5 + t_r21_c19_6;
  assign t_r21_c19_10 = t_r21_c19_7 + t_r21_c19_8;
  assign t_r21_c19_11 = t_r21_c19_9 + t_r21_c19_10;
  assign t_r21_c19_12 = t_r21_c19_11 + p_22_20;
  assign out_21_19 = t_r21_c19_12 >> 4;

  assign t_r21_c20_0 = p_20_20 << 1;
  assign t_r21_c20_1 = p_21_19 << 1;
  assign t_r21_c20_2 = p_21_20 << 2;
  assign t_r21_c20_3 = p_21_21 << 1;
  assign t_r21_c20_4 = p_22_20 << 1;
  assign t_r21_c20_5 = t_r21_c20_0 + p_20_19;
  assign t_r21_c20_6 = t_r21_c20_1 + p_20_21;
  assign t_r21_c20_7 = t_r21_c20_2 + t_r21_c20_3;
  assign t_r21_c20_8 = t_r21_c20_4 + p_22_19;
  assign t_r21_c20_9 = t_r21_c20_5 + t_r21_c20_6;
  assign t_r21_c20_10 = t_r21_c20_7 + t_r21_c20_8;
  assign t_r21_c20_11 = t_r21_c20_9 + t_r21_c20_10;
  assign t_r21_c20_12 = t_r21_c20_11 + p_22_21;
  assign out_21_20 = t_r21_c20_12 >> 4;

  assign t_r21_c21_0 = p_20_21 << 1;
  assign t_r21_c21_1 = p_21_20 << 1;
  assign t_r21_c21_2 = p_21_21 << 2;
  assign t_r21_c21_3 = p_21_22 << 1;
  assign t_r21_c21_4 = p_22_21 << 1;
  assign t_r21_c21_5 = t_r21_c21_0 + p_20_20;
  assign t_r21_c21_6 = t_r21_c21_1 + p_20_22;
  assign t_r21_c21_7 = t_r21_c21_2 + t_r21_c21_3;
  assign t_r21_c21_8 = t_r21_c21_4 + p_22_20;
  assign t_r21_c21_9 = t_r21_c21_5 + t_r21_c21_6;
  assign t_r21_c21_10 = t_r21_c21_7 + t_r21_c21_8;
  assign t_r21_c21_11 = t_r21_c21_9 + t_r21_c21_10;
  assign t_r21_c21_12 = t_r21_c21_11 + p_22_22;
  assign out_21_21 = t_r21_c21_12 >> 4;

  assign t_r21_c22_0 = p_20_22 << 1;
  assign t_r21_c22_1 = p_21_21 << 1;
  assign t_r21_c22_2 = p_21_22 << 2;
  assign t_r21_c22_3 = p_21_23 << 1;
  assign t_r21_c22_4 = p_22_22 << 1;
  assign t_r21_c22_5 = t_r21_c22_0 + p_20_21;
  assign t_r21_c22_6 = t_r21_c22_1 + p_20_23;
  assign t_r21_c22_7 = t_r21_c22_2 + t_r21_c22_3;
  assign t_r21_c22_8 = t_r21_c22_4 + p_22_21;
  assign t_r21_c22_9 = t_r21_c22_5 + t_r21_c22_6;
  assign t_r21_c22_10 = t_r21_c22_7 + t_r21_c22_8;
  assign t_r21_c22_11 = t_r21_c22_9 + t_r21_c22_10;
  assign t_r21_c22_12 = t_r21_c22_11 + p_22_23;
  assign out_21_22 = t_r21_c22_12 >> 4;

  assign t_r21_c23_0 = p_20_23 << 1;
  assign t_r21_c23_1 = p_21_22 << 1;
  assign t_r21_c23_2 = p_21_23 << 2;
  assign t_r21_c23_3 = p_21_24 << 1;
  assign t_r21_c23_4 = p_22_23 << 1;
  assign t_r21_c23_5 = t_r21_c23_0 + p_20_22;
  assign t_r21_c23_6 = t_r21_c23_1 + p_20_24;
  assign t_r21_c23_7 = t_r21_c23_2 + t_r21_c23_3;
  assign t_r21_c23_8 = t_r21_c23_4 + p_22_22;
  assign t_r21_c23_9 = t_r21_c23_5 + t_r21_c23_6;
  assign t_r21_c23_10 = t_r21_c23_7 + t_r21_c23_8;
  assign t_r21_c23_11 = t_r21_c23_9 + t_r21_c23_10;
  assign t_r21_c23_12 = t_r21_c23_11 + p_22_24;
  assign out_21_23 = t_r21_c23_12 >> 4;

  assign t_r21_c24_0 = p_20_24 << 1;
  assign t_r21_c24_1 = p_21_23 << 1;
  assign t_r21_c24_2 = p_21_24 << 2;
  assign t_r21_c24_3 = p_21_25 << 1;
  assign t_r21_c24_4 = p_22_24 << 1;
  assign t_r21_c24_5 = t_r21_c24_0 + p_20_23;
  assign t_r21_c24_6 = t_r21_c24_1 + p_20_25;
  assign t_r21_c24_7 = t_r21_c24_2 + t_r21_c24_3;
  assign t_r21_c24_8 = t_r21_c24_4 + p_22_23;
  assign t_r21_c24_9 = t_r21_c24_5 + t_r21_c24_6;
  assign t_r21_c24_10 = t_r21_c24_7 + t_r21_c24_8;
  assign t_r21_c24_11 = t_r21_c24_9 + t_r21_c24_10;
  assign t_r21_c24_12 = t_r21_c24_11 + p_22_25;
  assign out_21_24 = t_r21_c24_12 >> 4;

  assign t_r21_c25_0 = p_20_25 << 1;
  assign t_r21_c25_1 = p_21_24 << 1;
  assign t_r21_c25_2 = p_21_25 << 2;
  assign t_r21_c25_3 = p_21_26 << 1;
  assign t_r21_c25_4 = p_22_25 << 1;
  assign t_r21_c25_5 = t_r21_c25_0 + p_20_24;
  assign t_r21_c25_6 = t_r21_c25_1 + p_20_26;
  assign t_r21_c25_7 = t_r21_c25_2 + t_r21_c25_3;
  assign t_r21_c25_8 = t_r21_c25_4 + p_22_24;
  assign t_r21_c25_9 = t_r21_c25_5 + t_r21_c25_6;
  assign t_r21_c25_10 = t_r21_c25_7 + t_r21_c25_8;
  assign t_r21_c25_11 = t_r21_c25_9 + t_r21_c25_10;
  assign t_r21_c25_12 = t_r21_c25_11 + p_22_26;
  assign out_21_25 = t_r21_c25_12 >> 4;

  assign t_r21_c26_0 = p_20_26 << 1;
  assign t_r21_c26_1 = p_21_25 << 1;
  assign t_r21_c26_2 = p_21_26 << 2;
  assign t_r21_c26_3 = p_21_27 << 1;
  assign t_r21_c26_4 = p_22_26 << 1;
  assign t_r21_c26_5 = t_r21_c26_0 + p_20_25;
  assign t_r21_c26_6 = t_r21_c26_1 + p_20_27;
  assign t_r21_c26_7 = t_r21_c26_2 + t_r21_c26_3;
  assign t_r21_c26_8 = t_r21_c26_4 + p_22_25;
  assign t_r21_c26_9 = t_r21_c26_5 + t_r21_c26_6;
  assign t_r21_c26_10 = t_r21_c26_7 + t_r21_c26_8;
  assign t_r21_c26_11 = t_r21_c26_9 + t_r21_c26_10;
  assign t_r21_c26_12 = t_r21_c26_11 + p_22_27;
  assign out_21_26 = t_r21_c26_12 >> 4;

  assign t_r21_c27_0 = p_20_27 << 1;
  assign t_r21_c27_1 = p_21_26 << 1;
  assign t_r21_c27_2 = p_21_27 << 2;
  assign t_r21_c27_3 = p_21_28 << 1;
  assign t_r21_c27_4 = p_22_27 << 1;
  assign t_r21_c27_5 = t_r21_c27_0 + p_20_26;
  assign t_r21_c27_6 = t_r21_c27_1 + p_20_28;
  assign t_r21_c27_7 = t_r21_c27_2 + t_r21_c27_3;
  assign t_r21_c27_8 = t_r21_c27_4 + p_22_26;
  assign t_r21_c27_9 = t_r21_c27_5 + t_r21_c27_6;
  assign t_r21_c27_10 = t_r21_c27_7 + t_r21_c27_8;
  assign t_r21_c27_11 = t_r21_c27_9 + t_r21_c27_10;
  assign t_r21_c27_12 = t_r21_c27_11 + p_22_28;
  assign out_21_27 = t_r21_c27_12 >> 4;

  assign t_r21_c28_0 = p_20_28 << 1;
  assign t_r21_c28_1 = p_21_27 << 1;
  assign t_r21_c28_2 = p_21_28 << 2;
  assign t_r21_c28_3 = p_21_29 << 1;
  assign t_r21_c28_4 = p_22_28 << 1;
  assign t_r21_c28_5 = t_r21_c28_0 + p_20_27;
  assign t_r21_c28_6 = t_r21_c28_1 + p_20_29;
  assign t_r21_c28_7 = t_r21_c28_2 + t_r21_c28_3;
  assign t_r21_c28_8 = t_r21_c28_4 + p_22_27;
  assign t_r21_c28_9 = t_r21_c28_5 + t_r21_c28_6;
  assign t_r21_c28_10 = t_r21_c28_7 + t_r21_c28_8;
  assign t_r21_c28_11 = t_r21_c28_9 + t_r21_c28_10;
  assign t_r21_c28_12 = t_r21_c28_11 + p_22_29;
  assign out_21_28 = t_r21_c28_12 >> 4;

  assign t_r21_c29_0 = p_20_29 << 1;
  assign t_r21_c29_1 = p_21_28 << 1;
  assign t_r21_c29_2 = p_21_29 << 2;
  assign t_r21_c29_3 = p_21_30 << 1;
  assign t_r21_c29_4 = p_22_29 << 1;
  assign t_r21_c29_5 = t_r21_c29_0 + p_20_28;
  assign t_r21_c29_6 = t_r21_c29_1 + p_20_30;
  assign t_r21_c29_7 = t_r21_c29_2 + t_r21_c29_3;
  assign t_r21_c29_8 = t_r21_c29_4 + p_22_28;
  assign t_r21_c29_9 = t_r21_c29_5 + t_r21_c29_6;
  assign t_r21_c29_10 = t_r21_c29_7 + t_r21_c29_8;
  assign t_r21_c29_11 = t_r21_c29_9 + t_r21_c29_10;
  assign t_r21_c29_12 = t_r21_c29_11 + p_22_30;
  assign out_21_29 = t_r21_c29_12 >> 4;

  assign t_r21_c30_0 = p_20_30 << 1;
  assign t_r21_c30_1 = p_21_29 << 1;
  assign t_r21_c30_2 = p_21_30 << 2;
  assign t_r21_c30_3 = p_21_31 << 1;
  assign t_r21_c30_4 = p_22_30 << 1;
  assign t_r21_c30_5 = t_r21_c30_0 + p_20_29;
  assign t_r21_c30_6 = t_r21_c30_1 + p_20_31;
  assign t_r21_c30_7 = t_r21_c30_2 + t_r21_c30_3;
  assign t_r21_c30_8 = t_r21_c30_4 + p_22_29;
  assign t_r21_c30_9 = t_r21_c30_5 + t_r21_c30_6;
  assign t_r21_c30_10 = t_r21_c30_7 + t_r21_c30_8;
  assign t_r21_c30_11 = t_r21_c30_9 + t_r21_c30_10;
  assign t_r21_c30_12 = t_r21_c30_11 + p_22_31;
  assign out_21_30 = t_r21_c30_12 >> 4;

  assign t_r21_c31_0 = p_20_31 << 1;
  assign t_r21_c31_1 = p_21_30 << 1;
  assign t_r21_c31_2 = p_21_31 << 2;
  assign t_r21_c31_3 = p_21_32 << 1;
  assign t_r21_c31_4 = p_22_31 << 1;
  assign t_r21_c31_5 = t_r21_c31_0 + p_20_30;
  assign t_r21_c31_6 = t_r21_c31_1 + p_20_32;
  assign t_r21_c31_7 = t_r21_c31_2 + t_r21_c31_3;
  assign t_r21_c31_8 = t_r21_c31_4 + p_22_30;
  assign t_r21_c31_9 = t_r21_c31_5 + t_r21_c31_6;
  assign t_r21_c31_10 = t_r21_c31_7 + t_r21_c31_8;
  assign t_r21_c31_11 = t_r21_c31_9 + t_r21_c31_10;
  assign t_r21_c31_12 = t_r21_c31_11 + p_22_32;
  assign out_21_31 = t_r21_c31_12 >> 4;

  assign t_r21_c32_0 = p_20_32 << 1;
  assign t_r21_c32_1 = p_21_31 << 1;
  assign t_r21_c32_2 = p_21_32 << 2;
  assign t_r21_c32_3 = p_21_33 << 1;
  assign t_r21_c32_4 = p_22_32 << 1;
  assign t_r21_c32_5 = t_r21_c32_0 + p_20_31;
  assign t_r21_c32_6 = t_r21_c32_1 + p_20_33;
  assign t_r21_c32_7 = t_r21_c32_2 + t_r21_c32_3;
  assign t_r21_c32_8 = t_r21_c32_4 + p_22_31;
  assign t_r21_c32_9 = t_r21_c32_5 + t_r21_c32_6;
  assign t_r21_c32_10 = t_r21_c32_7 + t_r21_c32_8;
  assign t_r21_c32_11 = t_r21_c32_9 + t_r21_c32_10;
  assign t_r21_c32_12 = t_r21_c32_11 + p_22_33;
  assign out_21_32 = t_r21_c32_12 >> 4;

  assign t_r21_c33_0 = p_20_33 << 1;
  assign t_r21_c33_1 = p_21_32 << 1;
  assign t_r21_c33_2 = p_21_33 << 2;
  assign t_r21_c33_3 = p_21_34 << 1;
  assign t_r21_c33_4 = p_22_33 << 1;
  assign t_r21_c33_5 = t_r21_c33_0 + p_20_32;
  assign t_r21_c33_6 = t_r21_c33_1 + p_20_34;
  assign t_r21_c33_7 = t_r21_c33_2 + t_r21_c33_3;
  assign t_r21_c33_8 = t_r21_c33_4 + p_22_32;
  assign t_r21_c33_9 = t_r21_c33_5 + t_r21_c33_6;
  assign t_r21_c33_10 = t_r21_c33_7 + t_r21_c33_8;
  assign t_r21_c33_11 = t_r21_c33_9 + t_r21_c33_10;
  assign t_r21_c33_12 = t_r21_c33_11 + p_22_34;
  assign out_21_33 = t_r21_c33_12 >> 4;

  assign t_r21_c34_0 = p_20_34 << 1;
  assign t_r21_c34_1 = p_21_33 << 1;
  assign t_r21_c34_2 = p_21_34 << 2;
  assign t_r21_c34_3 = p_21_35 << 1;
  assign t_r21_c34_4 = p_22_34 << 1;
  assign t_r21_c34_5 = t_r21_c34_0 + p_20_33;
  assign t_r21_c34_6 = t_r21_c34_1 + p_20_35;
  assign t_r21_c34_7 = t_r21_c34_2 + t_r21_c34_3;
  assign t_r21_c34_8 = t_r21_c34_4 + p_22_33;
  assign t_r21_c34_9 = t_r21_c34_5 + t_r21_c34_6;
  assign t_r21_c34_10 = t_r21_c34_7 + t_r21_c34_8;
  assign t_r21_c34_11 = t_r21_c34_9 + t_r21_c34_10;
  assign t_r21_c34_12 = t_r21_c34_11 + p_22_35;
  assign out_21_34 = t_r21_c34_12 >> 4;

  assign t_r21_c35_0 = p_20_35 << 1;
  assign t_r21_c35_1 = p_21_34 << 1;
  assign t_r21_c35_2 = p_21_35 << 2;
  assign t_r21_c35_3 = p_21_36 << 1;
  assign t_r21_c35_4 = p_22_35 << 1;
  assign t_r21_c35_5 = t_r21_c35_0 + p_20_34;
  assign t_r21_c35_6 = t_r21_c35_1 + p_20_36;
  assign t_r21_c35_7 = t_r21_c35_2 + t_r21_c35_3;
  assign t_r21_c35_8 = t_r21_c35_4 + p_22_34;
  assign t_r21_c35_9 = t_r21_c35_5 + t_r21_c35_6;
  assign t_r21_c35_10 = t_r21_c35_7 + t_r21_c35_8;
  assign t_r21_c35_11 = t_r21_c35_9 + t_r21_c35_10;
  assign t_r21_c35_12 = t_r21_c35_11 + p_22_36;
  assign out_21_35 = t_r21_c35_12 >> 4;

  assign t_r21_c36_0 = p_20_36 << 1;
  assign t_r21_c36_1 = p_21_35 << 1;
  assign t_r21_c36_2 = p_21_36 << 2;
  assign t_r21_c36_3 = p_21_37 << 1;
  assign t_r21_c36_4 = p_22_36 << 1;
  assign t_r21_c36_5 = t_r21_c36_0 + p_20_35;
  assign t_r21_c36_6 = t_r21_c36_1 + p_20_37;
  assign t_r21_c36_7 = t_r21_c36_2 + t_r21_c36_3;
  assign t_r21_c36_8 = t_r21_c36_4 + p_22_35;
  assign t_r21_c36_9 = t_r21_c36_5 + t_r21_c36_6;
  assign t_r21_c36_10 = t_r21_c36_7 + t_r21_c36_8;
  assign t_r21_c36_11 = t_r21_c36_9 + t_r21_c36_10;
  assign t_r21_c36_12 = t_r21_c36_11 + p_22_37;
  assign out_21_36 = t_r21_c36_12 >> 4;

  assign t_r21_c37_0 = p_20_37 << 1;
  assign t_r21_c37_1 = p_21_36 << 1;
  assign t_r21_c37_2 = p_21_37 << 2;
  assign t_r21_c37_3 = p_21_38 << 1;
  assign t_r21_c37_4 = p_22_37 << 1;
  assign t_r21_c37_5 = t_r21_c37_0 + p_20_36;
  assign t_r21_c37_6 = t_r21_c37_1 + p_20_38;
  assign t_r21_c37_7 = t_r21_c37_2 + t_r21_c37_3;
  assign t_r21_c37_8 = t_r21_c37_4 + p_22_36;
  assign t_r21_c37_9 = t_r21_c37_5 + t_r21_c37_6;
  assign t_r21_c37_10 = t_r21_c37_7 + t_r21_c37_8;
  assign t_r21_c37_11 = t_r21_c37_9 + t_r21_c37_10;
  assign t_r21_c37_12 = t_r21_c37_11 + p_22_38;
  assign out_21_37 = t_r21_c37_12 >> 4;

  assign t_r21_c38_0 = p_20_38 << 1;
  assign t_r21_c38_1 = p_21_37 << 1;
  assign t_r21_c38_2 = p_21_38 << 2;
  assign t_r21_c38_3 = p_21_39 << 1;
  assign t_r21_c38_4 = p_22_38 << 1;
  assign t_r21_c38_5 = t_r21_c38_0 + p_20_37;
  assign t_r21_c38_6 = t_r21_c38_1 + p_20_39;
  assign t_r21_c38_7 = t_r21_c38_2 + t_r21_c38_3;
  assign t_r21_c38_8 = t_r21_c38_4 + p_22_37;
  assign t_r21_c38_9 = t_r21_c38_5 + t_r21_c38_6;
  assign t_r21_c38_10 = t_r21_c38_7 + t_r21_c38_8;
  assign t_r21_c38_11 = t_r21_c38_9 + t_r21_c38_10;
  assign t_r21_c38_12 = t_r21_c38_11 + p_22_39;
  assign out_21_38 = t_r21_c38_12 >> 4;

  assign t_r21_c39_0 = p_20_39 << 1;
  assign t_r21_c39_1 = p_21_38 << 1;
  assign t_r21_c39_2 = p_21_39 << 2;
  assign t_r21_c39_3 = p_21_40 << 1;
  assign t_r21_c39_4 = p_22_39 << 1;
  assign t_r21_c39_5 = t_r21_c39_0 + p_20_38;
  assign t_r21_c39_6 = t_r21_c39_1 + p_20_40;
  assign t_r21_c39_7 = t_r21_c39_2 + t_r21_c39_3;
  assign t_r21_c39_8 = t_r21_c39_4 + p_22_38;
  assign t_r21_c39_9 = t_r21_c39_5 + t_r21_c39_6;
  assign t_r21_c39_10 = t_r21_c39_7 + t_r21_c39_8;
  assign t_r21_c39_11 = t_r21_c39_9 + t_r21_c39_10;
  assign t_r21_c39_12 = t_r21_c39_11 + p_22_40;
  assign out_21_39 = t_r21_c39_12 >> 4;

  assign t_r21_c40_0 = p_20_40 << 1;
  assign t_r21_c40_1 = p_21_39 << 1;
  assign t_r21_c40_2 = p_21_40 << 2;
  assign t_r21_c40_3 = p_21_41 << 1;
  assign t_r21_c40_4 = p_22_40 << 1;
  assign t_r21_c40_5 = t_r21_c40_0 + p_20_39;
  assign t_r21_c40_6 = t_r21_c40_1 + p_20_41;
  assign t_r21_c40_7 = t_r21_c40_2 + t_r21_c40_3;
  assign t_r21_c40_8 = t_r21_c40_4 + p_22_39;
  assign t_r21_c40_9 = t_r21_c40_5 + t_r21_c40_6;
  assign t_r21_c40_10 = t_r21_c40_7 + t_r21_c40_8;
  assign t_r21_c40_11 = t_r21_c40_9 + t_r21_c40_10;
  assign t_r21_c40_12 = t_r21_c40_11 + p_22_41;
  assign out_21_40 = t_r21_c40_12 >> 4;

  assign t_r21_c41_0 = p_20_41 << 1;
  assign t_r21_c41_1 = p_21_40 << 1;
  assign t_r21_c41_2 = p_21_41 << 2;
  assign t_r21_c41_3 = p_21_42 << 1;
  assign t_r21_c41_4 = p_22_41 << 1;
  assign t_r21_c41_5 = t_r21_c41_0 + p_20_40;
  assign t_r21_c41_6 = t_r21_c41_1 + p_20_42;
  assign t_r21_c41_7 = t_r21_c41_2 + t_r21_c41_3;
  assign t_r21_c41_8 = t_r21_c41_4 + p_22_40;
  assign t_r21_c41_9 = t_r21_c41_5 + t_r21_c41_6;
  assign t_r21_c41_10 = t_r21_c41_7 + t_r21_c41_8;
  assign t_r21_c41_11 = t_r21_c41_9 + t_r21_c41_10;
  assign t_r21_c41_12 = t_r21_c41_11 + p_22_42;
  assign out_21_41 = t_r21_c41_12 >> 4;

  assign t_r21_c42_0 = p_20_42 << 1;
  assign t_r21_c42_1 = p_21_41 << 1;
  assign t_r21_c42_2 = p_21_42 << 2;
  assign t_r21_c42_3 = p_21_43 << 1;
  assign t_r21_c42_4 = p_22_42 << 1;
  assign t_r21_c42_5 = t_r21_c42_0 + p_20_41;
  assign t_r21_c42_6 = t_r21_c42_1 + p_20_43;
  assign t_r21_c42_7 = t_r21_c42_2 + t_r21_c42_3;
  assign t_r21_c42_8 = t_r21_c42_4 + p_22_41;
  assign t_r21_c42_9 = t_r21_c42_5 + t_r21_c42_6;
  assign t_r21_c42_10 = t_r21_c42_7 + t_r21_c42_8;
  assign t_r21_c42_11 = t_r21_c42_9 + t_r21_c42_10;
  assign t_r21_c42_12 = t_r21_c42_11 + p_22_43;
  assign out_21_42 = t_r21_c42_12 >> 4;

  assign t_r21_c43_0 = p_20_43 << 1;
  assign t_r21_c43_1 = p_21_42 << 1;
  assign t_r21_c43_2 = p_21_43 << 2;
  assign t_r21_c43_3 = p_21_44 << 1;
  assign t_r21_c43_4 = p_22_43 << 1;
  assign t_r21_c43_5 = t_r21_c43_0 + p_20_42;
  assign t_r21_c43_6 = t_r21_c43_1 + p_20_44;
  assign t_r21_c43_7 = t_r21_c43_2 + t_r21_c43_3;
  assign t_r21_c43_8 = t_r21_c43_4 + p_22_42;
  assign t_r21_c43_9 = t_r21_c43_5 + t_r21_c43_6;
  assign t_r21_c43_10 = t_r21_c43_7 + t_r21_c43_8;
  assign t_r21_c43_11 = t_r21_c43_9 + t_r21_c43_10;
  assign t_r21_c43_12 = t_r21_c43_11 + p_22_44;
  assign out_21_43 = t_r21_c43_12 >> 4;

  assign t_r21_c44_0 = p_20_44 << 1;
  assign t_r21_c44_1 = p_21_43 << 1;
  assign t_r21_c44_2 = p_21_44 << 2;
  assign t_r21_c44_3 = p_21_45 << 1;
  assign t_r21_c44_4 = p_22_44 << 1;
  assign t_r21_c44_5 = t_r21_c44_0 + p_20_43;
  assign t_r21_c44_6 = t_r21_c44_1 + p_20_45;
  assign t_r21_c44_7 = t_r21_c44_2 + t_r21_c44_3;
  assign t_r21_c44_8 = t_r21_c44_4 + p_22_43;
  assign t_r21_c44_9 = t_r21_c44_5 + t_r21_c44_6;
  assign t_r21_c44_10 = t_r21_c44_7 + t_r21_c44_8;
  assign t_r21_c44_11 = t_r21_c44_9 + t_r21_c44_10;
  assign t_r21_c44_12 = t_r21_c44_11 + p_22_45;
  assign out_21_44 = t_r21_c44_12 >> 4;

  assign t_r21_c45_0 = p_20_45 << 1;
  assign t_r21_c45_1 = p_21_44 << 1;
  assign t_r21_c45_2 = p_21_45 << 2;
  assign t_r21_c45_3 = p_21_46 << 1;
  assign t_r21_c45_4 = p_22_45 << 1;
  assign t_r21_c45_5 = t_r21_c45_0 + p_20_44;
  assign t_r21_c45_6 = t_r21_c45_1 + p_20_46;
  assign t_r21_c45_7 = t_r21_c45_2 + t_r21_c45_3;
  assign t_r21_c45_8 = t_r21_c45_4 + p_22_44;
  assign t_r21_c45_9 = t_r21_c45_5 + t_r21_c45_6;
  assign t_r21_c45_10 = t_r21_c45_7 + t_r21_c45_8;
  assign t_r21_c45_11 = t_r21_c45_9 + t_r21_c45_10;
  assign t_r21_c45_12 = t_r21_c45_11 + p_22_46;
  assign out_21_45 = t_r21_c45_12 >> 4;

  assign t_r21_c46_0 = p_20_46 << 1;
  assign t_r21_c46_1 = p_21_45 << 1;
  assign t_r21_c46_2 = p_21_46 << 2;
  assign t_r21_c46_3 = p_21_47 << 1;
  assign t_r21_c46_4 = p_22_46 << 1;
  assign t_r21_c46_5 = t_r21_c46_0 + p_20_45;
  assign t_r21_c46_6 = t_r21_c46_1 + p_20_47;
  assign t_r21_c46_7 = t_r21_c46_2 + t_r21_c46_3;
  assign t_r21_c46_8 = t_r21_c46_4 + p_22_45;
  assign t_r21_c46_9 = t_r21_c46_5 + t_r21_c46_6;
  assign t_r21_c46_10 = t_r21_c46_7 + t_r21_c46_8;
  assign t_r21_c46_11 = t_r21_c46_9 + t_r21_c46_10;
  assign t_r21_c46_12 = t_r21_c46_11 + p_22_47;
  assign out_21_46 = t_r21_c46_12 >> 4;

  assign t_r21_c47_0 = p_20_47 << 1;
  assign t_r21_c47_1 = p_21_46 << 1;
  assign t_r21_c47_2 = p_21_47 << 2;
  assign t_r21_c47_3 = p_21_48 << 1;
  assign t_r21_c47_4 = p_22_47 << 1;
  assign t_r21_c47_5 = t_r21_c47_0 + p_20_46;
  assign t_r21_c47_6 = t_r21_c47_1 + p_20_48;
  assign t_r21_c47_7 = t_r21_c47_2 + t_r21_c47_3;
  assign t_r21_c47_8 = t_r21_c47_4 + p_22_46;
  assign t_r21_c47_9 = t_r21_c47_5 + t_r21_c47_6;
  assign t_r21_c47_10 = t_r21_c47_7 + t_r21_c47_8;
  assign t_r21_c47_11 = t_r21_c47_9 + t_r21_c47_10;
  assign t_r21_c47_12 = t_r21_c47_11 + p_22_48;
  assign out_21_47 = t_r21_c47_12 >> 4;

  assign t_r21_c48_0 = p_20_48 << 1;
  assign t_r21_c48_1 = p_21_47 << 1;
  assign t_r21_c48_2 = p_21_48 << 2;
  assign t_r21_c48_3 = p_21_49 << 1;
  assign t_r21_c48_4 = p_22_48 << 1;
  assign t_r21_c48_5 = t_r21_c48_0 + p_20_47;
  assign t_r21_c48_6 = t_r21_c48_1 + p_20_49;
  assign t_r21_c48_7 = t_r21_c48_2 + t_r21_c48_3;
  assign t_r21_c48_8 = t_r21_c48_4 + p_22_47;
  assign t_r21_c48_9 = t_r21_c48_5 + t_r21_c48_6;
  assign t_r21_c48_10 = t_r21_c48_7 + t_r21_c48_8;
  assign t_r21_c48_11 = t_r21_c48_9 + t_r21_c48_10;
  assign t_r21_c48_12 = t_r21_c48_11 + p_22_49;
  assign out_21_48 = t_r21_c48_12 >> 4;

  assign t_r21_c49_0 = p_20_49 << 1;
  assign t_r21_c49_1 = p_21_48 << 1;
  assign t_r21_c49_2 = p_21_49 << 2;
  assign t_r21_c49_3 = p_21_50 << 1;
  assign t_r21_c49_4 = p_22_49 << 1;
  assign t_r21_c49_5 = t_r21_c49_0 + p_20_48;
  assign t_r21_c49_6 = t_r21_c49_1 + p_20_50;
  assign t_r21_c49_7 = t_r21_c49_2 + t_r21_c49_3;
  assign t_r21_c49_8 = t_r21_c49_4 + p_22_48;
  assign t_r21_c49_9 = t_r21_c49_5 + t_r21_c49_6;
  assign t_r21_c49_10 = t_r21_c49_7 + t_r21_c49_8;
  assign t_r21_c49_11 = t_r21_c49_9 + t_r21_c49_10;
  assign t_r21_c49_12 = t_r21_c49_11 + p_22_50;
  assign out_21_49 = t_r21_c49_12 >> 4;

  assign t_r21_c50_0 = p_20_50 << 1;
  assign t_r21_c50_1 = p_21_49 << 1;
  assign t_r21_c50_2 = p_21_50 << 2;
  assign t_r21_c50_3 = p_21_51 << 1;
  assign t_r21_c50_4 = p_22_50 << 1;
  assign t_r21_c50_5 = t_r21_c50_0 + p_20_49;
  assign t_r21_c50_6 = t_r21_c50_1 + p_20_51;
  assign t_r21_c50_7 = t_r21_c50_2 + t_r21_c50_3;
  assign t_r21_c50_8 = t_r21_c50_4 + p_22_49;
  assign t_r21_c50_9 = t_r21_c50_5 + t_r21_c50_6;
  assign t_r21_c50_10 = t_r21_c50_7 + t_r21_c50_8;
  assign t_r21_c50_11 = t_r21_c50_9 + t_r21_c50_10;
  assign t_r21_c50_12 = t_r21_c50_11 + p_22_51;
  assign out_21_50 = t_r21_c50_12 >> 4;

  assign t_r21_c51_0 = p_20_51 << 1;
  assign t_r21_c51_1 = p_21_50 << 1;
  assign t_r21_c51_2 = p_21_51 << 2;
  assign t_r21_c51_3 = p_21_52 << 1;
  assign t_r21_c51_4 = p_22_51 << 1;
  assign t_r21_c51_5 = t_r21_c51_0 + p_20_50;
  assign t_r21_c51_6 = t_r21_c51_1 + p_20_52;
  assign t_r21_c51_7 = t_r21_c51_2 + t_r21_c51_3;
  assign t_r21_c51_8 = t_r21_c51_4 + p_22_50;
  assign t_r21_c51_9 = t_r21_c51_5 + t_r21_c51_6;
  assign t_r21_c51_10 = t_r21_c51_7 + t_r21_c51_8;
  assign t_r21_c51_11 = t_r21_c51_9 + t_r21_c51_10;
  assign t_r21_c51_12 = t_r21_c51_11 + p_22_52;
  assign out_21_51 = t_r21_c51_12 >> 4;

  assign t_r21_c52_0 = p_20_52 << 1;
  assign t_r21_c52_1 = p_21_51 << 1;
  assign t_r21_c52_2 = p_21_52 << 2;
  assign t_r21_c52_3 = p_21_53 << 1;
  assign t_r21_c52_4 = p_22_52 << 1;
  assign t_r21_c52_5 = t_r21_c52_0 + p_20_51;
  assign t_r21_c52_6 = t_r21_c52_1 + p_20_53;
  assign t_r21_c52_7 = t_r21_c52_2 + t_r21_c52_3;
  assign t_r21_c52_8 = t_r21_c52_4 + p_22_51;
  assign t_r21_c52_9 = t_r21_c52_5 + t_r21_c52_6;
  assign t_r21_c52_10 = t_r21_c52_7 + t_r21_c52_8;
  assign t_r21_c52_11 = t_r21_c52_9 + t_r21_c52_10;
  assign t_r21_c52_12 = t_r21_c52_11 + p_22_53;
  assign out_21_52 = t_r21_c52_12 >> 4;

  assign t_r21_c53_0 = p_20_53 << 1;
  assign t_r21_c53_1 = p_21_52 << 1;
  assign t_r21_c53_2 = p_21_53 << 2;
  assign t_r21_c53_3 = p_21_54 << 1;
  assign t_r21_c53_4 = p_22_53 << 1;
  assign t_r21_c53_5 = t_r21_c53_0 + p_20_52;
  assign t_r21_c53_6 = t_r21_c53_1 + p_20_54;
  assign t_r21_c53_7 = t_r21_c53_2 + t_r21_c53_3;
  assign t_r21_c53_8 = t_r21_c53_4 + p_22_52;
  assign t_r21_c53_9 = t_r21_c53_5 + t_r21_c53_6;
  assign t_r21_c53_10 = t_r21_c53_7 + t_r21_c53_8;
  assign t_r21_c53_11 = t_r21_c53_9 + t_r21_c53_10;
  assign t_r21_c53_12 = t_r21_c53_11 + p_22_54;
  assign out_21_53 = t_r21_c53_12 >> 4;

  assign t_r21_c54_0 = p_20_54 << 1;
  assign t_r21_c54_1 = p_21_53 << 1;
  assign t_r21_c54_2 = p_21_54 << 2;
  assign t_r21_c54_3 = p_21_55 << 1;
  assign t_r21_c54_4 = p_22_54 << 1;
  assign t_r21_c54_5 = t_r21_c54_0 + p_20_53;
  assign t_r21_c54_6 = t_r21_c54_1 + p_20_55;
  assign t_r21_c54_7 = t_r21_c54_2 + t_r21_c54_3;
  assign t_r21_c54_8 = t_r21_c54_4 + p_22_53;
  assign t_r21_c54_9 = t_r21_c54_5 + t_r21_c54_6;
  assign t_r21_c54_10 = t_r21_c54_7 + t_r21_c54_8;
  assign t_r21_c54_11 = t_r21_c54_9 + t_r21_c54_10;
  assign t_r21_c54_12 = t_r21_c54_11 + p_22_55;
  assign out_21_54 = t_r21_c54_12 >> 4;

  assign t_r21_c55_0 = p_20_55 << 1;
  assign t_r21_c55_1 = p_21_54 << 1;
  assign t_r21_c55_2 = p_21_55 << 2;
  assign t_r21_c55_3 = p_21_56 << 1;
  assign t_r21_c55_4 = p_22_55 << 1;
  assign t_r21_c55_5 = t_r21_c55_0 + p_20_54;
  assign t_r21_c55_6 = t_r21_c55_1 + p_20_56;
  assign t_r21_c55_7 = t_r21_c55_2 + t_r21_c55_3;
  assign t_r21_c55_8 = t_r21_c55_4 + p_22_54;
  assign t_r21_c55_9 = t_r21_c55_5 + t_r21_c55_6;
  assign t_r21_c55_10 = t_r21_c55_7 + t_r21_c55_8;
  assign t_r21_c55_11 = t_r21_c55_9 + t_r21_c55_10;
  assign t_r21_c55_12 = t_r21_c55_11 + p_22_56;
  assign out_21_55 = t_r21_c55_12 >> 4;

  assign t_r21_c56_0 = p_20_56 << 1;
  assign t_r21_c56_1 = p_21_55 << 1;
  assign t_r21_c56_2 = p_21_56 << 2;
  assign t_r21_c56_3 = p_21_57 << 1;
  assign t_r21_c56_4 = p_22_56 << 1;
  assign t_r21_c56_5 = t_r21_c56_0 + p_20_55;
  assign t_r21_c56_6 = t_r21_c56_1 + p_20_57;
  assign t_r21_c56_7 = t_r21_c56_2 + t_r21_c56_3;
  assign t_r21_c56_8 = t_r21_c56_4 + p_22_55;
  assign t_r21_c56_9 = t_r21_c56_5 + t_r21_c56_6;
  assign t_r21_c56_10 = t_r21_c56_7 + t_r21_c56_8;
  assign t_r21_c56_11 = t_r21_c56_9 + t_r21_c56_10;
  assign t_r21_c56_12 = t_r21_c56_11 + p_22_57;
  assign out_21_56 = t_r21_c56_12 >> 4;

  assign t_r21_c57_0 = p_20_57 << 1;
  assign t_r21_c57_1 = p_21_56 << 1;
  assign t_r21_c57_2 = p_21_57 << 2;
  assign t_r21_c57_3 = p_21_58 << 1;
  assign t_r21_c57_4 = p_22_57 << 1;
  assign t_r21_c57_5 = t_r21_c57_0 + p_20_56;
  assign t_r21_c57_6 = t_r21_c57_1 + p_20_58;
  assign t_r21_c57_7 = t_r21_c57_2 + t_r21_c57_3;
  assign t_r21_c57_8 = t_r21_c57_4 + p_22_56;
  assign t_r21_c57_9 = t_r21_c57_5 + t_r21_c57_6;
  assign t_r21_c57_10 = t_r21_c57_7 + t_r21_c57_8;
  assign t_r21_c57_11 = t_r21_c57_9 + t_r21_c57_10;
  assign t_r21_c57_12 = t_r21_c57_11 + p_22_58;
  assign out_21_57 = t_r21_c57_12 >> 4;

  assign t_r21_c58_0 = p_20_58 << 1;
  assign t_r21_c58_1 = p_21_57 << 1;
  assign t_r21_c58_2 = p_21_58 << 2;
  assign t_r21_c58_3 = p_21_59 << 1;
  assign t_r21_c58_4 = p_22_58 << 1;
  assign t_r21_c58_5 = t_r21_c58_0 + p_20_57;
  assign t_r21_c58_6 = t_r21_c58_1 + p_20_59;
  assign t_r21_c58_7 = t_r21_c58_2 + t_r21_c58_3;
  assign t_r21_c58_8 = t_r21_c58_4 + p_22_57;
  assign t_r21_c58_9 = t_r21_c58_5 + t_r21_c58_6;
  assign t_r21_c58_10 = t_r21_c58_7 + t_r21_c58_8;
  assign t_r21_c58_11 = t_r21_c58_9 + t_r21_c58_10;
  assign t_r21_c58_12 = t_r21_c58_11 + p_22_59;
  assign out_21_58 = t_r21_c58_12 >> 4;

  assign t_r21_c59_0 = p_20_59 << 1;
  assign t_r21_c59_1 = p_21_58 << 1;
  assign t_r21_c59_2 = p_21_59 << 2;
  assign t_r21_c59_3 = p_21_60 << 1;
  assign t_r21_c59_4 = p_22_59 << 1;
  assign t_r21_c59_5 = t_r21_c59_0 + p_20_58;
  assign t_r21_c59_6 = t_r21_c59_1 + p_20_60;
  assign t_r21_c59_7 = t_r21_c59_2 + t_r21_c59_3;
  assign t_r21_c59_8 = t_r21_c59_4 + p_22_58;
  assign t_r21_c59_9 = t_r21_c59_5 + t_r21_c59_6;
  assign t_r21_c59_10 = t_r21_c59_7 + t_r21_c59_8;
  assign t_r21_c59_11 = t_r21_c59_9 + t_r21_c59_10;
  assign t_r21_c59_12 = t_r21_c59_11 + p_22_60;
  assign out_21_59 = t_r21_c59_12 >> 4;

  assign t_r21_c60_0 = p_20_60 << 1;
  assign t_r21_c60_1 = p_21_59 << 1;
  assign t_r21_c60_2 = p_21_60 << 2;
  assign t_r21_c60_3 = p_21_61 << 1;
  assign t_r21_c60_4 = p_22_60 << 1;
  assign t_r21_c60_5 = t_r21_c60_0 + p_20_59;
  assign t_r21_c60_6 = t_r21_c60_1 + p_20_61;
  assign t_r21_c60_7 = t_r21_c60_2 + t_r21_c60_3;
  assign t_r21_c60_8 = t_r21_c60_4 + p_22_59;
  assign t_r21_c60_9 = t_r21_c60_5 + t_r21_c60_6;
  assign t_r21_c60_10 = t_r21_c60_7 + t_r21_c60_8;
  assign t_r21_c60_11 = t_r21_c60_9 + t_r21_c60_10;
  assign t_r21_c60_12 = t_r21_c60_11 + p_22_61;
  assign out_21_60 = t_r21_c60_12 >> 4;

  assign t_r21_c61_0 = p_20_61 << 1;
  assign t_r21_c61_1 = p_21_60 << 1;
  assign t_r21_c61_2 = p_21_61 << 2;
  assign t_r21_c61_3 = p_21_62 << 1;
  assign t_r21_c61_4 = p_22_61 << 1;
  assign t_r21_c61_5 = t_r21_c61_0 + p_20_60;
  assign t_r21_c61_6 = t_r21_c61_1 + p_20_62;
  assign t_r21_c61_7 = t_r21_c61_2 + t_r21_c61_3;
  assign t_r21_c61_8 = t_r21_c61_4 + p_22_60;
  assign t_r21_c61_9 = t_r21_c61_5 + t_r21_c61_6;
  assign t_r21_c61_10 = t_r21_c61_7 + t_r21_c61_8;
  assign t_r21_c61_11 = t_r21_c61_9 + t_r21_c61_10;
  assign t_r21_c61_12 = t_r21_c61_11 + p_22_62;
  assign out_21_61 = t_r21_c61_12 >> 4;

  assign t_r21_c62_0 = p_20_62 << 1;
  assign t_r21_c62_1 = p_21_61 << 1;
  assign t_r21_c62_2 = p_21_62 << 2;
  assign t_r21_c62_3 = p_21_63 << 1;
  assign t_r21_c62_4 = p_22_62 << 1;
  assign t_r21_c62_5 = t_r21_c62_0 + p_20_61;
  assign t_r21_c62_6 = t_r21_c62_1 + p_20_63;
  assign t_r21_c62_7 = t_r21_c62_2 + t_r21_c62_3;
  assign t_r21_c62_8 = t_r21_c62_4 + p_22_61;
  assign t_r21_c62_9 = t_r21_c62_5 + t_r21_c62_6;
  assign t_r21_c62_10 = t_r21_c62_7 + t_r21_c62_8;
  assign t_r21_c62_11 = t_r21_c62_9 + t_r21_c62_10;
  assign t_r21_c62_12 = t_r21_c62_11 + p_22_63;
  assign out_21_62 = t_r21_c62_12 >> 4;

  assign t_r21_c63_0 = p_20_63 << 1;
  assign t_r21_c63_1 = p_21_62 << 1;
  assign t_r21_c63_2 = p_21_63 << 2;
  assign t_r21_c63_3 = p_21_64 << 1;
  assign t_r21_c63_4 = p_22_63 << 1;
  assign t_r21_c63_5 = t_r21_c63_0 + p_20_62;
  assign t_r21_c63_6 = t_r21_c63_1 + p_20_64;
  assign t_r21_c63_7 = t_r21_c63_2 + t_r21_c63_3;
  assign t_r21_c63_8 = t_r21_c63_4 + p_22_62;
  assign t_r21_c63_9 = t_r21_c63_5 + t_r21_c63_6;
  assign t_r21_c63_10 = t_r21_c63_7 + t_r21_c63_8;
  assign t_r21_c63_11 = t_r21_c63_9 + t_r21_c63_10;
  assign t_r21_c63_12 = t_r21_c63_11 + p_22_64;
  assign out_21_63 = t_r21_c63_12 >> 4;

  assign t_r21_c64_0 = p_20_64 << 1;
  assign t_r21_c64_1 = p_21_63 << 1;
  assign t_r21_c64_2 = p_21_64 << 2;
  assign t_r21_c64_3 = p_21_65 << 1;
  assign t_r21_c64_4 = p_22_64 << 1;
  assign t_r21_c64_5 = t_r21_c64_0 + p_20_63;
  assign t_r21_c64_6 = t_r21_c64_1 + p_20_65;
  assign t_r21_c64_7 = t_r21_c64_2 + t_r21_c64_3;
  assign t_r21_c64_8 = t_r21_c64_4 + p_22_63;
  assign t_r21_c64_9 = t_r21_c64_5 + t_r21_c64_6;
  assign t_r21_c64_10 = t_r21_c64_7 + t_r21_c64_8;
  assign t_r21_c64_11 = t_r21_c64_9 + t_r21_c64_10;
  assign t_r21_c64_12 = t_r21_c64_11 + p_22_65;
  assign out_21_64 = t_r21_c64_12 >> 4;

  assign t_r22_c1_0 = p_21_1 << 1;
  assign t_r22_c1_1 = p_22_0 << 1;
  assign t_r22_c1_2 = p_22_1 << 2;
  assign t_r22_c1_3 = p_22_2 << 1;
  assign t_r22_c1_4 = p_23_1 << 1;
  assign t_r22_c1_5 = t_r22_c1_0 + p_21_0;
  assign t_r22_c1_6 = t_r22_c1_1 + p_21_2;
  assign t_r22_c1_7 = t_r22_c1_2 + t_r22_c1_3;
  assign t_r22_c1_8 = t_r22_c1_4 + p_23_0;
  assign t_r22_c1_9 = t_r22_c1_5 + t_r22_c1_6;
  assign t_r22_c1_10 = t_r22_c1_7 + t_r22_c1_8;
  assign t_r22_c1_11 = t_r22_c1_9 + t_r22_c1_10;
  assign t_r22_c1_12 = t_r22_c1_11 + p_23_2;
  assign out_22_1 = t_r22_c1_12 >> 4;

  assign t_r22_c2_0 = p_21_2 << 1;
  assign t_r22_c2_1 = p_22_1 << 1;
  assign t_r22_c2_2 = p_22_2 << 2;
  assign t_r22_c2_3 = p_22_3 << 1;
  assign t_r22_c2_4 = p_23_2 << 1;
  assign t_r22_c2_5 = t_r22_c2_0 + p_21_1;
  assign t_r22_c2_6 = t_r22_c2_1 + p_21_3;
  assign t_r22_c2_7 = t_r22_c2_2 + t_r22_c2_3;
  assign t_r22_c2_8 = t_r22_c2_4 + p_23_1;
  assign t_r22_c2_9 = t_r22_c2_5 + t_r22_c2_6;
  assign t_r22_c2_10 = t_r22_c2_7 + t_r22_c2_8;
  assign t_r22_c2_11 = t_r22_c2_9 + t_r22_c2_10;
  assign t_r22_c2_12 = t_r22_c2_11 + p_23_3;
  assign out_22_2 = t_r22_c2_12 >> 4;

  assign t_r22_c3_0 = p_21_3 << 1;
  assign t_r22_c3_1 = p_22_2 << 1;
  assign t_r22_c3_2 = p_22_3 << 2;
  assign t_r22_c3_3 = p_22_4 << 1;
  assign t_r22_c3_4 = p_23_3 << 1;
  assign t_r22_c3_5 = t_r22_c3_0 + p_21_2;
  assign t_r22_c3_6 = t_r22_c3_1 + p_21_4;
  assign t_r22_c3_7 = t_r22_c3_2 + t_r22_c3_3;
  assign t_r22_c3_8 = t_r22_c3_4 + p_23_2;
  assign t_r22_c3_9 = t_r22_c3_5 + t_r22_c3_6;
  assign t_r22_c3_10 = t_r22_c3_7 + t_r22_c3_8;
  assign t_r22_c3_11 = t_r22_c3_9 + t_r22_c3_10;
  assign t_r22_c3_12 = t_r22_c3_11 + p_23_4;
  assign out_22_3 = t_r22_c3_12 >> 4;

  assign t_r22_c4_0 = p_21_4 << 1;
  assign t_r22_c4_1 = p_22_3 << 1;
  assign t_r22_c4_2 = p_22_4 << 2;
  assign t_r22_c4_3 = p_22_5 << 1;
  assign t_r22_c4_4 = p_23_4 << 1;
  assign t_r22_c4_5 = t_r22_c4_0 + p_21_3;
  assign t_r22_c4_6 = t_r22_c4_1 + p_21_5;
  assign t_r22_c4_7 = t_r22_c4_2 + t_r22_c4_3;
  assign t_r22_c4_8 = t_r22_c4_4 + p_23_3;
  assign t_r22_c4_9 = t_r22_c4_5 + t_r22_c4_6;
  assign t_r22_c4_10 = t_r22_c4_7 + t_r22_c4_8;
  assign t_r22_c4_11 = t_r22_c4_9 + t_r22_c4_10;
  assign t_r22_c4_12 = t_r22_c4_11 + p_23_5;
  assign out_22_4 = t_r22_c4_12 >> 4;

  assign t_r22_c5_0 = p_21_5 << 1;
  assign t_r22_c5_1 = p_22_4 << 1;
  assign t_r22_c5_2 = p_22_5 << 2;
  assign t_r22_c5_3 = p_22_6 << 1;
  assign t_r22_c5_4 = p_23_5 << 1;
  assign t_r22_c5_5 = t_r22_c5_0 + p_21_4;
  assign t_r22_c5_6 = t_r22_c5_1 + p_21_6;
  assign t_r22_c5_7 = t_r22_c5_2 + t_r22_c5_3;
  assign t_r22_c5_8 = t_r22_c5_4 + p_23_4;
  assign t_r22_c5_9 = t_r22_c5_5 + t_r22_c5_6;
  assign t_r22_c5_10 = t_r22_c5_7 + t_r22_c5_8;
  assign t_r22_c5_11 = t_r22_c5_9 + t_r22_c5_10;
  assign t_r22_c5_12 = t_r22_c5_11 + p_23_6;
  assign out_22_5 = t_r22_c5_12 >> 4;

  assign t_r22_c6_0 = p_21_6 << 1;
  assign t_r22_c6_1 = p_22_5 << 1;
  assign t_r22_c6_2 = p_22_6 << 2;
  assign t_r22_c6_3 = p_22_7 << 1;
  assign t_r22_c6_4 = p_23_6 << 1;
  assign t_r22_c6_5 = t_r22_c6_0 + p_21_5;
  assign t_r22_c6_6 = t_r22_c6_1 + p_21_7;
  assign t_r22_c6_7 = t_r22_c6_2 + t_r22_c6_3;
  assign t_r22_c6_8 = t_r22_c6_4 + p_23_5;
  assign t_r22_c6_9 = t_r22_c6_5 + t_r22_c6_6;
  assign t_r22_c6_10 = t_r22_c6_7 + t_r22_c6_8;
  assign t_r22_c6_11 = t_r22_c6_9 + t_r22_c6_10;
  assign t_r22_c6_12 = t_r22_c6_11 + p_23_7;
  assign out_22_6 = t_r22_c6_12 >> 4;

  assign t_r22_c7_0 = p_21_7 << 1;
  assign t_r22_c7_1 = p_22_6 << 1;
  assign t_r22_c7_2 = p_22_7 << 2;
  assign t_r22_c7_3 = p_22_8 << 1;
  assign t_r22_c7_4 = p_23_7 << 1;
  assign t_r22_c7_5 = t_r22_c7_0 + p_21_6;
  assign t_r22_c7_6 = t_r22_c7_1 + p_21_8;
  assign t_r22_c7_7 = t_r22_c7_2 + t_r22_c7_3;
  assign t_r22_c7_8 = t_r22_c7_4 + p_23_6;
  assign t_r22_c7_9 = t_r22_c7_5 + t_r22_c7_6;
  assign t_r22_c7_10 = t_r22_c7_7 + t_r22_c7_8;
  assign t_r22_c7_11 = t_r22_c7_9 + t_r22_c7_10;
  assign t_r22_c7_12 = t_r22_c7_11 + p_23_8;
  assign out_22_7 = t_r22_c7_12 >> 4;

  assign t_r22_c8_0 = p_21_8 << 1;
  assign t_r22_c8_1 = p_22_7 << 1;
  assign t_r22_c8_2 = p_22_8 << 2;
  assign t_r22_c8_3 = p_22_9 << 1;
  assign t_r22_c8_4 = p_23_8 << 1;
  assign t_r22_c8_5 = t_r22_c8_0 + p_21_7;
  assign t_r22_c8_6 = t_r22_c8_1 + p_21_9;
  assign t_r22_c8_7 = t_r22_c8_2 + t_r22_c8_3;
  assign t_r22_c8_8 = t_r22_c8_4 + p_23_7;
  assign t_r22_c8_9 = t_r22_c8_5 + t_r22_c8_6;
  assign t_r22_c8_10 = t_r22_c8_7 + t_r22_c8_8;
  assign t_r22_c8_11 = t_r22_c8_9 + t_r22_c8_10;
  assign t_r22_c8_12 = t_r22_c8_11 + p_23_9;
  assign out_22_8 = t_r22_c8_12 >> 4;

  assign t_r22_c9_0 = p_21_9 << 1;
  assign t_r22_c9_1 = p_22_8 << 1;
  assign t_r22_c9_2 = p_22_9 << 2;
  assign t_r22_c9_3 = p_22_10 << 1;
  assign t_r22_c9_4 = p_23_9 << 1;
  assign t_r22_c9_5 = t_r22_c9_0 + p_21_8;
  assign t_r22_c9_6 = t_r22_c9_1 + p_21_10;
  assign t_r22_c9_7 = t_r22_c9_2 + t_r22_c9_3;
  assign t_r22_c9_8 = t_r22_c9_4 + p_23_8;
  assign t_r22_c9_9 = t_r22_c9_5 + t_r22_c9_6;
  assign t_r22_c9_10 = t_r22_c9_7 + t_r22_c9_8;
  assign t_r22_c9_11 = t_r22_c9_9 + t_r22_c9_10;
  assign t_r22_c9_12 = t_r22_c9_11 + p_23_10;
  assign out_22_9 = t_r22_c9_12 >> 4;

  assign t_r22_c10_0 = p_21_10 << 1;
  assign t_r22_c10_1 = p_22_9 << 1;
  assign t_r22_c10_2 = p_22_10 << 2;
  assign t_r22_c10_3 = p_22_11 << 1;
  assign t_r22_c10_4 = p_23_10 << 1;
  assign t_r22_c10_5 = t_r22_c10_0 + p_21_9;
  assign t_r22_c10_6 = t_r22_c10_1 + p_21_11;
  assign t_r22_c10_7 = t_r22_c10_2 + t_r22_c10_3;
  assign t_r22_c10_8 = t_r22_c10_4 + p_23_9;
  assign t_r22_c10_9 = t_r22_c10_5 + t_r22_c10_6;
  assign t_r22_c10_10 = t_r22_c10_7 + t_r22_c10_8;
  assign t_r22_c10_11 = t_r22_c10_9 + t_r22_c10_10;
  assign t_r22_c10_12 = t_r22_c10_11 + p_23_11;
  assign out_22_10 = t_r22_c10_12 >> 4;

  assign t_r22_c11_0 = p_21_11 << 1;
  assign t_r22_c11_1 = p_22_10 << 1;
  assign t_r22_c11_2 = p_22_11 << 2;
  assign t_r22_c11_3 = p_22_12 << 1;
  assign t_r22_c11_4 = p_23_11 << 1;
  assign t_r22_c11_5 = t_r22_c11_0 + p_21_10;
  assign t_r22_c11_6 = t_r22_c11_1 + p_21_12;
  assign t_r22_c11_7 = t_r22_c11_2 + t_r22_c11_3;
  assign t_r22_c11_8 = t_r22_c11_4 + p_23_10;
  assign t_r22_c11_9 = t_r22_c11_5 + t_r22_c11_6;
  assign t_r22_c11_10 = t_r22_c11_7 + t_r22_c11_8;
  assign t_r22_c11_11 = t_r22_c11_9 + t_r22_c11_10;
  assign t_r22_c11_12 = t_r22_c11_11 + p_23_12;
  assign out_22_11 = t_r22_c11_12 >> 4;

  assign t_r22_c12_0 = p_21_12 << 1;
  assign t_r22_c12_1 = p_22_11 << 1;
  assign t_r22_c12_2 = p_22_12 << 2;
  assign t_r22_c12_3 = p_22_13 << 1;
  assign t_r22_c12_4 = p_23_12 << 1;
  assign t_r22_c12_5 = t_r22_c12_0 + p_21_11;
  assign t_r22_c12_6 = t_r22_c12_1 + p_21_13;
  assign t_r22_c12_7 = t_r22_c12_2 + t_r22_c12_3;
  assign t_r22_c12_8 = t_r22_c12_4 + p_23_11;
  assign t_r22_c12_9 = t_r22_c12_5 + t_r22_c12_6;
  assign t_r22_c12_10 = t_r22_c12_7 + t_r22_c12_8;
  assign t_r22_c12_11 = t_r22_c12_9 + t_r22_c12_10;
  assign t_r22_c12_12 = t_r22_c12_11 + p_23_13;
  assign out_22_12 = t_r22_c12_12 >> 4;

  assign t_r22_c13_0 = p_21_13 << 1;
  assign t_r22_c13_1 = p_22_12 << 1;
  assign t_r22_c13_2 = p_22_13 << 2;
  assign t_r22_c13_3 = p_22_14 << 1;
  assign t_r22_c13_4 = p_23_13 << 1;
  assign t_r22_c13_5 = t_r22_c13_0 + p_21_12;
  assign t_r22_c13_6 = t_r22_c13_1 + p_21_14;
  assign t_r22_c13_7 = t_r22_c13_2 + t_r22_c13_3;
  assign t_r22_c13_8 = t_r22_c13_4 + p_23_12;
  assign t_r22_c13_9 = t_r22_c13_5 + t_r22_c13_6;
  assign t_r22_c13_10 = t_r22_c13_7 + t_r22_c13_8;
  assign t_r22_c13_11 = t_r22_c13_9 + t_r22_c13_10;
  assign t_r22_c13_12 = t_r22_c13_11 + p_23_14;
  assign out_22_13 = t_r22_c13_12 >> 4;

  assign t_r22_c14_0 = p_21_14 << 1;
  assign t_r22_c14_1 = p_22_13 << 1;
  assign t_r22_c14_2 = p_22_14 << 2;
  assign t_r22_c14_3 = p_22_15 << 1;
  assign t_r22_c14_4 = p_23_14 << 1;
  assign t_r22_c14_5 = t_r22_c14_0 + p_21_13;
  assign t_r22_c14_6 = t_r22_c14_1 + p_21_15;
  assign t_r22_c14_7 = t_r22_c14_2 + t_r22_c14_3;
  assign t_r22_c14_8 = t_r22_c14_4 + p_23_13;
  assign t_r22_c14_9 = t_r22_c14_5 + t_r22_c14_6;
  assign t_r22_c14_10 = t_r22_c14_7 + t_r22_c14_8;
  assign t_r22_c14_11 = t_r22_c14_9 + t_r22_c14_10;
  assign t_r22_c14_12 = t_r22_c14_11 + p_23_15;
  assign out_22_14 = t_r22_c14_12 >> 4;

  assign t_r22_c15_0 = p_21_15 << 1;
  assign t_r22_c15_1 = p_22_14 << 1;
  assign t_r22_c15_2 = p_22_15 << 2;
  assign t_r22_c15_3 = p_22_16 << 1;
  assign t_r22_c15_4 = p_23_15 << 1;
  assign t_r22_c15_5 = t_r22_c15_0 + p_21_14;
  assign t_r22_c15_6 = t_r22_c15_1 + p_21_16;
  assign t_r22_c15_7 = t_r22_c15_2 + t_r22_c15_3;
  assign t_r22_c15_8 = t_r22_c15_4 + p_23_14;
  assign t_r22_c15_9 = t_r22_c15_5 + t_r22_c15_6;
  assign t_r22_c15_10 = t_r22_c15_7 + t_r22_c15_8;
  assign t_r22_c15_11 = t_r22_c15_9 + t_r22_c15_10;
  assign t_r22_c15_12 = t_r22_c15_11 + p_23_16;
  assign out_22_15 = t_r22_c15_12 >> 4;

  assign t_r22_c16_0 = p_21_16 << 1;
  assign t_r22_c16_1 = p_22_15 << 1;
  assign t_r22_c16_2 = p_22_16 << 2;
  assign t_r22_c16_3 = p_22_17 << 1;
  assign t_r22_c16_4 = p_23_16 << 1;
  assign t_r22_c16_5 = t_r22_c16_0 + p_21_15;
  assign t_r22_c16_6 = t_r22_c16_1 + p_21_17;
  assign t_r22_c16_7 = t_r22_c16_2 + t_r22_c16_3;
  assign t_r22_c16_8 = t_r22_c16_4 + p_23_15;
  assign t_r22_c16_9 = t_r22_c16_5 + t_r22_c16_6;
  assign t_r22_c16_10 = t_r22_c16_7 + t_r22_c16_8;
  assign t_r22_c16_11 = t_r22_c16_9 + t_r22_c16_10;
  assign t_r22_c16_12 = t_r22_c16_11 + p_23_17;
  assign out_22_16 = t_r22_c16_12 >> 4;

  assign t_r22_c17_0 = p_21_17 << 1;
  assign t_r22_c17_1 = p_22_16 << 1;
  assign t_r22_c17_2 = p_22_17 << 2;
  assign t_r22_c17_3 = p_22_18 << 1;
  assign t_r22_c17_4 = p_23_17 << 1;
  assign t_r22_c17_5 = t_r22_c17_0 + p_21_16;
  assign t_r22_c17_6 = t_r22_c17_1 + p_21_18;
  assign t_r22_c17_7 = t_r22_c17_2 + t_r22_c17_3;
  assign t_r22_c17_8 = t_r22_c17_4 + p_23_16;
  assign t_r22_c17_9 = t_r22_c17_5 + t_r22_c17_6;
  assign t_r22_c17_10 = t_r22_c17_7 + t_r22_c17_8;
  assign t_r22_c17_11 = t_r22_c17_9 + t_r22_c17_10;
  assign t_r22_c17_12 = t_r22_c17_11 + p_23_18;
  assign out_22_17 = t_r22_c17_12 >> 4;

  assign t_r22_c18_0 = p_21_18 << 1;
  assign t_r22_c18_1 = p_22_17 << 1;
  assign t_r22_c18_2 = p_22_18 << 2;
  assign t_r22_c18_3 = p_22_19 << 1;
  assign t_r22_c18_4 = p_23_18 << 1;
  assign t_r22_c18_5 = t_r22_c18_0 + p_21_17;
  assign t_r22_c18_6 = t_r22_c18_1 + p_21_19;
  assign t_r22_c18_7 = t_r22_c18_2 + t_r22_c18_3;
  assign t_r22_c18_8 = t_r22_c18_4 + p_23_17;
  assign t_r22_c18_9 = t_r22_c18_5 + t_r22_c18_6;
  assign t_r22_c18_10 = t_r22_c18_7 + t_r22_c18_8;
  assign t_r22_c18_11 = t_r22_c18_9 + t_r22_c18_10;
  assign t_r22_c18_12 = t_r22_c18_11 + p_23_19;
  assign out_22_18 = t_r22_c18_12 >> 4;

  assign t_r22_c19_0 = p_21_19 << 1;
  assign t_r22_c19_1 = p_22_18 << 1;
  assign t_r22_c19_2 = p_22_19 << 2;
  assign t_r22_c19_3 = p_22_20 << 1;
  assign t_r22_c19_4 = p_23_19 << 1;
  assign t_r22_c19_5 = t_r22_c19_0 + p_21_18;
  assign t_r22_c19_6 = t_r22_c19_1 + p_21_20;
  assign t_r22_c19_7 = t_r22_c19_2 + t_r22_c19_3;
  assign t_r22_c19_8 = t_r22_c19_4 + p_23_18;
  assign t_r22_c19_9 = t_r22_c19_5 + t_r22_c19_6;
  assign t_r22_c19_10 = t_r22_c19_7 + t_r22_c19_8;
  assign t_r22_c19_11 = t_r22_c19_9 + t_r22_c19_10;
  assign t_r22_c19_12 = t_r22_c19_11 + p_23_20;
  assign out_22_19 = t_r22_c19_12 >> 4;

  assign t_r22_c20_0 = p_21_20 << 1;
  assign t_r22_c20_1 = p_22_19 << 1;
  assign t_r22_c20_2 = p_22_20 << 2;
  assign t_r22_c20_3 = p_22_21 << 1;
  assign t_r22_c20_4 = p_23_20 << 1;
  assign t_r22_c20_5 = t_r22_c20_0 + p_21_19;
  assign t_r22_c20_6 = t_r22_c20_1 + p_21_21;
  assign t_r22_c20_7 = t_r22_c20_2 + t_r22_c20_3;
  assign t_r22_c20_8 = t_r22_c20_4 + p_23_19;
  assign t_r22_c20_9 = t_r22_c20_5 + t_r22_c20_6;
  assign t_r22_c20_10 = t_r22_c20_7 + t_r22_c20_8;
  assign t_r22_c20_11 = t_r22_c20_9 + t_r22_c20_10;
  assign t_r22_c20_12 = t_r22_c20_11 + p_23_21;
  assign out_22_20 = t_r22_c20_12 >> 4;

  assign t_r22_c21_0 = p_21_21 << 1;
  assign t_r22_c21_1 = p_22_20 << 1;
  assign t_r22_c21_2 = p_22_21 << 2;
  assign t_r22_c21_3 = p_22_22 << 1;
  assign t_r22_c21_4 = p_23_21 << 1;
  assign t_r22_c21_5 = t_r22_c21_0 + p_21_20;
  assign t_r22_c21_6 = t_r22_c21_1 + p_21_22;
  assign t_r22_c21_7 = t_r22_c21_2 + t_r22_c21_3;
  assign t_r22_c21_8 = t_r22_c21_4 + p_23_20;
  assign t_r22_c21_9 = t_r22_c21_5 + t_r22_c21_6;
  assign t_r22_c21_10 = t_r22_c21_7 + t_r22_c21_8;
  assign t_r22_c21_11 = t_r22_c21_9 + t_r22_c21_10;
  assign t_r22_c21_12 = t_r22_c21_11 + p_23_22;
  assign out_22_21 = t_r22_c21_12 >> 4;

  assign t_r22_c22_0 = p_21_22 << 1;
  assign t_r22_c22_1 = p_22_21 << 1;
  assign t_r22_c22_2 = p_22_22 << 2;
  assign t_r22_c22_3 = p_22_23 << 1;
  assign t_r22_c22_4 = p_23_22 << 1;
  assign t_r22_c22_5 = t_r22_c22_0 + p_21_21;
  assign t_r22_c22_6 = t_r22_c22_1 + p_21_23;
  assign t_r22_c22_7 = t_r22_c22_2 + t_r22_c22_3;
  assign t_r22_c22_8 = t_r22_c22_4 + p_23_21;
  assign t_r22_c22_9 = t_r22_c22_5 + t_r22_c22_6;
  assign t_r22_c22_10 = t_r22_c22_7 + t_r22_c22_8;
  assign t_r22_c22_11 = t_r22_c22_9 + t_r22_c22_10;
  assign t_r22_c22_12 = t_r22_c22_11 + p_23_23;
  assign out_22_22 = t_r22_c22_12 >> 4;

  assign t_r22_c23_0 = p_21_23 << 1;
  assign t_r22_c23_1 = p_22_22 << 1;
  assign t_r22_c23_2 = p_22_23 << 2;
  assign t_r22_c23_3 = p_22_24 << 1;
  assign t_r22_c23_4 = p_23_23 << 1;
  assign t_r22_c23_5 = t_r22_c23_0 + p_21_22;
  assign t_r22_c23_6 = t_r22_c23_1 + p_21_24;
  assign t_r22_c23_7 = t_r22_c23_2 + t_r22_c23_3;
  assign t_r22_c23_8 = t_r22_c23_4 + p_23_22;
  assign t_r22_c23_9 = t_r22_c23_5 + t_r22_c23_6;
  assign t_r22_c23_10 = t_r22_c23_7 + t_r22_c23_8;
  assign t_r22_c23_11 = t_r22_c23_9 + t_r22_c23_10;
  assign t_r22_c23_12 = t_r22_c23_11 + p_23_24;
  assign out_22_23 = t_r22_c23_12 >> 4;

  assign t_r22_c24_0 = p_21_24 << 1;
  assign t_r22_c24_1 = p_22_23 << 1;
  assign t_r22_c24_2 = p_22_24 << 2;
  assign t_r22_c24_3 = p_22_25 << 1;
  assign t_r22_c24_4 = p_23_24 << 1;
  assign t_r22_c24_5 = t_r22_c24_0 + p_21_23;
  assign t_r22_c24_6 = t_r22_c24_1 + p_21_25;
  assign t_r22_c24_7 = t_r22_c24_2 + t_r22_c24_3;
  assign t_r22_c24_8 = t_r22_c24_4 + p_23_23;
  assign t_r22_c24_9 = t_r22_c24_5 + t_r22_c24_6;
  assign t_r22_c24_10 = t_r22_c24_7 + t_r22_c24_8;
  assign t_r22_c24_11 = t_r22_c24_9 + t_r22_c24_10;
  assign t_r22_c24_12 = t_r22_c24_11 + p_23_25;
  assign out_22_24 = t_r22_c24_12 >> 4;

  assign t_r22_c25_0 = p_21_25 << 1;
  assign t_r22_c25_1 = p_22_24 << 1;
  assign t_r22_c25_2 = p_22_25 << 2;
  assign t_r22_c25_3 = p_22_26 << 1;
  assign t_r22_c25_4 = p_23_25 << 1;
  assign t_r22_c25_5 = t_r22_c25_0 + p_21_24;
  assign t_r22_c25_6 = t_r22_c25_1 + p_21_26;
  assign t_r22_c25_7 = t_r22_c25_2 + t_r22_c25_3;
  assign t_r22_c25_8 = t_r22_c25_4 + p_23_24;
  assign t_r22_c25_9 = t_r22_c25_5 + t_r22_c25_6;
  assign t_r22_c25_10 = t_r22_c25_7 + t_r22_c25_8;
  assign t_r22_c25_11 = t_r22_c25_9 + t_r22_c25_10;
  assign t_r22_c25_12 = t_r22_c25_11 + p_23_26;
  assign out_22_25 = t_r22_c25_12 >> 4;

  assign t_r22_c26_0 = p_21_26 << 1;
  assign t_r22_c26_1 = p_22_25 << 1;
  assign t_r22_c26_2 = p_22_26 << 2;
  assign t_r22_c26_3 = p_22_27 << 1;
  assign t_r22_c26_4 = p_23_26 << 1;
  assign t_r22_c26_5 = t_r22_c26_0 + p_21_25;
  assign t_r22_c26_6 = t_r22_c26_1 + p_21_27;
  assign t_r22_c26_7 = t_r22_c26_2 + t_r22_c26_3;
  assign t_r22_c26_8 = t_r22_c26_4 + p_23_25;
  assign t_r22_c26_9 = t_r22_c26_5 + t_r22_c26_6;
  assign t_r22_c26_10 = t_r22_c26_7 + t_r22_c26_8;
  assign t_r22_c26_11 = t_r22_c26_9 + t_r22_c26_10;
  assign t_r22_c26_12 = t_r22_c26_11 + p_23_27;
  assign out_22_26 = t_r22_c26_12 >> 4;

  assign t_r22_c27_0 = p_21_27 << 1;
  assign t_r22_c27_1 = p_22_26 << 1;
  assign t_r22_c27_2 = p_22_27 << 2;
  assign t_r22_c27_3 = p_22_28 << 1;
  assign t_r22_c27_4 = p_23_27 << 1;
  assign t_r22_c27_5 = t_r22_c27_0 + p_21_26;
  assign t_r22_c27_6 = t_r22_c27_1 + p_21_28;
  assign t_r22_c27_7 = t_r22_c27_2 + t_r22_c27_3;
  assign t_r22_c27_8 = t_r22_c27_4 + p_23_26;
  assign t_r22_c27_9 = t_r22_c27_5 + t_r22_c27_6;
  assign t_r22_c27_10 = t_r22_c27_7 + t_r22_c27_8;
  assign t_r22_c27_11 = t_r22_c27_9 + t_r22_c27_10;
  assign t_r22_c27_12 = t_r22_c27_11 + p_23_28;
  assign out_22_27 = t_r22_c27_12 >> 4;

  assign t_r22_c28_0 = p_21_28 << 1;
  assign t_r22_c28_1 = p_22_27 << 1;
  assign t_r22_c28_2 = p_22_28 << 2;
  assign t_r22_c28_3 = p_22_29 << 1;
  assign t_r22_c28_4 = p_23_28 << 1;
  assign t_r22_c28_5 = t_r22_c28_0 + p_21_27;
  assign t_r22_c28_6 = t_r22_c28_1 + p_21_29;
  assign t_r22_c28_7 = t_r22_c28_2 + t_r22_c28_3;
  assign t_r22_c28_8 = t_r22_c28_4 + p_23_27;
  assign t_r22_c28_9 = t_r22_c28_5 + t_r22_c28_6;
  assign t_r22_c28_10 = t_r22_c28_7 + t_r22_c28_8;
  assign t_r22_c28_11 = t_r22_c28_9 + t_r22_c28_10;
  assign t_r22_c28_12 = t_r22_c28_11 + p_23_29;
  assign out_22_28 = t_r22_c28_12 >> 4;

  assign t_r22_c29_0 = p_21_29 << 1;
  assign t_r22_c29_1 = p_22_28 << 1;
  assign t_r22_c29_2 = p_22_29 << 2;
  assign t_r22_c29_3 = p_22_30 << 1;
  assign t_r22_c29_4 = p_23_29 << 1;
  assign t_r22_c29_5 = t_r22_c29_0 + p_21_28;
  assign t_r22_c29_6 = t_r22_c29_1 + p_21_30;
  assign t_r22_c29_7 = t_r22_c29_2 + t_r22_c29_3;
  assign t_r22_c29_8 = t_r22_c29_4 + p_23_28;
  assign t_r22_c29_9 = t_r22_c29_5 + t_r22_c29_6;
  assign t_r22_c29_10 = t_r22_c29_7 + t_r22_c29_8;
  assign t_r22_c29_11 = t_r22_c29_9 + t_r22_c29_10;
  assign t_r22_c29_12 = t_r22_c29_11 + p_23_30;
  assign out_22_29 = t_r22_c29_12 >> 4;

  assign t_r22_c30_0 = p_21_30 << 1;
  assign t_r22_c30_1 = p_22_29 << 1;
  assign t_r22_c30_2 = p_22_30 << 2;
  assign t_r22_c30_3 = p_22_31 << 1;
  assign t_r22_c30_4 = p_23_30 << 1;
  assign t_r22_c30_5 = t_r22_c30_0 + p_21_29;
  assign t_r22_c30_6 = t_r22_c30_1 + p_21_31;
  assign t_r22_c30_7 = t_r22_c30_2 + t_r22_c30_3;
  assign t_r22_c30_8 = t_r22_c30_4 + p_23_29;
  assign t_r22_c30_9 = t_r22_c30_5 + t_r22_c30_6;
  assign t_r22_c30_10 = t_r22_c30_7 + t_r22_c30_8;
  assign t_r22_c30_11 = t_r22_c30_9 + t_r22_c30_10;
  assign t_r22_c30_12 = t_r22_c30_11 + p_23_31;
  assign out_22_30 = t_r22_c30_12 >> 4;

  assign t_r22_c31_0 = p_21_31 << 1;
  assign t_r22_c31_1 = p_22_30 << 1;
  assign t_r22_c31_2 = p_22_31 << 2;
  assign t_r22_c31_3 = p_22_32 << 1;
  assign t_r22_c31_4 = p_23_31 << 1;
  assign t_r22_c31_5 = t_r22_c31_0 + p_21_30;
  assign t_r22_c31_6 = t_r22_c31_1 + p_21_32;
  assign t_r22_c31_7 = t_r22_c31_2 + t_r22_c31_3;
  assign t_r22_c31_8 = t_r22_c31_4 + p_23_30;
  assign t_r22_c31_9 = t_r22_c31_5 + t_r22_c31_6;
  assign t_r22_c31_10 = t_r22_c31_7 + t_r22_c31_8;
  assign t_r22_c31_11 = t_r22_c31_9 + t_r22_c31_10;
  assign t_r22_c31_12 = t_r22_c31_11 + p_23_32;
  assign out_22_31 = t_r22_c31_12 >> 4;

  assign t_r22_c32_0 = p_21_32 << 1;
  assign t_r22_c32_1 = p_22_31 << 1;
  assign t_r22_c32_2 = p_22_32 << 2;
  assign t_r22_c32_3 = p_22_33 << 1;
  assign t_r22_c32_4 = p_23_32 << 1;
  assign t_r22_c32_5 = t_r22_c32_0 + p_21_31;
  assign t_r22_c32_6 = t_r22_c32_1 + p_21_33;
  assign t_r22_c32_7 = t_r22_c32_2 + t_r22_c32_3;
  assign t_r22_c32_8 = t_r22_c32_4 + p_23_31;
  assign t_r22_c32_9 = t_r22_c32_5 + t_r22_c32_6;
  assign t_r22_c32_10 = t_r22_c32_7 + t_r22_c32_8;
  assign t_r22_c32_11 = t_r22_c32_9 + t_r22_c32_10;
  assign t_r22_c32_12 = t_r22_c32_11 + p_23_33;
  assign out_22_32 = t_r22_c32_12 >> 4;

  assign t_r22_c33_0 = p_21_33 << 1;
  assign t_r22_c33_1 = p_22_32 << 1;
  assign t_r22_c33_2 = p_22_33 << 2;
  assign t_r22_c33_3 = p_22_34 << 1;
  assign t_r22_c33_4 = p_23_33 << 1;
  assign t_r22_c33_5 = t_r22_c33_0 + p_21_32;
  assign t_r22_c33_6 = t_r22_c33_1 + p_21_34;
  assign t_r22_c33_7 = t_r22_c33_2 + t_r22_c33_3;
  assign t_r22_c33_8 = t_r22_c33_4 + p_23_32;
  assign t_r22_c33_9 = t_r22_c33_5 + t_r22_c33_6;
  assign t_r22_c33_10 = t_r22_c33_7 + t_r22_c33_8;
  assign t_r22_c33_11 = t_r22_c33_9 + t_r22_c33_10;
  assign t_r22_c33_12 = t_r22_c33_11 + p_23_34;
  assign out_22_33 = t_r22_c33_12 >> 4;

  assign t_r22_c34_0 = p_21_34 << 1;
  assign t_r22_c34_1 = p_22_33 << 1;
  assign t_r22_c34_2 = p_22_34 << 2;
  assign t_r22_c34_3 = p_22_35 << 1;
  assign t_r22_c34_4 = p_23_34 << 1;
  assign t_r22_c34_5 = t_r22_c34_0 + p_21_33;
  assign t_r22_c34_6 = t_r22_c34_1 + p_21_35;
  assign t_r22_c34_7 = t_r22_c34_2 + t_r22_c34_3;
  assign t_r22_c34_8 = t_r22_c34_4 + p_23_33;
  assign t_r22_c34_9 = t_r22_c34_5 + t_r22_c34_6;
  assign t_r22_c34_10 = t_r22_c34_7 + t_r22_c34_8;
  assign t_r22_c34_11 = t_r22_c34_9 + t_r22_c34_10;
  assign t_r22_c34_12 = t_r22_c34_11 + p_23_35;
  assign out_22_34 = t_r22_c34_12 >> 4;

  assign t_r22_c35_0 = p_21_35 << 1;
  assign t_r22_c35_1 = p_22_34 << 1;
  assign t_r22_c35_2 = p_22_35 << 2;
  assign t_r22_c35_3 = p_22_36 << 1;
  assign t_r22_c35_4 = p_23_35 << 1;
  assign t_r22_c35_5 = t_r22_c35_0 + p_21_34;
  assign t_r22_c35_6 = t_r22_c35_1 + p_21_36;
  assign t_r22_c35_7 = t_r22_c35_2 + t_r22_c35_3;
  assign t_r22_c35_8 = t_r22_c35_4 + p_23_34;
  assign t_r22_c35_9 = t_r22_c35_5 + t_r22_c35_6;
  assign t_r22_c35_10 = t_r22_c35_7 + t_r22_c35_8;
  assign t_r22_c35_11 = t_r22_c35_9 + t_r22_c35_10;
  assign t_r22_c35_12 = t_r22_c35_11 + p_23_36;
  assign out_22_35 = t_r22_c35_12 >> 4;

  assign t_r22_c36_0 = p_21_36 << 1;
  assign t_r22_c36_1 = p_22_35 << 1;
  assign t_r22_c36_2 = p_22_36 << 2;
  assign t_r22_c36_3 = p_22_37 << 1;
  assign t_r22_c36_4 = p_23_36 << 1;
  assign t_r22_c36_5 = t_r22_c36_0 + p_21_35;
  assign t_r22_c36_6 = t_r22_c36_1 + p_21_37;
  assign t_r22_c36_7 = t_r22_c36_2 + t_r22_c36_3;
  assign t_r22_c36_8 = t_r22_c36_4 + p_23_35;
  assign t_r22_c36_9 = t_r22_c36_5 + t_r22_c36_6;
  assign t_r22_c36_10 = t_r22_c36_7 + t_r22_c36_8;
  assign t_r22_c36_11 = t_r22_c36_9 + t_r22_c36_10;
  assign t_r22_c36_12 = t_r22_c36_11 + p_23_37;
  assign out_22_36 = t_r22_c36_12 >> 4;

  assign t_r22_c37_0 = p_21_37 << 1;
  assign t_r22_c37_1 = p_22_36 << 1;
  assign t_r22_c37_2 = p_22_37 << 2;
  assign t_r22_c37_3 = p_22_38 << 1;
  assign t_r22_c37_4 = p_23_37 << 1;
  assign t_r22_c37_5 = t_r22_c37_0 + p_21_36;
  assign t_r22_c37_6 = t_r22_c37_1 + p_21_38;
  assign t_r22_c37_7 = t_r22_c37_2 + t_r22_c37_3;
  assign t_r22_c37_8 = t_r22_c37_4 + p_23_36;
  assign t_r22_c37_9 = t_r22_c37_5 + t_r22_c37_6;
  assign t_r22_c37_10 = t_r22_c37_7 + t_r22_c37_8;
  assign t_r22_c37_11 = t_r22_c37_9 + t_r22_c37_10;
  assign t_r22_c37_12 = t_r22_c37_11 + p_23_38;
  assign out_22_37 = t_r22_c37_12 >> 4;

  assign t_r22_c38_0 = p_21_38 << 1;
  assign t_r22_c38_1 = p_22_37 << 1;
  assign t_r22_c38_2 = p_22_38 << 2;
  assign t_r22_c38_3 = p_22_39 << 1;
  assign t_r22_c38_4 = p_23_38 << 1;
  assign t_r22_c38_5 = t_r22_c38_0 + p_21_37;
  assign t_r22_c38_6 = t_r22_c38_1 + p_21_39;
  assign t_r22_c38_7 = t_r22_c38_2 + t_r22_c38_3;
  assign t_r22_c38_8 = t_r22_c38_4 + p_23_37;
  assign t_r22_c38_9 = t_r22_c38_5 + t_r22_c38_6;
  assign t_r22_c38_10 = t_r22_c38_7 + t_r22_c38_8;
  assign t_r22_c38_11 = t_r22_c38_9 + t_r22_c38_10;
  assign t_r22_c38_12 = t_r22_c38_11 + p_23_39;
  assign out_22_38 = t_r22_c38_12 >> 4;

  assign t_r22_c39_0 = p_21_39 << 1;
  assign t_r22_c39_1 = p_22_38 << 1;
  assign t_r22_c39_2 = p_22_39 << 2;
  assign t_r22_c39_3 = p_22_40 << 1;
  assign t_r22_c39_4 = p_23_39 << 1;
  assign t_r22_c39_5 = t_r22_c39_0 + p_21_38;
  assign t_r22_c39_6 = t_r22_c39_1 + p_21_40;
  assign t_r22_c39_7 = t_r22_c39_2 + t_r22_c39_3;
  assign t_r22_c39_8 = t_r22_c39_4 + p_23_38;
  assign t_r22_c39_9 = t_r22_c39_5 + t_r22_c39_6;
  assign t_r22_c39_10 = t_r22_c39_7 + t_r22_c39_8;
  assign t_r22_c39_11 = t_r22_c39_9 + t_r22_c39_10;
  assign t_r22_c39_12 = t_r22_c39_11 + p_23_40;
  assign out_22_39 = t_r22_c39_12 >> 4;

  assign t_r22_c40_0 = p_21_40 << 1;
  assign t_r22_c40_1 = p_22_39 << 1;
  assign t_r22_c40_2 = p_22_40 << 2;
  assign t_r22_c40_3 = p_22_41 << 1;
  assign t_r22_c40_4 = p_23_40 << 1;
  assign t_r22_c40_5 = t_r22_c40_0 + p_21_39;
  assign t_r22_c40_6 = t_r22_c40_1 + p_21_41;
  assign t_r22_c40_7 = t_r22_c40_2 + t_r22_c40_3;
  assign t_r22_c40_8 = t_r22_c40_4 + p_23_39;
  assign t_r22_c40_9 = t_r22_c40_5 + t_r22_c40_6;
  assign t_r22_c40_10 = t_r22_c40_7 + t_r22_c40_8;
  assign t_r22_c40_11 = t_r22_c40_9 + t_r22_c40_10;
  assign t_r22_c40_12 = t_r22_c40_11 + p_23_41;
  assign out_22_40 = t_r22_c40_12 >> 4;

  assign t_r22_c41_0 = p_21_41 << 1;
  assign t_r22_c41_1 = p_22_40 << 1;
  assign t_r22_c41_2 = p_22_41 << 2;
  assign t_r22_c41_3 = p_22_42 << 1;
  assign t_r22_c41_4 = p_23_41 << 1;
  assign t_r22_c41_5 = t_r22_c41_0 + p_21_40;
  assign t_r22_c41_6 = t_r22_c41_1 + p_21_42;
  assign t_r22_c41_7 = t_r22_c41_2 + t_r22_c41_3;
  assign t_r22_c41_8 = t_r22_c41_4 + p_23_40;
  assign t_r22_c41_9 = t_r22_c41_5 + t_r22_c41_6;
  assign t_r22_c41_10 = t_r22_c41_7 + t_r22_c41_8;
  assign t_r22_c41_11 = t_r22_c41_9 + t_r22_c41_10;
  assign t_r22_c41_12 = t_r22_c41_11 + p_23_42;
  assign out_22_41 = t_r22_c41_12 >> 4;

  assign t_r22_c42_0 = p_21_42 << 1;
  assign t_r22_c42_1 = p_22_41 << 1;
  assign t_r22_c42_2 = p_22_42 << 2;
  assign t_r22_c42_3 = p_22_43 << 1;
  assign t_r22_c42_4 = p_23_42 << 1;
  assign t_r22_c42_5 = t_r22_c42_0 + p_21_41;
  assign t_r22_c42_6 = t_r22_c42_1 + p_21_43;
  assign t_r22_c42_7 = t_r22_c42_2 + t_r22_c42_3;
  assign t_r22_c42_8 = t_r22_c42_4 + p_23_41;
  assign t_r22_c42_9 = t_r22_c42_5 + t_r22_c42_6;
  assign t_r22_c42_10 = t_r22_c42_7 + t_r22_c42_8;
  assign t_r22_c42_11 = t_r22_c42_9 + t_r22_c42_10;
  assign t_r22_c42_12 = t_r22_c42_11 + p_23_43;
  assign out_22_42 = t_r22_c42_12 >> 4;

  assign t_r22_c43_0 = p_21_43 << 1;
  assign t_r22_c43_1 = p_22_42 << 1;
  assign t_r22_c43_2 = p_22_43 << 2;
  assign t_r22_c43_3 = p_22_44 << 1;
  assign t_r22_c43_4 = p_23_43 << 1;
  assign t_r22_c43_5 = t_r22_c43_0 + p_21_42;
  assign t_r22_c43_6 = t_r22_c43_1 + p_21_44;
  assign t_r22_c43_7 = t_r22_c43_2 + t_r22_c43_3;
  assign t_r22_c43_8 = t_r22_c43_4 + p_23_42;
  assign t_r22_c43_9 = t_r22_c43_5 + t_r22_c43_6;
  assign t_r22_c43_10 = t_r22_c43_7 + t_r22_c43_8;
  assign t_r22_c43_11 = t_r22_c43_9 + t_r22_c43_10;
  assign t_r22_c43_12 = t_r22_c43_11 + p_23_44;
  assign out_22_43 = t_r22_c43_12 >> 4;

  assign t_r22_c44_0 = p_21_44 << 1;
  assign t_r22_c44_1 = p_22_43 << 1;
  assign t_r22_c44_2 = p_22_44 << 2;
  assign t_r22_c44_3 = p_22_45 << 1;
  assign t_r22_c44_4 = p_23_44 << 1;
  assign t_r22_c44_5 = t_r22_c44_0 + p_21_43;
  assign t_r22_c44_6 = t_r22_c44_1 + p_21_45;
  assign t_r22_c44_7 = t_r22_c44_2 + t_r22_c44_3;
  assign t_r22_c44_8 = t_r22_c44_4 + p_23_43;
  assign t_r22_c44_9 = t_r22_c44_5 + t_r22_c44_6;
  assign t_r22_c44_10 = t_r22_c44_7 + t_r22_c44_8;
  assign t_r22_c44_11 = t_r22_c44_9 + t_r22_c44_10;
  assign t_r22_c44_12 = t_r22_c44_11 + p_23_45;
  assign out_22_44 = t_r22_c44_12 >> 4;

  assign t_r22_c45_0 = p_21_45 << 1;
  assign t_r22_c45_1 = p_22_44 << 1;
  assign t_r22_c45_2 = p_22_45 << 2;
  assign t_r22_c45_3 = p_22_46 << 1;
  assign t_r22_c45_4 = p_23_45 << 1;
  assign t_r22_c45_5 = t_r22_c45_0 + p_21_44;
  assign t_r22_c45_6 = t_r22_c45_1 + p_21_46;
  assign t_r22_c45_7 = t_r22_c45_2 + t_r22_c45_3;
  assign t_r22_c45_8 = t_r22_c45_4 + p_23_44;
  assign t_r22_c45_9 = t_r22_c45_5 + t_r22_c45_6;
  assign t_r22_c45_10 = t_r22_c45_7 + t_r22_c45_8;
  assign t_r22_c45_11 = t_r22_c45_9 + t_r22_c45_10;
  assign t_r22_c45_12 = t_r22_c45_11 + p_23_46;
  assign out_22_45 = t_r22_c45_12 >> 4;

  assign t_r22_c46_0 = p_21_46 << 1;
  assign t_r22_c46_1 = p_22_45 << 1;
  assign t_r22_c46_2 = p_22_46 << 2;
  assign t_r22_c46_3 = p_22_47 << 1;
  assign t_r22_c46_4 = p_23_46 << 1;
  assign t_r22_c46_5 = t_r22_c46_0 + p_21_45;
  assign t_r22_c46_6 = t_r22_c46_1 + p_21_47;
  assign t_r22_c46_7 = t_r22_c46_2 + t_r22_c46_3;
  assign t_r22_c46_8 = t_r22_c46_4 + p_23_45;
  assign t_r22_c46_9 = t_r22_c46_5 + t_r22_c46_6;
  assign t_r22_c46_10 = t_r22_c46_7 + t_r22_c46_8;
  assign t_r22_c46_11 = t_r22_c46_9 + t_r22_c46_10;
  assign t_r22_c46_12 = t_r22_c46_11 + p_23_47;
  assign out_22_46 = t_r22_c46_12 >> 4;

  assign t_r22_c47_0 = p_21_47 << 1;
  assign t_r22_c47_1 = p_22_46 << 1;
  assign t_r22_c47_2 = p_22_47 << 2;
  assign t_r22_c47_3 = p_22_48 << 1;
  assign t_r22_c47_4 = p_23_47 << 1;
  assign t_r22_c47_5 = t_r22_c47_0 + p_21_46;
  assign t_r22_c47_6 = t_r22_c47_1 + p_21_48;
  assign t_r22_c47_7 = t_r22_c47_2 + t_r22_c47_3;
  assign t_r22_c47_8 = t_r22_c47_4 + p_23_46;
  assign t_r22_c47_9 = t_r22_c47_5 + t_r22_c47_6;
  assign t_r22_c47_10 = t_r22_c47_7 + t_r22_c47_8;
  assign t_r22_c47_11 = t_r22_c47_9 + t_r22_c47_10;
  assign t_r22_c47_12 = t_r22_c47_11 + p_23_48;
  assign out_22_47 = t_r22_c47_12 >> 4;

  assign t_r22_c48_0 = p_21_48 << 1;
  assign t_r22_c48_1 = p_22_47 << 1;
  assign t_r22_c48_2 = p_22_48 << 2;
  assign t_r22_c48_3 = p_22_49 << 1;
  assign t_r22_c48_4 = p_23_48 << 1;
  assign t_r22_c48_5 = t_r22_c48_0 + p_21_47;
  assign t_r22_c48_6 = t_r22_c48_1 + p_21_49;
  assign t_r22_c48_7 = t_r22_c48_2 + t_r22_c48_3;
  assign t_r22_c48_8 = t_r22_c48_4 + p_23_47;
  assign t_r22_c48_9 = t_r22_c48_5 + t_r22_c48_6;
  assign t_r22_c48_10 = t_r22_c48_7 + t_r22_c48_8;
  assign t_r22_c48_11 = t_r22_c48_9 + t_r22_c48_10;
  assign t_r22_c48_12 = t_r22_c48_11 + p_23_49;
  assign out_22_48 = t_r22_c48_12 >> 4;

  assign t_r22_c49_0 = p_21_49 << 1;
  assign t_r22_c49_1 = p_22_48 << 1;
  assign t_r22_c49_2 = p_22_49 << 2;
  assign t_r22_c49_3 = p_22_50 << 1;
  assign t_r22_c49_4 = p_23_49 << 1;
  assign t_r22_c49_5 = t_r22_c49_0 + p_21_48;
  assign t_r22_c49_6 = t_r22_c49_1 + p_21_50;
  assign t_r22_c49_7 = t_r22_c49_2 + t_r22_c49_3;
  assign t_r22_c49_8 = t_r22_c49_4 + p_23_48;
  assign t_r22_c49_9 = t_r22_c49_5 + t_r22_c49_6;
  assign t_r22_c49_10 = t_r22_c49_7 + t_r22_c49_8;
  assign t_r22_c49_11 = t_r22_c49_9 + t_r22_c49_10;
  assign t_r22_c49_12 = t_r22_c49_11 + p_23_50;
  assign out_22_49 = t_r22_c49_12 >> 4;

  assign t_r22_c50_0 = p_21_50 << 1;
  assign t_r22_c50_1 = p_22_49 << 1;
  assign t_r22_c50_2 = p_22_50 << 2;
  assign t_r22_c50_3 = p_22_51 << 1;
  assign t_r22_c50_4 = p_23_50 << 1;
  assign t_r22_c50_5 = t_r22_c50_0 + p_21_49;
  assign t_r22_c50_6 = t_r22_c50_1 + p_21_51;
  assign t_r22_c50_7 = t_r22_c50_2 + t_r22_c50_3;
  assign t_r22_c50_8 = t_r22_c50_4 + p_23_49;
  assign t_r22_c50_9 = t_r22_c50_5 + t_r22_c50_6;
  assign t_r22_c50_10 = t_r22_c50_7 + t_r22_c50_8;
  assign t_r22_c50_11 = t_r22_c50_9 + t_r22_c50_10;
  assign t_r22_c50_12 = t_r22_c50_11 + p_23_51;
  assign out_22_50 = t_r22_c50_12 >> 4;

  assign t_r22_c51_0 = p_21_51 << 1;
  assign t_r22_c51_1 = p_22_50 << 1;
  assign t_r22_c51_2 = p_22_51 << 2;
  assign t_r22_c51_3 = p_22_52 << 1;
  assign t_r22_c51_4 = p_23_51 << 1;
  assign t_r22_c51_5 = t_r22_c51_0 + p_21_50;
  assign t_r22_c51_6 = t_r22_c51_1 + p_21_52;
  assign t_r22_c51_7 = t_r22_c51_2 + t_r22_c51_3;
  assign t_r22_c51_8 = t_r22_c51_4 + p_23_50;
  assign t_r22_c51_9 = t_r22_c51_5 + t_r22_c51_6;
  assign t_r22_c51_10 = t_r22_c51_7 + t_r22_c51_8;
  assign t_r22_c51_11 = t_r22_c51_9 + t_r22_c51_10;
  assign t_r22_c51_12 = t_r22_c51_11 + p_23_52;
  assign out_22_51 = t_r22_c51_12 >> 4;

  assign t_r22_c52_0 = p_21_52 << 1;
  assign t_r22_c52_1 = p_22_51 << 1;
  assign t_r22_c52_2 = p_22_52 << 2;
  assign t_r22_c52_3 = p_22_53 << 1;
  assign t_r22_c52_4 = p_23_52 << 1;
  assign t_r22_c52_5 = t_r22_c52_0 + p_21_51;
  assign t_r22_c52_6 = t_r22_c52_1 + p_21_53;
  assign t_r22_c52_7 = t_r22_c52_2 + t_r22_c52_3;
  assign t_r22_c52_8 = t_r22_c52_4 + p_23_51;
  assign t_r22_c52_9 = t_r22_c52_5 + t_r22_c52_6;
  assign t_r22_c52_10 = t_r22_c52_7 + t_r22_c52_8;
  assign t_r22_c52_11 = t_r22_c52_9 + t_r22_c52_10;
  assign t_r22_c52_12 = t_r22_c52_11 + p_23_53;
  assign out_22_52 = t_r22_c52_12 >> 4;

  assign t_r22_c53_0 = p_21_53 << 1;
  assign t_r22_c53_1 = p_22_52 << 1;
  assign t_r22_c53_2 = p_22_53 << 2;
  assign t_r22_c53_3 = p_22_54 << 1;
  assign t_r22_c53_4 = p_23_53 << 1;
  assign t_r22_c53_5 = t_r22_c53_0 + p_21_52;
  assign t_r22_c53_6 = t_r22_c53_1 + p_21_54;
  assign t_r22_c53_7 = t_r22_c53_2 + t_r22_c53_3;
  assign t_r22_c53_8 = t_r22_c53_4 + p_23_52;
  assign t_r22_c53_9 = t_r22_c53_5 + t_r22_c53_6;
  assign t_r22_c53_10 = t_r22_c53_7 + t_r22_c53_8;
  assign t_r22_c53_11 = t_r22_c53_9 + t_r22_c53_10;
  assign t_r22_c53_12 = t_r22_c53_11 + p_23_54;
  assign out_22_53 = t_r22_c53_12 >> 4;

  assign t_r22_c54_0 = p_21_54 << 1;
  assign t_r22_c54_1 = p_22_53 << 1;
  assign t_r22_c54_2 = p_22_54 << 2;
  assign t_r22_c54_3 = p_22_55 << 1;
  assign t_r22_c54_4 = p_23_54 << 1;
  assign t_r22_c54_5 = t_r22_c54_0 + p_21_53;
  assign t_r22_c54_6 = t_r22_c54_1 + p_21_55;
  assign t_r22_c54_7 = t_r22_c54_2 + t_r22_c54_3;
  assign t_r22_c54_8 = t_r22_c54_4 + p_23_53;
  assign t_r22_c54_9 = t_r22_c54_5 + t_r22_c54_6;
  assign t_r22_c54_10 = t_r22_c54_7 + t_r22_c54_8;
  assign t_r22_c54_11 = t_r22_c54_9 + t_r22_c54_10;
  assign t_r22_c54_12 = t_r22_c54_11 + p_23_55;
  assign out_22_54 = t_r22_c54_12 >> 4;

  assign t_r22_c55_0 = p_21_55 << 1;
  assign t_r22_c55_1 = p_22_54 << 1;
  assign t_r22_c55_2 = p_22_55 << 2;
  assign t_r22_c55_3 = p_22_56 << 1;
  assign t_r22_c55_4 = p_23_55 << 1;
  assign t_r22_c55_5 = t_r22_c55_0 + p_21_54;
  assign t_r22_c55_6 = t_r22_c55_1 + p_21_56;
  assign t_r22_c55_7 = t_r22_c55_2 + t_r22_c55_3;
  assign t_r22_c55_8 = t_r22_c55_4 + p_23_54;
  assign t_r22_c55_9 = t_r22_c55_5 + t_r22_c55_6;
  assign t_r22_c55_10 = t_r22_c55_7 + t_r22_c55_8;
  assign t_r22_c55_11 = t_r22_c55_9 + t_r22_c55_10;
  assign t_r22_c55_12 = t_r22_c55_11 + p_23_56;
  assign out_22_55 = t_r22_c55_12 >> 4;

  assign t_r22_c56_0 = p_21_56 << 1;
  assign t_r22_c56_1 = p_22_55 << 1;
  assign t_r22_c56_2 = p_22_56 << 2;
  assign t_r22_c56_3 = p_22_57 << 1;
  assign t_r22_c56_4 = p_23_56 << 1;
  assign t_r22_c56_5 = t_r22_c56_0 + p_21_55;
  assign t_r22_c56_6 = t_r22_c56_1 + p_21_57;
  assign t_r22_c56_7 = t_r22_c56_2 + t_r22_c56_3;
  assign t_r22_c56_8 = t_r22_c56_4 + p_23_55;
  assign t_r22_c56_9 = t_r22_c56_5 + t_r22_c56_6;
  assign t_r22_c56_10 = t_r22_c56_7 + t_r22_c56_8;
  assign t_r22_c56_11 = t_r22_c56_9 + t_r22_c56_10;
  assign t_r22_c56_12 = t_r22_c56_11 + p_23_57;
  assign out_22_56 = t_r22_c56_12 >> 4;

  assign t_r22_c57_0 = p_21_57 << 1;
  assign t_r22_c57_1 = p_22_56 << 1;
  assign t_r22_c57_2 = p_22_57 << 2;
  assign t_r22_c57_3 = p_22_58 << 1;
  assign t_r22_c57_4 = p_23_57 << 1;
  assign t_r22_c57_5 = t_r22_c57_0 + p_21_56;
  assign t_r22_c57_6 = t_r22_c57_1 + p_21_58;
  assign t_r22_c57_7 = t_r22_c57_2 + t_r22_c57_3;
  assign t_r22_c57_8 = t_r22_c57_4 + p_23_56;
  assign t_r22_c57_9 = t_r22_c57_5 + t_r22_c57_6;
  assign t_r22_c57_10 = t_r22_c57_7 + t_r22_c57_8;
  assign t_r22_c57_11 = t_r22_c57_9 + t_r22_c57_10;
  assign t_r22_c57_12 = t_r22_c57_11 + p_23_58;
  assign out_22_57 = t_r22_c57_12 >> 4;

  assign t_r22_c58_0 = p_21_58 << 1;
  assign t_r22_c58_1 = p_22_57 << 1;
  assign t_r22_c58_2 = p_22_58 << 2;
  assign t_r22_c58_3 = p_22_59 << 1;
  assign t_r22_c58_4 = p_23_58 << 1;
  assign t_r22_c58_5 = t_r22_c58_0 + p_21_57;
  assign t_r22_c58_6 = t_r22_c58_1 + p_21_59;
  assign t_r22_c58_7 = t_r22_c58_2 + t_r22_c58_3;
  assign t_r22_c58_8 = t_r22_c58_4 + p_23_57;
  assign t_r22_c58_9 = t_r22_c58_5 + t_r22_c58_6;
  assign t_r22_c58_10 = t_r22_c58_7 + t_r22_c58_8;
  assign t_r22_c58_11 = t_r22_c58_9 + t_r22_c58_10;
  assign t_r22_c58_12 = t_r22_c58_11 + p_23_59;
  assign out_22_58 = t_r22_c58_12 >> 4;

  assign t_r22_c59_0 = p_21_59 << 1;
  assign t_r22_c59_1 = p_22_58 << 1;
  assign t_r22_c59_2 = p_22_59 << 2;
  assign t_r22_c59_3 = p_22_60 << 1;
  assign t_r22_c59_4 = p_23_59 << 1;
  assign t_r22_c59_5 = t_r22_c59_0 + p_21_58;
  assign t_r22_c59_6 = t_r22_c59_1 + p_21_60;
  assign t_r22_c59_7 = t_r22_c59_2 + t_r22_c59_3;
  assign t_r22_c59_8 = t_r22_c59_4 + p_23_58;
  assign t_r22_c59_9 = t_r22_c59_5 + t_r22_c59_6;
  assign t_r22_c59_10 = t_r22_c59_7 + t_r22_c59_8;
  assign t_r22_c59_11 = t_r22_c59_9 + t_r22_c59_10;
  assign t_r22_c59_12 = t_r22_c59_11 + p_23_60;
  assign out_22_59 = t_r22_c59_12 >> 4;

  assign t_r22_c60_0 = p_21_60 << 1;
  assign t_r22_c60_1 = p_22_59 << 1;
  assign t_r22_c60_2 = p_22_60 << 2;
  assign t_r22_c60_3 = p_22_61 << 1;
  assign t_r22_c60_4 = p_23_60 << 1;
  assign t_r22_c60_5 = t_r22_c60_0 + p_21_59;
  assign t_r22_c60_6 = t_r22_c60_1 + p_21_61;
  assign t_r22_c60_7 = t_r22_c60_2 + t_r22_c60_3;
  assign t_r22_c60_8 = t_r22_c60_4 + p_23_59;
  assign t_r22_c60_9 = t_r22_c60_5 + t_r22_c60_6;
  assign t_r22_c60_10 = t_r22_c60_7 + t_r22_c60_8;
  assign t_r22_c60_11 = t_r22_c60_9 + t_r22_c60_10;
  assign t_r22_c60_12 = t_r22_c60_11 + p_23_61;
  assign out_22_60 = t_r22_c60_12 >> 4;

  assign t_r22_c61_0 = p_21_61 << 1;
  assign t_r22_c61_1 = p_22_60 << 1;
  assign t_r22_c61_2 = p_22_61 << 2;
  assign t_r22_c61_3 = p_22_62 << 1;
  assign t_r22_c61_4 = p_23_61 << 1;
  assign t_r22_c61_5 = t_r22_c61_0 + p_21_60;
  assign t_r22_c61_6 = t_r22_c61_1 + p_21_62;
  assign t_r22_c61_7 = t_r22_c61_2 + t_r22_c61_3;
  assign t_r22_c61_8 = t_r22_c61_4 + p_23_60;
  assign t_r22_c61_9 = t_r22_c61_5 + t_r22_c61_6;
  assign t_r22_c61_10 = t_r22_c61_7 + t_r22_c61_8;
  assign t_r22_c61_11 = t_r22_c61_9 + t_r22_c61_10;
  assign t_r22_c61_12 = t_r22_c61_11 + p_23_62;
  assign out_22_61 = t_r22_c61_12 >> 4;

  assign t_r22_c62_0 = p_21_62 << 1;
  assign t_r22_c62_1 = p_22_61 << 1;
  assign t_r22_c62_2 = p_22_62 << 2;
  assign t_r22_c62_3 = p_22_63 << 1;
  assign t_r22_c62_4 = p_23_62 << 1;
  assign t_r22_c62_5 = t_r22_c62_0 + p_21_61;
  assign t_r22_c62_6 = t_r22_c62_1 + p_21_63;
  assign t_r22_c62_7 = t_r22_c62_2 + t_r22_c62_3;
  assign t_r22_c62_8 = t_r22_c62_4 + p_23_61;
  assign t_r22_c62_9 = t_r22_c62_5 + t_r22_c62_6;
  assign t_r22_c62_10 = t_r22_c62_7 + t_r22_c62_8;
  assign t_r22_c62_11 = t_r22_c62_9 + t_r22_c62_10;
  assign t_r22_c62_12 = t_r22_c62_11 + p_23_63;
  assign out_22_62 = t_r22_c62_12 >> 4;

  assign t_r22_c63_0 = p_21_63 << 1;
  assign t_r22_c63_1 = p_22_62 << 1;
  assign t_r22_c63_2 = p_22_63 << 2;
  assign t_r22_c63_3 = p_22_64 << 1;
  assign t_r22_c63_4 = p_23_63 << 1;
  assign t_r22_c63_5 = t_r22_c63_0 + p_21_62;
  assign t_r22_c63_6 = t_r22_c63_1 + p_21_64;
  assign t_r22_c63_7 = t_r22_c63_2 + t_r22_c63_3;
  assign t_r22_c63_8 = t_r22_c63_4 + p_23_62;
  assign t_r22_c63_9 = t_r22_c63_5 + t_r22_c63_6;
  assign t_r22_c63_10 = t_r22_c63_7 + t_r22_c63_8;
  assign t_r22_c63_11 = t_r22_c63_9 + t_r22_c63_10;
  assign t_r22_c63_12 = t_r22_c63_11 + p_23_64;
  assign out_22_63 = t_r22_c63_12 >> 4;

  assign t_r22_c64_0 = p_21_64 << 1;
  assign t_r22_c64_1 = p_22_63 << 1;
  assign t_r22_c64_2 = p_22_64 << 2;
  assign t_r22_c64_3 = p_22_65 << 1;
  assign t_r22_c64_4 = p_23_64 << 1;
  assign t_r22_c64_5 = t_r22_c64_0 + p_21_63;
  assign t_r22_c64_6 = t_r22_c64_1 + p_21_65;
  assign t_r22_c64_7 = t_r22_c64_2 + t_r22_c64_3;
  assign t_r22_c64_8 = t_r22_c64_4 + p_23_63;
  assign t_r22_c64_9 = t_r22_c64_5 + t_r22_c64_6;
  assign t_r22_c64_10 = t_r22_c64_7 + t_r22_c64_8;
  assign t_r22_c64_11 = t_r22_c64_9 + t_r22_c64_10;
  assign t_r22_c64_12 = t_r22_c64_11 + p_23_65;
  assign out_22_64 = t_r22_c64_12 >> 4;

  assign t_r23_c1_0 = p_22_1 << 1;
  assign t_r23_c1_1 = p_23_0 << 1;
  assign t_r23_c1_2 = p_23_1 << 2;
  assign t_r23_c1_3 = p_23_2 << 1;
  assign t_r23_c1_4 = p_24_1 << 1;
  assign t_r23_c1_5 = t_r23_c1_0 + p_22_0;
  assign t_r23_c1_6 = t_r23_c1_1 + p_22_2;
  assign t_r23_c1_7 = t_r23_c1_2 + t_r23_c1_3;
  assign t_r23_c1_8 = t_r23_c1_4 + p_24_0;
  assign t_r23_c1_9 = t_r23_c1_5 + t_r23_c1_6;
  assign t_r23_c1_10 = t_r23_c1_7 + t_r23_c1_8;
  assign t_r23_c1_11 = t_r23_c1_9 + t_r23_c1_10;
  assign t_r23_c1_12 = t_r23_c1_11 + p_24_2;
  assign out_23_1 = t_r23_c1_12 >> 4;

  assign t_r23_c2_0 = p_22_2 << 1;
  assign t_r23_c2_1 = p_23_1 << 1;
  assign t_r23_c2_2 = p_23_2 << 2;
  assign t_r23_c2_3 = p_23_3 << 1;
  assign t_r23_c2_4 = p_24_2 << 1;
  assign t_r23_c2_5 = t_r23_c2_0 + p_22_1;
  assign t_r23_c2_6 = t_r23_c2_1 + p_22_3;
  assign t_r23_c2_7 = t_r23_c2_2 + t_r23_c2_3;
  assign t_r23_c2_8 = t_r23_c2_4 + p_24_1;
  assign t_r23_c2_9 = t_r23_c2_5 + t_r23_c2_6;
  assign t_r23_c2_10 = t_r23_c2_7 + t_r23_c2_8;
  assign t_r23_c2_11 = t_r23_c2_9 + t_r23_c2_10;
  assign t_r23_c2_12 = t_r23_c2_11 + p_24_3;
  assign out_23_2 = t_r23_c2_12 >> 4;

  assign t_r23_c3_0 = p_22_3 << 1;
  assign t_r23_c3_1 = p_23_2 << 1;
  assign t_r23_c3_2 = p_23_3 << 2;
  assign t_r23_c3_3 = p_23_4 << 1;
  assign t_r23_c3_4 = p_24_3 << 1;
  assign t_r23_c3_5 = t_r23_c3_0 + p_22_2;
  assign t_r23_c3_6 = t_r23_c3_1 + p_22_4;
  assign t_r23_c3_7 = t_r23_c3_2 + t_r23_c3_3;
  assign t_r23_c3_8 = t_r23_c3_4 + p_24_2;
  assign t_r23_c3_9 = t_r23_c3_5 + t_r23_c3_6;
  assign t_r23_c3_10 = t_r23_c3_7 + t_r23_c3_8;
  assign t_r23_c3_11 = t_r23_c3_9 + t_r23_c3_10;
  assign t_r23_c3_12 = t_r23_c3_11 + p_24_4;
  assign out_23_3 = t_r23_c3_12 >> 4;

  assign t_r23_c4_0 = p_22_4 << 1;
  assign t_r23_c4_1 = p_23_3 << 1;
  assign t_r23_c4_2 = p_23_4 << 2;
  assign t_r23_c4_3 = p_23_5 << 1;
  assign t_r23_c4_4 = p_24_4 << 1;
  assign t_r23_c4_5 = t_r23_c4_0 + p_22_3;
  assign t_r23_c4_6 = t_r23_c4_1 + p_22_5;
  assign t_r23_c4_7 = t_r23_c4_2 + t_r23_c4_3;
  assign t_r23_c4_8 = t_r23_c4_4 + p_24_3;
  assign t_r23_c4_9 = t_r23_c4_5 + t_r23_c4_6;
  assign t_r23_c4_10 = t_r23_c4_7 + t_r23_c4_8;
  assign t_r23_c4_11 = t_r23_c4_9 + t_r23_c4_10;
  assign t_r23_c4_12 = t_r23_c4_11 + p_24_5;
  assign out_23_4 = t_r23_c4_12 >> 4;

  assign t_r23_c5_0 = p_22_5 << 1;
  assign t_r23_c5_1 = p_23_4 << 1;
  assign t_r23_c5_2 = p_23_5 << 2;
  assign t_r23_c5_3 = p_23_6 << 1;
  assign t_r23_c5_4 = p_24_5 << 1;
  assign t_r23_c5_5 = t_r23_c5_0 + p_22_4;
  assign t_r23_c5_6 = t_r23_c5_1 + p_22_6;
  assign t_r23_c5_7 = t_r23_c5_2 + t_r23_c5_3;
  assign t_r23_c5_8 = t_r23_c5_4 + p_24_4;
  assign t_r23_c5_9 = t_r23_c5_5 + t_r23_c5_6;
  assign t_r23_c5_10 = t_r23_c5_7 + t_r23_c5_8;
  assign t_r23_c5_11 = t_r23_c5_9 + t_r23_c5_10;
  assign t_r23_c5_12 = t_r23_c5_11 + p_24_6;
  assign out_23_5 = t_r23_c5_12 >> 4;

  assign t_r23_c6_0 = p_22_6 << 1;
  assign t_r23_c6_1 = p_23_5 << 1;
  assign t_r23_c6_2 = p_23_6 << 2;
  assign t_r23_c6_3 = p_23_7 << 1;
  assign t_r23_c6_4 = p_24_6 << 1;
  assign t_r23_c6_5 = t_r23_c6_0 + p_22_5;
  assign t_r23_c6_6 = t_r23_c6_1 + p_22_7;
  assign t_r23_c6_7 = t_r23_c6_2 + t_r23_c6_3;
  assign t_r23_c6_8 = t_r23_c6_4 + p_24_5;
  assign t_r23_c6_9 = t_r23_c6_5 + t_r23_c6_6;
  assign t_r23_c6_10 = t_r23_c6_7 + t_r23_c6_8;
  assign t_r23_c6_11 = t_r23_c6_9 + t_r23_c6_10;
  assign t_r23_c6_12 = t_r23_c6_11 + p_24_7;
  assign out_23_6 = t_r23_c6_12 >> 4;

  assign t_r23_c7_0 = p_22_7 << 1;
  assign t_r23_c7_1 = p_23_6 << 1;
  assign t_r23_c7_2 = p_23_7 << 2;
  assign t_r23_c7_3 = p_23_8 << 1;
  assign t_r23_c7_4 = p_24_7 << 1;
  assign t_r23_c7_5 = t_r23_c7_0 + p_22_6;
  assign t_r23_c7_6 = t_r23_c7_1 + p_22_8;
  assign t_r23_c7_7 = t_r23_c7_2 + t_r23_c7_3;
  assign t_r23_c7_8 = t_r23_c7_4 + p_24_6;
  assign t_r23_c7_9 = t_r23_c7_5 + t_r23_c7_6;
  assign t_r23_c7_10 = t_r23_c7_7 + t_r23_c7_8;
  assign t_r23_c7_11 = t_r23_c7_9 + t_r23_c7_10;
  assign t_r23_c7_12 = t_r23_c7_11 + p_24_8;
  assign out_23_7 = t_r23_c7_12 >> 4;

  assign t_r23_c8_0 = p_22_8 << 1;
  assign t_r23_c8_1 = p_23_7 << 1;
  assign t_r23_c8_2 = p_23_8 << 2;
  assign t_r23_c8_3 = p_23_9 << 1;
  assign t_r23_c8_4 = p_24_8 << 1;
  assign t_r23_c8_5 = t_r23_c8_0 + p_22_7;
  assign t_r23_c8_6 = t_r23_c8_1 + p_22_9;
  assign t_r23_c8_7 = t_r23_c8_2 + t_r23_c8_3;
  assign t_r23_c8_8 = t_r23_c8_4 + p_24_7;
  assign t_r23_c8_9 = t_r23_c8_5 + t_r23_c8_6;
  assign t_r23_c8_10 = t_r23_c8_7 + t_r23_c8_8;
  assign t_r23_c8_11 = t_r23_c8_9 + t_r23_c8_10;
  assign t_r23_c8_12 = t_r23_c8_11 + p_24_9;
  assign out_23_8 = t_r23_c8_12 >> 4;

  assign t_r23_c9_0 = p_22_9 << 1;
  assign t_r23_c9_1 = p_23_8 << 1;
  assign t_r23_c9_2 = p_23_9 << 2;
  assign t_r23_c9_3 = p_23_10 << 1;
  assign t_r23_c9_4 = p_24_9 << 1;
  assign t_r23_c9_5 = t_r23_c9_0 + p_22_8;
  assign t_r23_c9_6 = t_r23_c9_1 + p_22_10;
  assign t_r23_c9_7 = t_r23_c9_2 + t_r23_c9_3;
  assign t_r23_c9_8 = t_r23_c9_4 + p_24_8;
  assign t_r23_c9_9 = t_r23_c9_5 + t_r23_c9_6;
  assign t_r23_c9_10 = t_r23_c9_7 + t_r23_c9_8;
  assign t_r23_c9_11 = t_r23_c9_9 + t_r23_c9_10;
  assign t_r23_c9_12 = t_r23_c9_11 + p_24_10;
  assign out_23_9 = t_r23_c9_12 >> 4;

  assign t_r23_c10_0 = p_22_10 << 1;
  assign t_r23_c10_1 = p_23_9 << 1;
  assign t_r23_c10_2 = p_23_10 << 2;
  assign t_r23_c10_3 = p_23_11 << 1;
  assign t_r23_c10_4 = p_24_10 << 1;
  assign t_r23_c10_5 = t_r23_c10_0 + p_22_9;
  assign t_r23_c10_6 = t_r23_c10_1 + p_22_11;
  assign t_r23_c10_7 = t_r23_c10_2 + t_r23_c10_3;
  assign t_r23_c10_8 = t_r23_c10_4 + p_24_9;
  assign t_r23_c10_9 = t_r23_c10_5 + t_r23_c10_6;
  assign t_r23_c10_10 = t_r23_c10_7 + t_r23_c10_8;
  assign t_r23_c10_11 = t_r23_c10_9 + t_r23_c10_10;
  assign t_r23_c10_12 = t_r23_c10_11 + p_24_11;
  assign out_23_10 = t_r23_c10_12 >> 4;

  assign t_r23_c11_0 = p_22_11 << 1;
  assign t_r23_c11_1 = p_23_10 << 1;
  assign t_r23_c11_2 = p_23_11 << 2;
  assign t_r23_c11_3 = p_23_12 << 1;
  assign t_r23_c11_4 = p_24_11 << 1;
  assign t_r23_c11_5 = t_r23_c11_0 + p_22_10;
  assign t_r23_c11_6 = t_r23_c11_1 + p_22_12;
  assign t_r23_c11_7 = t_r23_c11_2 + t_r23_c11_3;
  assign t_r23_c11_8 = t_r23_c11_4 + p_24_10;
  assign t_r23_c11_9 = t_r23_c11_5 + t_r23_c11_6;
  assign t_r23_c11_10 = t_r23_c11_7 + t_r23_c11_8;
  assign t_r23_c11_11 = t_r23_c11_9 + t_r23_c11_10;
  assign t_r23_c11_12 = t_r23_c11_11 + p_24_12;
  assign out_23_11 = t_r23_c11_12 >> 4;

  assign t_r23_c12_0 = p_22_12 << 1;
  assign t_r23_c12_1 = p_23_11 << 1;
  assign t_r23_c12_2 = p_23_12 << 2;
  assign t_r23_c12_3 = p_23_13 << 1;
  assign t_r23_c12_4 = p_24_12 << 1;
  assign t_r23_c12_5 = t_r23_c12_0 + p_22_11;
  assign t_r23_c12_6 = t_r23_c12_1 + p_22_13;
  assign t_r23_c12_7 = t_r23_c12_2 + t_r23_c12_3;
  assign t_r23_c12_8 = t_r23_c12_4 + p_24_11;
  assign t_r23_c12_9 = t_r23_c12_5 + t_r23_c12_6;
  assign t_r23_c12_10 = t_r23_c12_7 + t_r23_c12_8;
  assign t_r23_c12_11 = t_r23_c12_9 + t_r23_c12_10;
  assign t_r23_c12_12 = t_r23_c12_11 + p_24_13;
  assign out_23_12 = t_r23_c12_12 >> 4;

  assign t_r23_c13_0 = p_22_13 << 1;
  assign t_r23_c13_1 = p_23_12 << 1;
  assign t_r23_c13_2 = p_23_13 << 2;
  assign t_r23_c13_3 = p_23_14 << 1;
  assign t_r23_c13_4 = p_24_13 << 1;
  assign t_r23_c13_5 = t_r23_c13_0 + p_22_12;
  assign t_r23_c13_6 = t_r23_c13_1 + p_22_14;
  assign t_r23_c13_7 = t_r23_c13_2 + t_r23_c13_3;
  assign t_r23_c13_8 = t_r23_c13_4 + p_24_12;
  assign t_r23_c13_9 = t_r23_c13_5 + t_r23_c13_6;
  assign t_r23_c13_10 = t_r23_c13_7 + t_r23_c13_8;
  assign t_r23_c13_11 = t_r23_c13_9 + t_r23_c13_10;
  assign t_r23_c13_12 = t_r23_c13_11 + p_24_14;
  assign out_23_13 = t_r23_c13_12 >> 4;

  assign t_r23_c14_0 = p_22_14 << 1;
  assign t_r23_c14_1 = p_23_13 << 1;
  assign t_r23_c14_2 = p_23_14 << 2;
  assign t_r23_c14_3 = p_23_15 << 1;
  assign t_r23_c14_4 = p_24_14 << 1;
  assign t_r23_c14_5 = t_r23_c14_0 + p_22_13;
  assign t_r23_c14_6 = t_r23_c14_1 + p_22_15;
  assign t_r23_c14_7 = t_r23_c14_2 + t_r23_c14_3;
  assign t_r23_c14_8 = t_r23_c14_4 + p_24_13;
  assign t_r23_c14_9 = t_r23_c14_5 + t_r23_c14_6;
  assign t_r23_c14_10 = t_r23_c14_7 + t_r23_c14_8;
  assign t_r23_c14_11 = t_r23_c14_9 + t_r23_c14_10;
  assign t_r23_c14_12 = t_r23_c14_11 + p_24_15;
  assign out_23_14 = t_r23_c14_12 >> 4;

  assign t_r23_c15_0 = p_22_15 << 1;
  assign t_r23_c15_1 = p_23_14 << 1;
  assign t_r23_c15_2 = p_23_15 << 2;
  assign t_r23_c15_3 = p_23_16 << 1;
  assign t_r23_c15_4 = p_24_15 << 1;
  assign t_r23_c15_5 = t_r23_c15_0 + p_22_14;
  assign t_r23_c15_6 = t_r23_c15_1 + p_22_16;
  assign t_r23_c15_7 = t_r23_c15_2 + t_r23_c15_3;
  assign t_r23_c15_8 = t_r23_c15_4 + p_24_14;
  assign t_r23_c15_9 = t_r23_c15_5 + t_r23_c15_6;
  assign t_r23_c15_10 = t_r23_c15_7 + t_r23_c15_8;
  assign t_r23_c15_11 = t_r23_c15_9 + t_r23_c15_10;
  assign t_r23_c15_12 = t_r23_c15_11 + p_24_16;
  assign out_23_15 = t_r23_c15_12 >> 4;

  assign t_r23_c16_0 = p_22_16 << 1;
  assign t_r23_c16_1 = p_23_15 << 1;
  assign t_r23_c16_2 = p_23_16 << 2;
  assign t_r23_c16_3 = p_23_17 << 1;
  assign t_r23_c16_4 = p_24_16 << 1;
  assign t_r23_c16_5 = t_r23_c16_0 + p_22_15;
  assign t_r23_c16_6 = t_r23_c16_1 + p_22_17;
  assign t_r23_c16_7 = t_r23_c16_2 + t_r23_c16_3;
  assign t_r23_c16_8 = t_r23_c16_4 + p_24_15;
  assign t_r23_c16_9 = t_r23_c16_5 + t_r23_c16_6;
  assign t_r23_c16_10 = t_r23_c16_7 + t_r23_c16_8;
  assign t_r23_c16_11 = t_r23_c16_9 + t_r23_c16_10;
  assign t_r23_c16_12 = t_r23_c16_11 + p_24_17;
  assign out_23_16 = t_r23_c16_12 >> 4;

  assign t_r23_c17_0 = p_22_17 << 1;
  assign t_r23_c17_1 = p_23_16 << 1;
  assign t_r23_c17_2 = p_23_17 << 2;
  assign t_r23_c17_3 = p_23_18 << 1;
  assign t_r23_c17_4 = p_24_17 << 1;
  assign t_r23_c17_5 = t_r23_c17_0 + p_22_16;
  assign t_r23_c17_6 = t_r23_c17_1 + p_22_18;
  assign t_r23_c17_7 = t_r23_c17_2 + t_r23_c17_3;
  assign t_r23_c17_8 = t_r23_c17_4 + p_24_16;
  assign t_r23_c17_9 = t_r23_c17_5 + t_r23_c17_6;
  assign t_r23_c17_10 = t_r23_c17_7 + t_r23_c17_8;
  assign t_r23_c17_11 = t_r23_c17_9 + t_r23_c17_10;
  assign t_r23_c17_12 = t_r23_c17_11 + p_24_18;
  assign out_23_17 = t_r23_c17_12 >> 4;

  assign t_r23_c18_0 = p_22_18 << 1;
  assign t_r23_c18_1 = p_23_17 << 1;
  assign t_r23_c18_2 = p_23_18 << 2;
  assign t_r23_c18_3 = p_23_19 << 1;
  assign t_r23_c18_4 = p_24_18 << 1;
  assign t_r23_c18_5 = t_r23_c18_0 + p_22_17;
  assign t_r23_c18_6 = t_r23_c18_1 + p_22_19;
  assign t_r23_c18_7 = t_r23_c18_2 + t_r23_c18_3;
  assign t_r23_c18_8 = t_r23_c18_4 + p_24_17;
  assign t_r23_c18_9 = t_r23_c18_5 + t_r23_c18_6;
  assign t_r23_c18_10 = t_r23_c18_7 + t_r23_c18_8;
  assign t_r23_c18_11 = t_r23_c18_9 + t_r23_c18_10;
  assign t_r23_c18_12 = t_r23_c18_11 + p_24_19;
  assign out_23_18 = t_r23_c18_12 >> 4;

  assign t_r23_c19_0 = p_22_19 << 1;
  assign t_r23_c19_1 = p_23_18 << 1;
  assign t_r23_c19_2 = p_23_19 << 2;
  assign t_r23_c19_3 = p_23_20 << 1;
  assign t_r23_c19_4 = p_24_19 << 1;
  assign t_r23_c19_5 = t_r23_c19_0 + p_22_18;
  assign t_r23_c19_6 = t_r23_c19_1 + p_22_20;
  assign t_r23_c19_7 = t_r23_c19_2 + t_r23_c19_3;
  assign t_r23_c19_8 = t_r23_c19_4 + p_24_18;
  assign t_r23_c19_9 = t_r23_c19_5 + t_r23_c19_6;
  assign t_r23_c19_10 = t_r23_c19_7 + t_r23_c19_8;
  assign t_r23_c19_11 = t_r23_c19_9 + t_r23_c19_10;
  assign t_r23_c19_12 = t_r23_c19_11 + p_24_20;
  assign out_23_19 = t_r23_c19_12 >> 4;

  assign t_r23_c20_0 = p_22_20 << 1;
  assign t_r23_c20_1 = p_23_19 << 1;
  assign t_r23_c20_2 = p_23_20 << 2;
  assign t_r23_c20_3 = p_23_21 << 1;
  assign t_r23_c20_4 = p_24_20 << 1;
  assign t_r23_c20_5 = t_r23_c20_0 + p_22_19;
  assign t_r23_c20_6 = t_r23_c20_1 + p_22_21;
  assign t_r23_c20_7 = t_r23_c20_2 + t_r23_c20_3;
  assign t_r23_c20_8 = t_r23_c20_4 + p_24_19;
  assign t_r23_c20_9 = t_r23_c20_5 + t_r23_c20_6;
  assign t_r23_c20_10 = t_r23_c20_7 + t_r23_c20_8;
  assign t_r23_c20_11 = t_r23_c20_9 + t_r23_c20_10;
  assign t_r23_c20_12 = t_r23_c20_11 + p_24_21;
  assign out_23_20 = t_r23_c20_12 >> 4;

  assign t_r23_c21_0 = p_22_21 << 1;
  assign t_r23_c21_1 = p_23_20 << 1;
  assign t_r23_c21_2 = p_23_21 << 2;
  assign t_r23_c21_3 = p_23_22 << 1;
  assign t_r23_c21_4 = p_24_21 << 1;
  assign t_r23_c21_5 = t_r23_c21_0 + p_22_20;
  assign t_r23_c21_6 = t_r23_c21_1 + p_22_22;
  assign t_r23_c21_7 = t_r23_c21_2 + t_r23_c21_3;
  assign t_r23_c21_8 = t_r23_c21_4 + p_24_20;
  assign t_r23_c21_9 = t_r23_c21_5 + t_r23_c21_6;
  assign t_r23_c21_10 = t_r23_c21_7 + t_r23_c21_8;
  assign t_r23_c21_11 = t_r23_c21_9 + t_r23_c21_10;
  assign t_r23_c21_12 = t_r23_c21_11 + p_24_22;
  assign out_23_21 = t_r23_c21_12 >> 4;

  assign t_r23_c22_0 = p_22_22 << 1;
  assign t_r23_c22_1 = p_23_21 << 1;
  assign t_r23_c22_2 = p_23_22 << 2;
  assign t_r23_c22_3 = p_23_23 << 1;
  assign t_r23_c22_4 = p_24_22 << 1;
  assign t_r23_c22_5 = t_r23_c22_0 + p_22_21;
  assign t_r23_c22_6 = t_r23_c22_1 + p_22_23;
  assign t_r23_c22_7 = t_r23_c22_2 + t_r23_c22_3;
  assign t_r23_c22_8 = t_r23_c22_4 + p_24_21;
  assign t_r23_c22_9 = t_r23_c22_5 + t_r23_c22_6;
  assign t_r23_c22_10 = t_r23_c22_7 + t_r23_c22_8;
  assign t_r23_c22_11 = t_r23_c22_9 + t_r23_c22_10;
  assign t_r23_c22_12 = t_r23_c22_11 + p_24_23;
  assign out_23_22 = t_r23_c22_12 >> 4;

  assign t_r23_c23_0 = p_22_23 << 1;
  assign t_r23_c23_1 = p_23_22 << 1;
  assign t_r23_c23_2 = p_23_23 << 2;
  assign t_r23_c23_3 = p_23_24 << 1;
  assign t_r23_c23_4 = p_24_23 << 1;
  assign t_r23_c23_5 = t_r23_c23_0 + p_22_22;
  assign t_r23_c23_6 = t_r23_c23_1 + p_22_24;
  assign t_r23_c23_7 = t_r23_c23_2 + t_r23_c23_3;
  assign t_r23_c23_8 = t_r23_c23_4 + p_24_22;
  assign t_r23_c23_9 = t_r23_c23_5 + t_r23_c23_6;
  assign t_r23_c23_10 = t_r23_c23_7 + t_r23_c23_8;
  assign t_r23_c23_11 = t_r23_c23_9 + t_r23_c23_10;
  assign t_r23_c23_12 = t_r23_c23_11 + p_24_24;
  assign out_23_23 = t_r23_c23_12 >> 4;

  assign t_r23_c24_0 = p_22_24 << 1;
  assign t_r23_c24_1 = p_23_23 << 1;
  assign t_r23_c24_2 = p_23_24 << 2;
  assign t_r23_c24_3 = p_23_25 << 1;
  assign t_r23_c24_4 = p_24_24 << 1;
  assign t_r23_c24_5 = t_r23_c24_0 + p_22_23;
  assign t_r23_c24_6 = t_r23_c24_1 + p_22_25;
  assign t_r23_c24_7 = t_r23_c24_2 + t_r23_c24_3;
  assign t_r23_c24_8 = t_r23_c24_4 + p_24_23;
  assign t_r23_c24_9 = t_r23_c24_5 + t_r23_c24_6;
  assign t_r23_c24_10 = t_r23_c24_7 + t_r23_c24_8;
  assign t_r23_c24_11 = t_r23_c24_9 + t_r23_c24_10;
  assign t_r23_c24_12 = t_r23_c24_11 + p_24_25;
  assign out_23_24 = t_r23_c24_12 >> 4;

  assign t_r23_c25_0 = p_22_25 << 1;
  assign t_r23_c25_1 = p_23_24 << 1;
  assign t_r23_c25_2 = p_23_25 << 2;
  assign t_r23_c25_3 = p_23_26 << 1;
  assign t_r23_c25_4 = p_24_25 << 1;
  assign t_r23_c25_5 = t_r23_c25_0 + p_22_24;
  assign t_r23_c25_6 = t_r23_c25_1 + p_22_26;
  assign t_r23_c25_7 = t_r23_c25_2 + t_r23_c25_3;
  assign t_r23_c25_8 = t_r23_c25_4 + p_24_24;
  assign t_r23_c25_9 = t_r23_c25_5 + t_r23_c25_6;
  assign t_r23_c25_10 = t_r23_c25_7 + t_r23_c25_8;
  assign t_r23_c25_11 = t_r23_c25_9 + t_r23_c25_10;
  assign t_r23_c25_12 = t_r23_c25_11 + p_24_26;
  assign out_23_25 = t_r23_c25_12 >> 4;

  assign t_r23_c26_0 = p_22_26 << 1;
  assign t_r23_c26_1 = p_23_25 << 1;
  assign t_r23_c26_2 = p_23_26 << 2;
  assign t_r23_c26_3 = p_23_27 << 1;
  assign t_r23_c26_4 = p_24_26 << 1;
  assign t_r23_c26_5 = t_r23_c26_0 + p_22_25;
  assign t_r23_c26_6 = t_r23_c26_1 + p_22_27;
  assign t_r23_c26_7 = t_r23_c26_2 + t_r23_c26_3;
  assign t_r23_c26_8 = t_r23_c26_4 + p_24_25;
  assign t_r23_c26_9 = t_r23_c26_5 + t_r23_c26_6;
  assign t_r23_c26_10 = t_r23_c26_7 + t_r23_c26_8;
  assign t_r23_c26_11 = t_r23_c26_9 + t_r23_c26_10;
  assign t_r23_c26_12 = t_r23_c26_11 + p_24_27;
  assign out_23_26 = t_r23_c26_12 >> 4;

  assign t_r23_c27_0 = p_22_27 << 1;
  assign t_r23_c27_1 = p_23_26 << 1;
  assign t_r23_c27_2 = p_23_27 << 2;
  assign t_r23_c27_3 = p_23_28 << 1;
  assign t_r23_c27_4 = p_24_27 << 1;
  assign t_r23_c27_5 = t_r23_c27_0 + p_22_26;
  assign t_r23_c27_6 = t_r23_c27_1 + p_22_28;
  assign t_r23_c27_7 = t_r23_c27_2 + t_r23_c27_3;
  assign t_r23_c27_8 = t_r23_c27_4 + p_24_26;
  assign t_r23_c27_9 = t_r23_c27_5 + t_r23_c27_6;
  assign t_r23_c27_10 = t_r23_c27_7 + t_r23_c27_8;
  assign t_r23_c27_11 = t_r23_c27_9 + t_r23_c27_10;
  assign t_r23_c27_12 = t_r23_c27_11 + p_24_28;
  assign out_23_27 = t_r23_c27_12 >> 4;

  assign t_r23_c28_0 = p_22_28 << 1;
  assign t_r23_c28_1 = p_23_27 << 1;
  assign t_r23_c28_2 = p_23_28 << 2;
  assign t_r23_c28_3 = p_23_29 << 1;
  assign t_r23_c28_4 = p_24_28 << 1;
  assign t_r23_c28_5 = t_r23_c28_0 + p_22_27;
  assign t_r23_c28_6 = t_r23_c28_1 + p_22_29;
  assign t_r23_c28_7 = t_r23_c28_2 + t_r23_c28_3;
  assign t_r23_c28_8 = t_r23_c28_4 + p_24_27;
  assign t_r23_c28_9 = t_r23_c28_5 + t_r23_c28_6;
  assign t_r23_c28_10 = t_r23_c28_7 + t_r23_c28_8;
  assign t_r23_c28_11 = t_r23_c28_9 + t_r23_c28_10;
  assign t_r23_c28_12 = t_r23_c28_11 + p_24_29;
  assign out_23_28 = t_r23_c28_12 >> 4;

  assign t_r23_c29_0 = p_22_29 << 1;
  assign t_r23_c29_1 = p_23_28 << 1;
  assign t_r23_c29_2 = p_23_29 << 2;
  assign t_r23_c29_3 = p_23_30 << 1;
  assign t_r23_c29_4 = p_24_29 << 1;
  assign t_r23_c29_5 = t_r23_c29_0 + p_22_28;
  assign t_r23_c29_6 = t_r23_c29_1 + p_22_30;
  assign t_r23_c29_7 = t_r23_c29_2 + t_r23_c29_3;
  assign t_r23_c29_8 = t_r23_c29_4 + p_24_28;
  assign t_r23_c29_9 = t_r23_c29_5 + t_r23_c29_6;
  assign t_r23_c29_10 = t_r23_c29_7 + t_r23_c29_8;
  assign t_r23_c29_11 = t_r23_c29_9 + t_r23_c29_10;
  assign t_r23_c29_12 = t_r23_c29_11 + p_24_30;
  assign out_23_29 = t_r23_c29_12 >> 4;

  assign t_r23_c30_0 = p_22_30 << 1;
  assign t_r23_c30_1 = p_23_29 << 1;
  assign t_r23_c30_2 = p_23_30 << 2;
  assign t_r23_c30_3 = p_23_31 << 1;
  assign t_r23_c30_4 = p_24_30 << 1;
  assign t_r23_c30_5 = t_r23_c30_0 + p_22_29;
  assign t_r23_c30_6 = t_r23_c30_1 + p_22_31;
  assign t_r23_c30_7 = t_r23_c30_2 + t_r23_c30_3;
  assign t_r23_c30_8 = t_r23_c30_4 + p_24_29;
  assign t_r23_c30_9 = t_r23_c30_5 + t_r23_c30_6;
  assign t_r23_c30_10 = t_r23_c30_7 + t_r23_c30_8;
  assign t_r23_c30_11 = t_r23_c30_9 + t_r23_c30_10;
  assign t_r23_c30_12 = t_r23_c30_11 + p_24_31;
  assign out_23_30 = t_r23_c30_12 >> 4;

  assign t_r23_c31_0 = p_22_31 << 1;
  assign t_r23_c31_1 = p_23_30 << 1;
  assign t_r23_c31_2 = p_23_31 << 2;
  assign t_r23_c31_3 = p_23_32 << 1;
  assign t_r23_c31_4 = p_24_31 << 1;
  assign t_r23_c31_5 = t_r23_c31_0 + p_22_30;
  assign t_r23_c31_6 = t_r23_c31_1 + p_22_32;
  assign t_r23_c31_7 = t_r23_c31_2 + t_r23_c31_3;
  assign t_r23_c31_8 = t_r23_c31_4 + p_24_30;
  assign t_r23_c31_9 = t_r23_c31_5 + t_r23_c31_6;
  assign t_r23_c31_10 = t_r23_c31_7 + t_r23_c31_8;
  assign t_r23_c31_11 = t_r23_c31_9 + t_r23_c31_10;
  assign t_r23_c31_12 = t_r23_c31_11 + p_24_32;
  assign out_23_31 = t_r23_c31_12 >> 4;

  assign t_r23_c32_0 = p_22_32 << 1;
  assign t_r23_c32_1 = p_23_31 << 1;
  assign t_r23_c32_2 = p_23_32 << 2;
  assign t_r23_c32_3 = p_23_33 << 1;
  assign t_r23_c32_4 = p_24_32 << 1;
  assign t_r23_c32_5 = t_r23_c32_0 + p_22_31;
  assign t_r23_c32_6 = t_r23_c32_1 + p_22_33;
  assign t_r23_c32_7 = t_r23_c32_2 + t_r23_c32_3;
  assign t_r23_c32_8 = t_r23_c32_4 + p_24_31;
  assign t_r23_c32_9 = t_r23_c32_5 + t_r23_c32_6;
  assign t_r23_c32_10 = t_r23_c32_7 + t_r23_c32_8;
  assign t_r23_c32_11 = t_r23_c32_9 + t_r23_c32_10;
  assign t_r23_c32_12 = t_r23_c32_11 + p_24_33;
  assign out_23_32 = t_r23_c32_12 >> 4;

  assign t_r23_c33_0 = p_22_33 << 1;
  assign t_r23_c33_1 = p_23_32 << 1;
  assign t_r23_c33_2 = p_23_33 << 2;
  assign t_r23_c33_3 = p_23_34 << 1;
  assign t_r23_c33_4 = p_24_33 << 1;
  assign t_r23_c33_5 = t_r23_c33_0 + p_22_32;
  assign t_r23_c33_6 = t_r23_c33_1 + p_22_34;
  assign t_r23_c33_7 = t_r23_c33_2 + t_r23_c33_3;
  assign t_r23_c33_8 = t_r23_c33_4 + p_24_32;
  assign t_r23_c33_9 = t_r23_c33_5 + t_r23_c33_6;
  assign t_r23_c33_10 = t_r23_c33_7 + t_r23_c33_8;
  assign t_r23_c33_11 = t_r23_c33_9 + t_r23_c33_10;
  assign t_r23_c33_12 = t_r23_c33_11 + p_24_34;
  assign out_23_33 = t_r23_c33_12 >> 4;

  assign t_r23_c34_0 = p_22_34 << 1;
  assign t_r23_c34_1 = p_23_33 << 1;
  assign t_r23_c34_2 = p_23_34 << 2;
  assign t_r23_c34_3 = p_23_35 << 1;
  assign t_r23_c34_4 = p_24_34 << 1;
  assign t_r23_c34_5 = t_r23_c34_0 + p_22_33;
  assign t_r23_c34_6 = t_r23_c34_1 + p_22_35;
  assign t_r23_c34_7 = t_r23_c34_2 + t_r23_c34_3;
  assign t_r23_c34_8 = t_r23_c34_4 + p_24_33;
  assign t_r23_c34_9 = t_r23_c34_5 + t_r23_c34_6;
  assign t_r23_c34_10 = t_r23_c34_7 + t_r23_c34_8;
  assign t_r23_c34_11 = t_r23_c34_9 + t_r23_c34_10;
  assign t_r23_c34_12 = t_r23_c34_11 + p_24_35;
  assign out_23_34 = t_r23_c34_12 >> 4;

  assign t_r23_c35_0 = p_22_35 << 1;
  assign t_r23_c35_1 = p_23_34 << 1;
  assign t_r23_c35_2 = p_23_35 << 2;
  assign t_r23_c35_3 = p_23_36 << 1;
  assign t_r23_c35_4 = p_24_35 << 1;
  assign t_r23_c35_5 = t_r23_c35_0 + p_22_34;
  assign t_r23_c35_6 = t_r23_c35_1 + p_22_36;
  assign t_r23_c35_7 = t_r23_c35_2 + t_r23_c35_3;
  assign t_r23_c35_8 = t_r23_c35_4 + p_24_34;
  assign t_r23_c35_9 = t_r23_c35_5 + t_r23_c35_6;
  assign t_r23_c35_10 = t_r23_c35_7 + t_r23_c35_8;
  assign t_r23_c35_11 = t_r23_c35_9 + t_r23_c35_10;
  assign t_r23_c35_12 = t_r23_c35_11 + p_24_36;
  assign out_23_35 = t_r23_c35_12 >> 4;

  assign t_r23_c36_0 = p_22_36 << 1;
  assign t_r23_c36_1 = p_23_35 << 1;
  assign t_r23_c36_2 = p_23_36 << 2;
  assign t_r23_c36_3 = p_23_37 << 1;
  assign t_r23_c36_4 = p_24_36 << 1;
  assign t_r23_c36_5 = t_r23_c36_0 + p_22_35;
  assign t_r23_c36_6 = t_r23_c36_1 + p_22_37;
  assign t_r23_c36_7 = t_r23_c36_2 + t_r23_c36_3;
  assign t_r23_c36_8 = t_r23_c36_4 + p_24_35;
  assign t_r23_c36_9 = t_r23_c36_5 + t_r23_c36_6;
  assign t_r23_c36_10 = t_r23_c36_7 + t_r23_c36_8;
  assign t_r23_c36_11 = t_r23_c36_9 + t_r23_c36_10;
  assign t_r23_c36_12 = t_r23_c36_11 + p_24_37;
  assign out_23_36 = t_r23_c36_12 >> 4;

  assign t_r23_c37_0 = p_22_37 << 1;
  assign t_r23_c37_1 = p_23_36 << 1;
  assign t_r23_c37_2 = p_23_37 << 2;
  assign t_r23_c37_3 = p_23_38 << 1;
  assign t_r23_c37_4 = p_24_37 << 1;
  assign t_r23_c37_5 = t_r23_c37_0 + p_22_36;
  assign t_r23_c37_6 = t_r23_c37_1 + p_22_38;
  assign t_r23_c37_7 = t_r23_c37_2 + t_r23_c37_3;
  assign t_r23_c37_8 = t_r23_c37_4 + p_24_36;
  assign t_r23_c37_9 = t_r23_c37_5 + t_r23_c37_6;
  assign t_r23_c37_10 = t_r23_c37_7 + t_r23_c37_8;
  assign t_r23_c37_11 = t_r23_c37_9 + t_r23_c37_10;
  assign t_r23_c37_12 = t_r23_c37_11 + p_24_38;
  assign out_23_37 = t_r23_c37_12 >> 4;

  assign t_r23_c38_0 = p_22_38 << 1;
  assign t_r23_c38_1 = p_23_37 << 1;
  assign t_r23_c38_2 = p_23_38 << 2;
  assign t_r23_c38_3 = p_23_39 << 1;
  assign t_r23_c38_4 = p_24_38 << 1;
  assign t_r23_c38_5 = t_r23_c38_0 + p_22_37;
  assign t_r23_c38_6 = t_r23_c38_1 + p_22_39;
  assign t_r23_c38_7 = t_r23_c38_2 + t_r23_c38_3;
  assign t_r23_c38_8 = t_r23_c38_4 + p_24_37;
  assign t_r23_c38_9 = t_r23_c38_5 + t_r23_c38_6;
  assign t_r23_c38_10 = t_r23_c38_7 + t_r23_c38_8;
  assign t_r23_c38_11 = t_r23_c38_9 + t_r23_c38_10;
  assign t_r23_c38_12 = t_r23_c38_11 + p_24_39;
  assign out_23_38 = t_r23_c38_12 >> 4;

  assign t_r23_c39_0 = p_22_39 << 1;
  assign t_r23_c39_1 = p_23_38 << 1;
  assign t_r23_c39_2 = p_23_39 << 2;
  assign t_r23_c39_3 = p_23_40 << 1;
  assign t_r23_c39_4 = p_24_39 << 1;
  assign t_r23_c39_5 = t_r23_c39_0 + p_22_38;
  assign t_r23_c39_6 = t_r23_c39_1 + p_22_40;
  assign t_r23_c39_7 = t_r23_c39_2 + t_r23_c39_3;
  assign t_r23_c39_8 = t_r23_c39_4 + p_24_38;
  assign t_r23_c39_9 = t_r23_c39_5 + t_r23_c39_6;
  assign t_r23_c39_10 = t_r23_c39_7 + t_r23_c39_8;
  assign t_r23_c39_11 = t_r23_c39_9 + t_r23_c39_10;
  assign t_r23_c39_12 = t_r23_c39_11 + p_24_40;
  assign out_23_39 = t_r23_c39_12 >> 4;

  assign t_r23_c40_0 = p_22_40 << 1;
  assign t_r23_c40_1 = p_23_39 << 1;
  assign t_r23_c40_2 = p_23_40 << 2;
  assign t_r23_c40_3 = p_23_41 << 1;
  assign t_r23_c40_4 = p_24_40 << 1;
  assign t_r23_c40_5 = t_r23_c40_0 + p_22_39;
  assign t_r23_c40_6 = t_r23_c40_1 + p_22_41;
  assign t_r23_c40_7 = t_r23_c40_2 + t_r23_c40_3;
  assign t_r23_c40_8 = t_r23_c40_4 + p_24_39;
  assign t_r23_c40_9 = t_r23_c40_5 + t_r23_c40_6;
  assign t_r23_c40_10 = t_r23_c40_7 + t_r23_c40_8;
  assign t_r23_c40_11 = t_r23_c40_9 + t_r23_c40_10;
  assign t_r23_c40_12 = t_r23_c40_11 + p_24_41;
  assign out_23_40 = t_r23_c40_12 >> 4;

  assign t_r23_c41_0 = p_22_41 << 1;
  assign t_r23_c41_1 = p_23_40 << 1;
  assign t_r23_c41_2 = p_23_41 << 2;
  assign t_r23_c41_3 = p_23_42 << 1;
  assign t_r23_c41_4 = p_24_41 << 1;
  assign t_r23_c41_5 = t_r23_c41_0 + p_22_40;
  assign t_r23_c41_6 = t_r23_c41_1 + p_22_42;
  assign t_r23_c41_7 = t_r23_c41_2 + t_r23_c41_3;
  assign t_r23_c41_8 = t_r23_c41_4 + p_24_40;
  assign t_r23_c41_9 = t_r23_c41_5 + t_r23_c41_6;
  assign t_r23_c41_10 = t_r23_c41_7 + t_r23_c41_8;
  assign t_r23_c41_11 = t_r23_c41_9 + t_r23_c41_10;
  assign t_r23_c41_12 = t_r23_c41_11 + p_24_42;
  assign out_23_41 = t_r23_c41_12 >> 4;

  assign t_r23_c42_0 = p_22_42 << 1;
  assign t_r23_c42_1 = p_23_41 << 1;
  assign t_r23_c42_2 = p_23_42 << 2;
  assign t_r23_c42_3 = p_23_43 << 1;
  assign t_r23_c42_4 = p_24_42 << 1;
  assign t_r23_c42_5 = t_r23_c42_0 + p_22_41;
  assign t_r23_c42_6 = t_r23_c42_1 + p_22_43;
  assign t_r23_c42_7 = t_r23_c42_2 + t_r23_c42_3;
  assign t_r23_c42_8 = t_r23_c42_4 + p_24_41;
  assign t_r23_c42_9 = t_r23_c42_5 + t_r23_c42_6;
  assign t_r23_c42_10 = t_r23_c42_7 + t_r23_c42_8;
  assign t_r23_c42_11 = t_r23_c42_9 + t_r23_c42_10;
  assign t_r23_c42_12 = t_r23_c42_11 + p_24_43;
  assign out_23_42 = t_r23_c42_12 >> 4;

  assign t_r23_c43_0 = p_22_43 << 1;
  assign t_r23_c43_1 = p_23_42 << 1;
  assign t_r23_c43_2 = p_23_43 << 2;
  assign t_r23_c43_3 = p_23_44 << 1;
  assign t_r23_c43_4 = p_24_43 << 1;
  assign t_r23_c43_5 = t_r23_c43_0 + p_22_42;
  assign t_r23_c43_6 = t_r23_c43_1 + p_22_44;
  assign t_r23_c43_7 = t_r23_c43_2 + t_r23_c43_3;
  assign t_r23_c43_8 = t_r23_c43_4 + p_24_42;
  assign t_r23_c43_9 = t_r23_c43_5 + t_r23_c43_6;
  assign t_r23_c43_10 = t_r23_c43_7 + t_r23_c43_8;
  assign t_r23_c43_11 = t_r23_c43_9 + t_r23_c43_10;
  assign t_r23_c43_12 = t_r23_c43_11 + p_24_44;
  assign out_23_43 = t_r23_c43_12 >> 4;

  assign t_r23_c44_0 = p_22_44 << 1;
  assign t_r23_c44_1 = p_23_43 << 1;
  assign t_r23_c44_2 = p_23_44 << 2;
  assign t_r23_c44_3 = p_23_45 << 1;
  assign t_r23_c44_4 = p_24_44 << 1;
  assign t_r23_c44_5 = t_r23_c44_0 + p_22_43;
  assign t_r23_c44_6 = t_r23_c44_1 + p_22_45;
  assign t_r23_c44_7 = t_r23_c44_2 + t_r23_c44_3;
  assign t_r23_c44_8 = t_r23_c44_4 + p_24_43;
  assign t_r23_c44_9 = t_r23_c44_5 + t_r23_c44_6;
  assign t_r23_c44_10 = t_r23_c44_7 + t_r23_c44_8;
  assign t_r23_c44_11 = t_r23_c44_9 + t_r23_c44_10;
  assign t_r23_c44_12 = t_r23_c44_11 + p_24_45;
  assign out_23_44 = t_r23_c44_12 >> 4;

  assign t_r23_c45_0 = p_22_45 << 1;
  assign t_r23_c45_1 = p_23_44 << 1;
  assign t_r23_c45_2 = p_23_45 << 2;
  assign t_r23_c45_3 = p_23_46 << 1;
  assign t_r23_c45_4 = p_24_45 << 1;
  assign t_r23_c45_5 = t_r23_c45_0 + p_22_44;
  assign t_r23_c45_6 = t_r23_c45_1 + p_22_46;
  assign t_r23_c45_7 = t_r23_c45_2 + t_r23_c45_3;
  assign t_r23_c45_8 = t_r23_c45_4 + p_24_44;
  assign t_r23_c45_9 = t_r23_c45_5 + t_r23_c45_6;
  assign t_r23_c45_10 = t_r23_c45_7 + t_r23_c45_8;
  assign t_r23_c45_11 = t_r23_c45_9 + t_r23_c45_10;
  assign t_r23_c45_12 = t_r23_c45_11 + p_24_46;
  assign out_23_45 = t_r23_c45_12 >> 4;

  assign t_r23_c46_0 = p_22_46 << 1;
  assign t_r23_c46_1 = p_23_45 << 1;
  assign t_r23_c46_2 = p_23_46 << 2;
  assign t_r23_c46_3 = p_23_47 << 1;
  assign t_r23_c46_4 = p_24_46 << 1;
  assign t_r23_c46_5 = t_r23_c46_0 + p_22_45;
  assign t_r23_c46_6 = t_r23_c46_1 + p_22_47;
  assign t_r23_c46_7 = t_r23_c46_2 + t_r23_c46_3;
  assign t_r23_c46_8 = t_r23_c46_4 + p_24_45;
  assign t_r23_c46_9 = t_r23_c46_5 + t_r23_c46_6;
  assign t_r23_c46_10 = t_r23_c46_7 + t_r23_c46_8;
  assign t_r23_c46_11 = t_r23_c46_9 + t_r23_c46_10;
  assign t_r23_c46_12 = t_r23_c46_11 + p_24_47;
  assign out_23_46 = t_r23_c46_12 >> 4;

  assign t_r23_c47_0 = p_22_47 << 1;
  assign t_r23_c47_1 = p_23_46 << 1;
  assign t_r23_c47_2 = p_23_47 << 2;
  assign t_r23_c47_3 = p_23_48 << 1;
  assign t_r23_c47_4 = p_24_47 << 1;
  assign t_r23_c47_5 = t_r23_c47_0 + p_22_46;
  assign t_r23_c47_6 = t_r23_c47_1 + p_22_48;
  assign t_r23_c47_7 = t_r23_c47_2 + t_r23_c47_3;
  assign t_r23_c47_8 = t_r23_c47_4 + p_24_46;
  assign t_r23_c47_9 = t_r23_c47_5 + t_r23_c47_6;
  assign t_r23_c47_10 = t_r23_c47_7 + t_r23_c47_8;
  assign t_r23_c47_11 = t_r23_c47_9 + t_r23_c47_10;
  assign t_r23_c47_12 = t_r23_c47_11 + p_24_48;
  assign out_23_47 = t_r23_c47_12 >> 4;

  assign t_r23_c48_0 = p_22_48 << 1;
  assign t_r23_c48_1 = p_23_47 << 1;
  assign t_r23_c48_2 = p_23_48 << 2;
  assign t_r23_c48_3 = p_23_49 << 1;
  assign t_r23_c48_4 = p_24_48 << 1;
  assign t_r23_c48_5 = t_r23_c48_0 + p_22_47;
  assign t_r23_c48_6 = t_r23_c48_1 + p_22_49;
  assign t_r23_c48_7 = t_r23_c48_2 + t_r23_c48_3;
  assign t_r23_c48_8 = t_r23_c48_4 + p_24_47;
  assign t_r23_c48_9 = t_r23_c48_5 + t_r23_c48_6;
  assign t_r23_c48_10 = t_r23_c48_7 + t_r23_c48_8;
  assign t_r23_c48_11 = t_r23_c48_9 + t_r23_c48_10;
  assign t_r23_c48_12 = t_r23_c48_11 + p_24_49;
  assign out_23_48 = t_r23_c48_12 >> 4;

  assign t_r23_c49_0 = p_22_49 << 1;
  assign t_r23_c49_1 = p_23_48 << 1;
  assign t_r23_c49_2 = p_23_49 << 2;
  assign t_r23_c49_3 = p_23_50 << 1;
  assign t_r23_c49_4 = p_24_49 << 1;
  assign t_r23_c49_5 = t_r23_c49_0 + p_22_48;
  assign t_r23_c49_6 = t_r23_c49_1 + p_22_50;
  assign t_r23_c49_7 = t_r23_c49_2 + t_r23_c49_3;
  assign t_r23_c49_8 = t_r23_c49_4 + p_24_48;
  assign t_r23_c49_9 = t_r23_c49_5 + t_r23_c49_6;
  assign t_r23_c49_10 = t_r23_c49_7 + t_r23_c49_8;
  assign t_r23_c49_11 = t_r23_c49_9 + t_r23_c49_10;
  assign t_r23_c49_12 = t_r23_c49_11 + p_24_50;
  assign out_23_49 = t_r23_c49_12 >> 4;

  assign t_r23_c50_0 = p_22_50 << 1;
  assign t_r23_c50_1 = p_23_49 << 1;
  assign t_r23_c50_2 = p_23_50 << 2;
  assign t_r23_c50_3 = p_23_51 << 1;
  assign t_r23_c50_4 = p_24_50 << 1;
  assign t_r23_c50_5 = t_r23_c50_0 + p_22_49;
  assign t_r23_c50_6 = t_r23_c50_1 + p_22_51;
  assign t_r23_c50_7 = t_r23_c50_2 + t_r23_c50_3;
  assign t_r23_c50_8 = t_r23_c50_4 + p_24_49;
  assign t_r23_c50_9 = t_r23_c50_5 + t_r23_c50_6;
  assign t_r23_c50_10 = t_r23_c50_7 + t_r23_c50_8;
  assign t_r23_c50_11 = t_r23_c50_9 + t_r23_c50_10;
  assign t_r23_c50_12 = t_r23_c50_11 + p_24_51;
  assign out_23_50 = t_r23_c50_12 >> 4;

  assign t_r23_c51_0 = p_22_51 << 1;
  assign t_r23_c51_1 = p_23_50 << 1;
  assign t_r23_c51_2 = p_23_51 << 2;
  assign t_r23_c51_3 = p_23_52 << 1;
  assign t_r23_c51_4 = p_24_51 << 1;
  assign t_r23_c51_5 = t_r23_c51_0 + p_22_50;
  assign t_r23_c51_6 = t_r23_c51_1 + p_22_52;
  assign t_r23_c51_7 = t_r23_c51_2 + t_r23_c51_3;
  assign t_r23_c51_8 = t_r23_c51_4 + p_24_50;
  assign t_r23_c51_9 = t_r23_c51_5 + t_r23_c51_6;
  assign t_r23_c51_10 = t_r23_c51_7 + t_r23_c51_8;
  assign t_r23_c51_11 = t_r23_c51_9 + t_r23_c51_10;
  assign t_r23_c51_12 = t_r23_c51_11 + p_24_52;
  assign out_23_51 = t_r23_c51_12 >> 4;

  assign t_r23_c52_0 = p_22_52 << 1;
  assign t_r23_c52_1 = p_23_51 << 1;
  assign t_r23_c52_2 = p_23_52 << 2;
  assign t_r23_c52_3 = p_23_53 << 1;
  assign t_r23_c52_4 = p_24_52 << 1;
  assign t_r23_c52_5 = t_r23_c52_0 + p_22_51;
  assign t_r23_c52_6 = t_r23_c52_1 + p_22_53;
  assign t_r23_c52_7 = t_r23_c52_2 + t_r23_c52_3;
  assign t_r23_c52_8 = t_r23_c52_4 + p_24_51;
  assign t_r23_c52_9 = t_r23_c52_5 + t_r23_c52_6;
  assign t_r23_c52_10 = t_r23_c52_7 + t_r23_c52_8;
  assign t_r23_c52_11 = t_r23_c52_9 + t_r23_c52_10;
  assign t_r23_c52_12 = t_r23_c52_11 + p_24_53;
  assign out_23_52 = t_r23_c52_12 >> 4;

  assign t_r23_c53_0 = p_22_53 << 1;
  assign t_r23_c53_1 = p_23_52 << 1;
  assign t_r23_c53_2 = p_23_53 << 2;
  assign t_r23_c53_3 = p_23_54 << 1;
  assign t_r23_c53_4 = p_24_53 << 1;
  assign t_r23_c53_5 = t_r23_c53_0 + p_22_52;
  assign t_r23_c53_6 = t_r23_c53_1 + p_22_54;
  assign t_r23_c53_7 = t_r23_c53_2 + t_r23_c53_3;
  assign t_r23_c53_8 = t_r23_c53_4 + p_24_52;
  assign t_r23_c53_9 = t_r23_c53_5 + t_r23_c53_6;
  assign t_r23_c53_10 = t_r23_c53_7 + t_r23_c53_8;
  assign t_r23_c53_11 = t_r23_c53_9 + t_r23_c53_10;
  assign t_r23_c53_12 = t_r23_c53_11 + p_24_54;
  assign out_23_53 = t_r23_c53_12 >> 4;

  assign t_r23_c54_0 = p_22_54 << 1;
  assign t_r23_c54_1 = p_23_53 << 1;
  assign t_r23_c54_2 = p_23_54 << 2;
  assign t_r23_c54_3 = p_23_55 << 1;
  assign t_r23_c54_4 = p_24_54 << 1;
  assign t_r23_c54_5 = t_r23_c54_0 + p_22_53;
  assign t_r23_c54_6 = t_r23_c54_1 + p_22_55;
  assign t_r23_c54_7 = t_r23_c54_2 + t_r23_c54_3;
  assign t_r23_c54_8 = t_r23_c54_4 + p_24_53;
  assign t_r23_c54_9 = t_r23_c54_5 + t_r23_c54_6;
  assign t_r23_c54_10 = t_r23_c54_7 + t_r23_c54_8;
  assign t_r23_c54_11 = t_r23_c54_9 + t_r23_c54_10;
  assign t_r23_c54_12 = t_r23_c54_11 + p_24_55;
  assign out_23_54 = t_r23_c54_12 >> 4;

  assign t_r23_c55_0 = p_22_55 << 1;
  assign t_r23_c55_1 = p_23_54 << 1;
  assign t_r23_c55_2 = p_23_55 << 2;
  assign t_r23_c55_3 = p_23_56 << 1;
  assign t_r23_c55_4 = p_24_55 << 1;
  assign t_r23_c55_5 = t_r23_c55_0 + p_22_54;
  assign t_r23_c55_6 = t_r23_c55_1 + p_22_56;
  assign t_r23_c55_7 = t_r23_c55_2 + t_r23_c55_3;
  assign t_r23_c55_8 = t_r23_c55_4 + p_24_54;
  assign t_r23_c55_9 = t_r23_c55_5 + t_r23_c55_6;
  assign t_r23_c55_10 = t_r23_c55_7 + t_r23_c55_8;
  assign t_r23_c55_11 = t_r23_c55_9 + t_r23_c55_10;
  assign t_r23_c55_12 = t_r23_c55_11 + p_24_56;
  assign out_23_55 = t_r23_c55_12 >> 4;

  assign t_r23_c56_0 = p_22_56 << 1;
  assign t_r23_c56_1 = p_23_55 << 1;
  assign t_r23_c56_2 = p_23_56 << 2;
  assign t_r23_c56_3 = p_23_57 << 1;
  assign t_r23_c56_4 = p_24_56 << 1;
  assign t_r23_c56_5 = t_r23_c56_0 + p_22_55;
  assign t_r23_c56_6 = t_r23_c56_1 + p_22_57;
  assign t_r23_c56_7 = t_r23_c56_2 + t_r23_c56_3;
  assign t_r23_c56_8 = t_r23_c56_4 + p_24_55;
  assign t_r23_c56_9 = t_r23_c56_5 + t_r23_c56_6;
  assign t_r23_c56_10 = t_r23_c56_7 + t_r23_c56_8;
  assign t_r23_c56_11 = t_r23_c56_9 + t_r23_c56_10;
  assign t_r23_c56_12 = t_r23_c56_11 + p_24_57;
  assign out_23_56 = t_r23_c56_12 >> 4;

  assign t_r23_c57_0 = p_22_57 << 1;
  assign t_r23_c57_1 = p_23_56 << 1;
  assign t_r23_c57_2 = p_23_57 << 2;
  assign t_r23_c57_3 = p_23_58 << 1;
  assign t_r23_c57_4 = p_24_57 << 1;
  assign t_r23_c57_5 = t_r23_c57_0 + p_22_56;
  assign t_r23_c57_6 = t_r23_c57_1 + p_22_58;
  assign t_r23_c57_7 = t_r23_c57_2 + t_r23_c57_3;
  assign t_r23_c57_8 = t_r23_c57_4 + p_24_56;
  assign t_r23_c57_9 = t_r23_c57_5 + t_r23_c57_6;
  assign t_r23_c57_10 = t_r23_c57_7 + t_r23_c57_8;
  assign t_r23_c57_11 = t_r23_c57_9 + t_r23_c57_10;
  assign t_r23_c57_12 = t_r23_c57_11 + p_24_58;
  assign out_23_57 = t_r23_c57_12 >> 4;

  assign t_r23_c58_0 = p_22_58 << 1;
  assign t_r23_c58_1 = p_23_57 << 1;
  assign t_r23_c58_2 = p_23_58 << 2;
  assign t_r23_c58_3 = p_23_59 << 1;
  assign t_r23_c58_4 = p_24_58 << 1;
  assign t_r23_c58_5 = t_r23_c58_0 + p_22_57;
  assign t_r23_c58_6 = t_r23_c58_1 + p_22_59;
  assign t_r23_c58_7 = t_r23_c58_2 + t_r23_c58_3;
  assign t_r23_c58_8 = t_r23_c58_4 + p_24_57;
  assign t_r23_c58_9 = t_r23_c58_5 + t_r23_c58_6;
  assign t_r23_c58_10 = t_r23_c58_7 + t_r23_c58_8;
  assign t_r23_c58_11 = t_r23_c58_9 + t_r23_c58_10;
  assign t_r23_c58_12 = t_r23_c58_11 + p_24_59;
  assign out_23_58 = t_r23_c58_12 >> 4;

  assign t_r23_c59_0 = p_22_59 << 1;
  assign t_r23_c59_1 = p_23_58 << 1;
  assign t_r23_c59_2 = p_23_59 << 2;
  assign t_r23_c59_3 = p_23_60 << 1;
  assign t_r23_c59_4 = p_24_59 << 1;
  assign t_r23_c59_5 = t_r23_c59_0 + p_22_58;
  assign t_r23_c59_6 = t_r23_c59_1 + p_22_60;
  assign t_r23_c59_7 = t_r23_c59_2 + t_r23_c59_3;
  assign t_r23_c59_8 = t_r23_c59_4 + p_24_58;
  assign t_r23_c59_9 = t_r23_c59_5 + t_r23_c59_6;
  assign t_r23_c59_10 = t_r23_c59_7 + t_r23_c59_8;
  assign t_r23_c59_11 = t_r23_c59_9 + t_r23_c59_10;
  assign t_r23_c59_12 = t_r23_c59_11 + p_24_60;
  assign out_23_59 = t_r23_c59_12 >> 4;

  assign t_r23_c60_0 = p_22_60 << 1;
  assign t_r23_c60_1 = p_23_59 << 1;
  assign t_r23_c60_2 = p_23_60 << 2;
  assign t_r23_c60_3 = p_23_61 << 1;
  assign t_r23_c60_4 = p_24_60 << 1;
  assign t_r23_c60_5 = t_r23_c60_0 + p_22_59;
  assign t_r23_c60_6 = t_r23_c60_1 + p_22_61;
  assign t_r23_c60_7 = t_r23_c60_2 + t_r23_c60_3;
  assign t_r23_c60_8 = t_r23_c60_4 + p_24_59;
  assign t_r23_c60_9 = t_r23_c60_5 + t_r23_c60_6;
  assign t_r23_c60_10 = t_r23_c60_7 + t_r23_c60_8;
  assign t_r23_c60_11 = t_r23_c60_9 + t_r23_c60_10;
  assign t_r23_c60_12 = t_r23_c60_11 + p_24_61;
  assign out_23_60 = t_r23_c60_12 >> 4;

  assign t_r23_c61_0 = p_22_61 << 1;
  assign t_r23_c61_1 = p_23_60 << 1;
  assign t_r23_c61_2 = p_23_61 << 2;
  assign t_r23_c61_3 = p_23_62 << 1;
  assign t_r23_c61_4 = p_24_61 << 1;
  assign t_r23_c61_5 = t_r23_c61_0 + p_22_60;
  assign t_r23_c61_6 = t_r23_c61_1 + p_22_62;
  assign t_r23_c61_7 = t_r23_c61_2 + t_r23_c61_3;
  assign t_r23_c61_8 = t_r23_c61_4 + p_24_60;
  assign t_r23_c61_9 = t_r23_c61_5 + t_r23_c61_6;
  assign t_r23_c61_10 = t_r23_c61_7 + t_r23_c61_8;
  assign t_r23_c61_11 = t_r23_c61_9 + t_r23_c61_10;
  assign t_r23_c61_12 = t_r23_c61_11 + p_24_62;
  assign out_23_61 = t_r23_c61_12 >> 4;

  assign t_r23_c62_0 = p_22_62 << 1;
  assign t_r23_c62_1 = p_23_61 << 1;
  assign t_r23_c62_2 = p_23_62 << 2;
  assign t_r23_c62_3 = p_23_63 << 1;
  assign t_r23_c62_4 = p_24_62 << 1;
  assign t_r23_c62_5 = t_r23_c62_0 + p_22_61;
  assign t_r23_c62_6 = t_r23_c62_1 + p_22_63;
  assign t_r23_c62_7 = t_r23_c62_2 + t_r23_c62_3;
  assign t_r23_c62_8 = t_r23_c62_4 + p_24_61;
  assign t_r23_c62_9 = t_r23_c62_5 + t_r23_c62_6;
  assign t_r23_c62_10 = t_r23_c62_7 + t_r23_c62_8;
  assign t_r23_c62_11 = t_r23_c62_9 + t_r23_c62_10;
  assign t_r23_c62_12 = t_r23_c62_11 + p_24_63;
  assign out_23_62 = t_r23_c62_12 >> 4;

  assign t_r23_c63_0 = p_22_63 << 1;
  assign t_r23_c63_1 = p_23_62 << 1;
  assign t_r23_c63_2 = p_23_63 << 2;
  assign t_r23_c63_3 = p_23_64 << 1;
  assign t_r23_c63_4 = p_24_63 << 1;
  assign t_r23_c63_5 = t_r23_c63_0 + p_22_62;
  assign t_r23_c63_6 = t_r23_c63_1 + p_22_64;
  assign t_r23_c63_7 = t_r23_c63_2 + t_r23_c63_3;
  assign t_r23_c63_8 = t_r23_c63_4 + p_24_62;
  assign t_r23_c63_9 = t_r23_c63_5 + t_r23_c63_6;
  assign t_r23_c63_10 = t_r23_c63_7 + t_r23_c63_8;
  assign t_r23_c63_11 = t_r23_c63_9 + t_r23_c63_10;
  assign t_r23_c63_12 = t_r23_c63_11 + p_24_64;
  assign out_23_63 = t_r23_c63_12 >> 4;

  assign t_r23_c64_0 = p_22_64 << 1;
  assign t_r23_c64_1 = p_23_63 << 1;
  assign t_r23_c64_2 = p_23_64 << 2;
  assign t_r23_c64_3 = p_23_65 << 1;
  assign t_r23_c64_4 = p_24_64 << 1;
  assign t_r23_c64_5 = t_r23_c64_0 + p_22_63;
  assign t_r23_c64_6 = t_r23_c64_1 + p_22_65;
  assign t_r23_c64_7 = t_r23_c64_2 + t_r23_c64_3;
  assign t_r23_c64_8 = t_r23_c64_4 + p_24_63;
  assign t_r23_c64_9 = t_r23_c64_5 + t_r23_c64_6;
  assign t_r23_c64_10 = t_r23_c64_7 + t_r23_c64_8;
  assign t_r23_c64_11 = t_r23_c64_9 + t_r23_c64_10;
  assign t_r23_c64_12 = t_r23_c64_11 + p_24_65;
  assign out_23_64 = t_r23_c64_12 >> 4;

  assign t_r24_c1_0 = p_23_1 << 1;
  assign t_r24_c1_1 = p_24_0 << 1;
  assign t_r24_c1_2 = p_24_1 << 2;
  assign t_r24_c1_3 = p_24_2 << 1;
  assign t_r24_c1_4 = p_25_1 << 1;
  assign t_r24_c1_5 = t_r24_c1_0 + p_23_0;
  assign t_r24_c1_6 = t_r24_c1_1 + p_23_2;
  assign t_r24_c1_7 = t_r24_c1_2 + t_r24_c1_3;
  assign t_r24_c1_8 = t_r24_c1_4 + p_25_0;
  assign t_r24_c1_9 = t_r24_c1_5 + t_r24_c1_6;
  assign t_r24_c1_10 = t_r24_c1_7 + t_r24_c1_8;
  assign t_r24_c1_11 = t_r24_c1_9 + t_r24_c1_10;
  assign t_r24_c1_12 = t_r24_c1_11 + p_25_2;
  assign out_24_1 = t_r24_c1_12 >> 4;

  assign t_r24_c2_0 = p_23_2 << 1;
  assign t_r24_c2_1 = p_24_1 << 1;
  assign t_r24_c2_2 = p_24_2 << 2;
  assign t_r24_c2_3 = p_24_3 << 1;
  assign t_r24_c2_4 = p_25_2 << 1;
  assign t_r24_c2_5 = t_r24_c2_0 + p_23_1;
  assign t_r24_c2_6 = t_r24_c2_1 + p_23_3;
  assign t_r24_c2_7 = t_r24_c2_2 + t_r24_c2_3;
  assign t_r24_c2_8 = t_r24_c2_4 + p_25_1;
  assign t_r24_c2_9 = t_r24_c2_5 + t_r24_c2_6;
  assign t_r24_c2_10 = t_r24_c2_7 + t_r24_c2_8;
  assign t_r24_c2_11 = t_r24_c2_9 + t_r24_c2_10;
  assign t_r24_c2_12 = t_r24_c2_11 + p_25_3;
  assign out_24_2 = t_r24_c2_12 >> 4;

  assign t_r24_c3_0 = p_23_3 << 1;
  assign t_r24_c3_1 = p_24_2 << 1;
  assign t_r24_c3_2 = p_24_3 << 2;
  assign t_r24_c3_3 = p_24_4 << 1;
  assign t_r24_c3_4 = p_25_3 << 1;
  assign t_r24_c3_5 = t_r24_c3_0 + p_23_2;
  assign t_r24_c3_6 = t_r24_c3_1 + p_23_4;
  assign t_r24_c3_7 = t_r24_c3_2 + t_r24_c3_3;
  assign t_r24_c3_8 = t_r24_c3_4 + p_25_2;
  assign t_r24_c3_9 = t_r24_c3_5 + t_r24_c3_6;
  assign t_r24_c3_10 = t_r24_c3_7 + t_r24_c3_8;
  assign t_r24_c3_11 = t_r24_c3_9 + t_r24_c3_10;
  assign t_r24_c3_12 = t_r24_c3_11 + p_25_4;
  assign out_24_3 = t_r24_c3_12 >> 4;

  assign t_r24_c4_0 = p_23_4 << 1;
  assign t_r24_c4_1 = p_24_3 << 1;
  assign t_r24_c4_2 = p_24_4 << 2;
  assign t_r24_c4_3 = p_24_5 << 1;
  assign t_r24_c4_4 = p_25_4 << 1;
  assign t_r24_c4_5 = t_r24_c4_0 + p_23_3;
  assign t_r24_c4_6 = t_r24_c4_1 + p_23_5;
  assign t_r24_c4_7 = t_r24_c4_2 + t_r24_c4_3;
  assign t_r24_c4_8 = t_r24_c4_4 + p_25_3;
  assign t_r24_c4_9 = t_r24_c4_5 + t_r24_c4_6;
  assign t_r24_c4_10 = t_r24_c4_7 + t_r24_c4_8;
  assign t_r24_c4_11 = t_r24_c4_9 + t_r24_c4_10;
  assign t_r24_c4_12 = t_r24_c4_11 + p_25_5;
  assign out_24_4 = t_r24_c4_12 >> 4;

  assign t_r24_c5_0 = p_23_5 << 1;
  assign t_r24_c5_1 = p_24_4 << 1;
  assign t_r24_c5_2 = p_24_5 << 2;
  assign t_r24_c5_3 = p_24_6 << 1;
  assign t_r24_c5_4 = p_25_5 << 1;
  assign t_r24_c5_5 = t_r24_c5_0 + p_23_4;
  assign t_r24_c5_6 = t_r24_c5_1 + p_23_6;
  assign t_r24_c5_7 = t_r24_c5_2 + t_r24_c5_3;
  assign t_r24_c5_8 = t_r24_c5_4 + p_25_4;
  assign t_r24_c5_9 = t_r24_c5_5 + t_r24_c5_6;
  assign t_r24_c5_10 = t_r24_c5_7 + t_r24_c5_8;
  assign t_r24_c5_11 = t_r24_c5_9 + t_r24_c5_10;
  assign t_r24_c5_12 = t_r24_c5_11 + p_25_6;
  assign out_24_5 = t_r24_c5_12 >> 4;

  assign t_r24_c6_0 = p_23_6 << 1;
  assign t_r24_c6_1 = p_24_5 << 1;
  assign t_r24_c6_2 = p_24_6 << 2;
  assign t_r24_c6_3 = p_24_7 << 1;
  assign t_r24_c6_4 = p_25_6 << 1;
  assign t_r24_c6_5 = t_r24_c6_0 + p_23_5;
  assign t_r24_c6_6 = t_r24_c6_1 + p_23_7;
  assign t_r24_c6_7 = t_r24_c6_2 + t_r24_c6_3;
  assign t_r24_c6_8 = t_r24_c6_4 + p_25_5;
  assign t_r24_c6_9 = t_r24_c6_5 + t_r24_c6_6;
  assign t_r24_c6_10 = t_r24_c6_7 + t_r24_c6_8;
  assign t_r24_c6_11 = t_r24_c6_9 + t_r24_c6_10;
  assign t_r24_c6_12 = t_r24_c6_11 + p_25_7;
  assign out_24_6 = t_r24_c6_12 >> 4;

  assign t_r24_c7_0 = p_23_7 << 1;
  assign t_r24_c7_1 = p_24_6 << 1;
  assign t_r24_c7_2 = p_24_7 << 2;
  assign t_r24_c7_3 = p_24_8 << 1;
  assign t_r24_c7_4 = p_25_7 << 1;
  assign t_r24_c7_5 = t_r24_c7_0 + p_23_6;
  assign t_r24_c7_6 = t_r24_c7_1 + p_23_8;
  assign t_r24_c7_7 = t_r24_c7_2 + t_r24_c7_3;
  assign t_r24_c7_8 = t_r24_c7_4 + p_25_6;
  assign t_r24_c7_9 = t_r24_c7_5 + t_r24_c7_6;
  assign t_r24_c7_10 = t_r24_c7_7 + t_r24_c7_8;
  assign t_r24_c7_11 = t_r24_c7_9 + t_r24_c7_10;
  assign t_r24_c7_12 = t_r24_c7_11 + p_25_8;
  assign out_24_7 = t_r24_c7_12 >> 4;

  assign t_r24_c8_0 = p_23_8 << 1;
  assign t_r24_c8_1 = p_24_7 << 1;
  assign t_r24_c8_2 = p_24_8 << 2;
  assign t_r24_c8_3 = p_24_9 << 1;
  assign t_r24_c8_4 = p_25_8 << 1;
  assign t_r24_c8_5 = t_r24_c8_0 + p_23_7;
  assign t_r24_c8_6 = t_r24_c8_1 + p_23_9;
  assign t_r24_c8_7 = t_r24_c8_2 + t_r24_c8_3;
  assign t_r24_c8_8 = t_r24_c8_4 + p_25_7;
  assign t_r24_c8_9 = t_r24_c8_5 + t_r24_c8_6;
  assign t_r24_c8_10 = t_r24_c8_7 + t_r24_c8_8;
  assign t_r24_c8_11 = t_r24_c8_9 + t_r24_c8_10;
  assign t_r24_c8_12 = t_r24_c8_11 + p_25_9;
  assign out_24_8 = t_r24_c8_12 >> 4;

  assign t_r24_c9_0 = p_23_9 << 1;
  assign t_r24_c9_1 = p_24_8 << 1;
  assign t_r24_c9_2 = p_24_9 << 2;
  assign t_r24_c9_3 = p_24_10 << 1;
  assign t_r24_c9_4 = p_25_9 << 1;
  assign t_r24_c9_5 = t_r24_c9_0 + p_23_8;
  assign t_r24_c9_6 = t_r24_c9_1 + p_23_10;
  assign t_r24_c9_7 = t_r24_c9_2 + t_r24_c9_3;
  assign t_r24_c9_8 = t_r24_c9_4 + p_25_8;
  assign t_r24_c9_9 = t_r24_c9_5 + t_r24_c9_6;
  assign t_r24_c9_10 = t_r24_c9_7 + t_r24_c9_8;
  assign t_r24_c9_11 = t_r24_c9_9 + t_r24_c9_10;
  assign t_r24_c9_12 = t_r24_c9_11 + p_25_10;
  assign out_24_9 = t_r24_c9_12 >> 4;

  assign t_r24_c10_0 = p_23_10 << 1;
  assign t_r24_c10_1 = p_24_9 << 1;
  assign t_r24_c10_2 = p_24_10 << 2;
  assign t_r24_c10_3 = p_24_11 << 1;
  assign t_r24_c10_4 = p_25_10 << 1;
  assign t_r24_c10_5 = t_r24_c10_0 + p_23_9;
  assign t_r24_c10_6 = t_r24_c10_1 + p_23_11;
  assign t_r24_c10_7 = t_r24_c10_2 + t_r24_c10_3;
  assign t_r24_c10_8 = t_r24_c10_4 + p_25_9;
  assign t_r24_c10_9 = t_r24_c10_5 + t_r24_c10_6;
  assign t_r24_c10_10 = t_r24_c10_7 + t_r24_c10_8;
  assign t_r24_c10_11 = t_r24_c10_9 + t_r24_c10_10;
  assign t_r24_c10_12 = t_r24_c10_11 + p_25_11;
  assign out_24_10 = t_r24_c10_12 >> 4;

  assign t_r24_c11_0 = p_23_11 << 1;
  assign t_r24_c11_1 = p_24_10 << 1;
  assign t_r24_c11_2 = p_24_11 << 2;
  assign t_r24_c11_3 = p_24_12 << 1;
  assign t_r24_c11_4 = p_25_11 << 1;
  assign t_r24_c11_5 = t_r24_c11_0 + p_23_10;
  assign t_r24_c11_6 = t_r24_c11_1 + p_23_12;
  assign t_r24_c11_7 = t_r24_c11_2 + t_r24_c11_3;
  assign t_r24_c11_8 = t_r24_c11_4 + p_25_10;
  assign t_r24_c11_9 = t_r24_c11_5 + t_r24_c11_6;
  assign t_r24_c11_10 = t_r24_c11_7 + t_r24_c11_8;
  assign t_r24_c11_11 = t_r24_c11_9 + t_r24_c11_10;
  assign t_r24_c11_12 = t_r24_c11_11 + p_25_12;
  assign out_24_11 = t_r24_c11_12 >> 4;

  assign t_r24_c12_0 = p_23_12 << 1;
  assign t_r24_c12_1 = p_24_11 << 1;
  assign t_r24_c12_2 = p_24_12 << 2;
  assign t_r24_c12_3 = p_24_13 << 1;
  assign t_r24_c12_4 = p_25_12 << 1;
  assign t_r24_c12_5 = t_r24_c12_0 + p_23_11;
  assign t_r24_c12_6 = t_r24_c12_1 + p_23_13;
  assign t_r24_c12_7 = t_r24_c12_2 + t_r24_c12_3;
  assign t_r24_c12_8 = t_r24_c12_4 + p_25_11;
  assign t_r24_c12_9 = t_r24_c12_5 + t_r24_c12_6;
  assign t_r24_c12_10 = t_r24_c12_7 + t_r24_c12_8;
  assign t_r24_c12_11 = t_r24_c12_9 + t_r24_c12_10;
  assign t_r24_c12_12 = t_r24_c12_11 + p_25_13;
  assign out_24_12 = t_r24_c12_12 >> 4;

  assign t_r24_c13_0 = p_23_13 << 1;
  assign t_r24_c13_1 = p_24_12 << 1;
  assign t_r24_c13_2 = p_24_13 << 2;
  assign t_r24_c13_3 = p_24_14 << 1;
  assign t_r24_c13_4 = p_25_13 << 1;
  assign t_r24_c13_5 = t_r24_c13_0 + p_23_12;
  assign t_r24_c13_6 = t_r24_c13_1 + p_23_14;
  assign t_r24_c13_7 = t_r24_c13_2 + t_r24_c13_3;
  assign t_r24_c13_8 = t_r24_c13_4 + p_25_12;
  assign t_r24_c13_9 = t_r24_c13_5 + t_r24_c13_6;
  assign t_r24_c13_10 = t_r24_c13_7 + t_r24_c13_8;
  assign t_r24_c13_11 = t_r24_c13_9 + t_r24_c13_10;
  assign t_r24_c13_12 = t_r24_c13_11 + p_25_14;
  assign out_24_13 = t_r24_c13_12 >> 4;

  assign t_r24_c14_0 = p_23_14 << 1;
  assign t_r24_c14_1 = p_24_13 << 1;
  assign t_r24_c14_2 = p_24_14 << 2;
  assign t_r24_c14_3 = p_24_15 << 1;
  assign t_r24_c14_4 = p_25_14 << 1;
  assign t_r24_c14_5 = t_r24_c14_0 + p_23_13;
  assign t_r24_c14_6 = t_r24_c14_1 + p_23_15;
  assign t_r24_c14_7 = t_r24_c14_2 + t_r24_c14_3;
  assign t_r24_c14_8 = t_r24_c14_4 + p_25_13;
  assign t_r24_c14_9 = t_r24_c14_5 + t_r24_c14_6;
  assign t_r24_c14_10 = t_r24_c14_7 + t_r24_c14_8;
  assign t_r24_c14_11 = t_r24_c14_9 + t_r24_c14_10;
  assign t_r24_c14_12 = t_r24_c14_11 + p_25_15;
  assign out_24_14 = t_r24_c14_12 >> 4;

  assign t_r24_c15_0 = p_23_15 << 1;
  assign t_r24_c15_1 = p_24_14 << 1;
  assign t_r24_c15_2 = p_24_15 << 2;
  assign t_r24_c15_3 = p_24_16 << 1;
  assign t_r24_c15_4 = p_25_15 << 1;
  assign t_r24_c15_5 = t_r24_c15_0 + p_23_14;
  assign t_r24_c15_6 = t_r24_c15_1 + p_23_16;
  assign t_r24_c15_7 = t_r24_c15_2 + t_r24_c15_3;
  assign t_r24_c15_8 = t_r24_c15_4 + p_25_14;
  assign t_r24_c15_9 = t_r24_c15_5 + t_r24_c15_6;
  assign t_r24_c15_10 = t_r24_c15_7 + t_r24_c15_8;
  assign t_r24_c15_11 = t_r24_c15_9 + t_r24_c15_10;
  assign t_r24_c15_12 = t_r24_c15_11 + p_25_16;
  assign out_24_15 = t_r24_c15_12 >> 4;

  assign t_r24_c16_0 = p_23_16 << 1;
  assign t_r24_c16_1 = p_24_15 << 1;
  assign t_r24_c16_2 = p_24_16 << 2;
  assign t_r24_c16_3 = p_24_17 << 1;
  assign t_r24_c16_4 = p_25_16 << 1;
  assign t_r24_c16_5 = t_r24_c16_0 + p_23_15;
  assign t_r24_c16_6 = t_r24_c16_1 + p_23_17;
  assign t_r24_c16_7 = t_r24_c16_2 + t_r24_c16_3;
  assign t_r24_c16_8 = t_r24_c16_4 + p_25_15;
  assign t_r24_c16_9 = t_r24_c16_5 + t_r24_c16_6;
  assign t_r24_c16_10 = t_r24_c16_7 + t_r24_c16_8;
  assign t_r24_c16_11 = t_r24_c16_9 + t_r24_c16_10;
  assign t_r24_c16_12 = t_r24_c16_11 + p_25_17;
  assign out_24_16 = t_r24_c16_12 >> 4;

  assign t_r24_c17_0 = p_23_17 << 1;
  assign t_r24_c17_1 = p_24_16 << 1;
  assign t_r24_c17_2 = p_24_17 << 2;
  assign t_r24_c17_3 = p_24_18 << 1;
  assign t_r24_c17_4 = p_25_17 << 1;
  assign t_r24_c17_5 = t_r24_c17_0 + p_23_16;
  assign t_r24_c17_6 = t_r24_c17_1 + p_23_18;
  assign t_r24_c17_7 = t_r24_c17_2 + t_r24_c17_3;
  assign t_r24_c17_8 = t_r24_c17_4 + p_25_16;
  assign t_r24_c17_9 = t_r24_c17_5 + t_r24_c17_6;
  assign t_r24_c17_10 = t_r24_c17_7 + t_r24_c17_8;
  assign t_r24_c17_11 = t_r24_c17_9 + t_r24_c17_10;
  assign t_r24_c17_12 = t_r24_c17_11 + p_25_18;
  assign out_24_17 = t_r24_c17_12 >> 4;

  assign t_r24_c18_0 = p_23_18 << 1;
  assign t_r24_c18_1 = p_24_17 << 1;
  assign t_r24_c18_2 = p_24_18 << 2;
  assign t_r24_c18_3 = p_24_19 << 1;
  assign t_r24_c18_4 = p_25_18 << 1;
  assign t_r24_c18_5 = t_r24_c18_0 + p_23_17;
  assign t_r24_c18_6 = t_r24_c18_1 + p_23_19;
  assign t_r24_c18_7 = t_r24_c18_2 + t_r24_c18_3;
  assign t_r24_c18_8 = t_r24_c18_4 + p_25_17;
  assign t_r24_c18_9 = t_r24_c18_5 + t_r24_c18_6;
  assign t_r24_c18_10 = t_r24_c18_7 + t_r24_c18_8;
  assign t_r24_c18_11 = t_r24_c18_9 + t_r24_c18_10;
  assign t_r24_c18_12 = t_r24_c18_11 + p_25_19;
  assign out_24_18 = t_r24_c18_12 >> 4;

  assign t_r24_c19_0 = p_23_19 << 1;
  assign t_r24_c19_1 = p_24_18 << 1;
  assign t_r24_c19_2 = p_24_19 << 2;
  assign t_r24_c19_3 = p_24_20 << 1;
  assign t_r24_c19_4 = p_25_19 << 1;
  assign t_r24_c19_5 = t_r24_c19_0 + p_23_18;
  assign t_r24_c19_6 = t_r24_c19_1 + p_23_20;
  assign t_r24_c19_7 = t_r24_c19_2 + t_r24_c19_3;
  assign t_r24_c19_8 = t_r24_c19_4 + p_25_18;
  assign t_r24_c19_9 = t_r24_c19_5 + t_r24_c19_6;
  assign t_r24_c19_10 = t_r24_c19_7 + t_r24_c19_8;
  assign t_r24_c19_11 = t_r24_c19_9 + t_r24_c19_10;
  assign t_r24_c19_12 = t_r24_c19_11 + p_25_20;
  assign out_24_19 = t_r24_c19_12 >> 4;

  assign t_r24_c20_0 = p_23_20 << 1;
  assign t_r24_c20_1 = p_24_19 << 1;
  assign t_r24_c20_2 = p_24_20 << 2;
  assign t_r24_c20_3 = p_24_21 << 1;
  assign t_r24_c20_4 = p_25_20 << 1;
  assign t_r24_c20_5 = t_r24_c20_0 + p_23_19;
  assign t_r24_c20_6 = t_r24_c20_1 + p_23_21;
  assign t_r24_c20_7 = t_r24_c20_2 + t_r24_c20_3;
  assign t_r24_c20_8 = t_r24_c20_4 + p_25_19;
  assign t_r24_c20_9 = t_r24_c20_5 + t_r24_c20_6;
  assign t_r24_c20_10 = t_r24_c20_7 + t_r24_c20_8;
  assign t_r24_c20_11 = t_r24_c20_9 + t_r24_c20_10;
  assign t_r24_c20_12 = t_r24_c20_11 + p_25_21;
  assign out_24_20 = t_r24_c20_12 >> 4;

  assign t_r24_c21_0 = p_23_21 << 1;
  assign t_r24_c21_1 = p_24_20 << 1;
  assign t_r24_c21_2 = p_24_21 << 2;
  assign t_r24_c21_3 = p_24_22 << 1;
  assign t_r24_c21_4 = p_25_21 << 1;
  assign t_r24_c21_5 = t_r24_c21_0 + p_23_20;
  assign t_r24_c21_6 = t_r24_c21_1 + p_23_22;
  assign t_r24_c21_7 = t_r24_c21_2 + t_r24_c21_3;
  assign t_r24_c21_8 = t_r24_c21_4 + p_25_20;
  assign t_r24_c21_9 = t_r24_c21_5 + t_r24_c21_6;
  assign t_r24_c21_10 = t_r24_c21_7 + t_r24_c21_8;
  assign t_r24_c21_11 = t_r24_c21_9 + t_r24_c21_10;
  assign t_r24_c21_12 = t_r24_c21_11 + p_25_22;
  assign out_24_21 = t_r24_c21_12 >> 4;

  assign t_r24_c22_0 = p_23_22 << 1;
  assign t_r24_c22_1 = p_24_21 << 1;
  assign t_r24_c22_2 = p_24_22 << 2;
  assign t_r24_c22_3 = p_24_23 << 1;
  assign t_r24_c22_4 = p_25_22 << 1;
  assign t_r24_c22_5 = t_r24_c22_0 + p_23_21;
  assign t_r24_c22_6 = t_r24_c22_1 + p_23_23;
  assign t_r24_c22_7 = t_r24_c22_2 + t_r24_c22_3;
  assign t_r24_c22_8 = t_r24_c22_4 + p_25_21;
  assign t_r24_c22_9 = t_r24_c22_5 + t_r24_c22_6;
  assign t_r24_c22_10 = t_r24_c22_7 + t_r24_c22_8;
  assign t_r24_c22_11 = t_r24_c22_9 + t_r24_c22_10;
  assign t_r24_c22_12 = t_r24_c22_11 + p_25_23;
  assign out_24_22 = t_r24_c22_12 >> 4;

  assign t_r24_c23_0 = p_23_23 << 1;
  assign t_r24_c23_1 = p_24_22 << 1;
  assign t_r24_c23_2 = p_24_23 << 2;
  assign t_r24_c23_3 = p_24_24 << 1;
  assign t_r24_c23_4 = p_25_23 << 1;
  assign t_r24_c23_5 = t_r24_c23_0 + p_23_22;
  assign t_r24_c23_6 = t_r24_c23_1 + p_23_24;
  assign t_r24_c23_7 = t_r24_c23_2 + t_r24_c23_3;
  assign t_r24_c23_8 = t_r24_c23_4 + p_25_22;
  assign t_r24_c23_9 = t_r24_c23_5 + t_r24_c23_6;
  assign t_r24_c23_10 = t_r24_c23_7 + t_r24_c23_8;
  assign t_r24_c23_11 = t_r24_c23_9 + t_r24_c23_10;
  assign t_r24_c23_12 = t_r24_c23_11 + p_25_24;
  assign out_24_23 = t_r24_c23_12 >> 4;

  assign t_r24_c24_0 = p_23_24 << 1;
  assign t_r24_c24_1 = p_24_23 << 1;
  assign t_r24_c24_2 = p_24_24 << 2;
  assign t_r24_c24_3 = p_24_25 << 1;
  assign t_r24_c24_4 = p_25_24 << 1;
  assign t_r24_c24_5 = t_r24_c24_0 + p_23_23;
  assign t_r24_c24_6 = t_r24_c24_1 + p_23_25;
  assign t_r24_c24_7 = t_r24_c24_2 + t_r24_c24_3;
  assign t_r24_c24_8 = t_r24_c24_4 + p_25_23;
  assign t_r24_c24_9 = t_r24_c24_5 + t_r24_c24_6;
  assign t_r24_c24_10 = t_r24_c24_7 + t_r24_c24_8;
  assign t_r24_c24_11 = t_r24_c24_9 + t_r24_c24_10;
  assign t_r24_c24_12 = t_r24_c24_11 + p_25_25;
  assign out_24_24 = t_r24_c24_12 >> 4;

  assign t_r24_c25_0 = p_23_25 << 1;
  assign t_r24_c25_1 = p_24_24 << 1;
  assign t_r24_c25_2 = p_24_25 << 2;
  assign t_r24_c25_3 = p_24_26 << 1;
  assign t_r24_c25_4 = p_25_25 << 1;
  assign t_r24_c25_5 = t_r24_c25_0 + p_23_24;
  assign t_r24_c25_6 = t_r24_c25_1 + p_23_26;
  assign t_r24_c25_7 = t_r24_c25_2 + t_r24_c25_3;
  assign t_r24_c25_8 = t_r24_c25_4 + p_25_24;
  assign t_r24_c25_9 = t_r24_c25_5 + t_r24_c25_6;
  assign t_r24_c25_10 = t_r24_c25_7 + t_r24_c25_8;
  assign t_r24_c25_11 = t_r24_c25_9 + t_r24_c25_10;
  assign t_r24_c25_12 = t_r24_c25_11 + p_25_26;
  assign out_24_25 = t_r24_c25_12 >> 4;

  assign t_r24_c26_0 = p_23_26 << 1;
  assign t_r24_c26_1 = p_24_25 << 1;
  assign t_r24_c26_2 = p_24_26 << 2;
  assign t_r24_c26_3 = p_24_27 << 1;
  assign t_r24_c26_4 = p_25_26 << 1;
  assign t_r24_c26_5 = t_r24_c26_0 + p_23_25;
  assign t_r24_c26_6 = t_r24_c26_1 + p_23_27;
  assign t_r24_c26_7 = t_r24_c26_2 + t_r24_c26_3;
  assign t_r24_c26_8 = t_r24_c26_4 + p_25_25;
  assign t_r24_c26_9 = t_r24_c26_5 + t_r24_c26_6;
  assign t_r24_c26_10 = t_r24_c26_7 + t_r24_c26_8;
  assign t_r24_c26_11 = t_r24_c26_9 + t_r24_c26_10;
  assign t_r24_c26_12 = t_r24_c26_11 + p_25_27;
  assign out_24_26 = t_r24_c26_12 >> 4;

  assign t_r24_c27_0 = p_23_27 << 1;
  assign t_r24_c27_1 = p_24_26 << 1;
  assign t_r24_c27_2 = p_24_27 << 2;
  assign t_r24_c27_3 = p_24_28 << 1;
  assign t_r24_c27_4 = p_25_27 << 1;
  assign t_r24_c27_5 = t_r24_c27_0 + p_23_26;
  assign t_r24_c27_6 = t_r24_c27_1 + p_23_28;
  assign t_r24_c27_7 = t_r24_c27_2 + t_r24_c27_3;
  assign t_r24_c27_8 = t_r24_c27_4 + p_25_26;
  assign t_r24_c27_9 = t_r24_c27_5 + t_r24_c27_6;
  assign t_r24_c27_10 = t_r24_c27_7 + t_r24_c27_8;
  assign t_r24_c27_11 = t_r24_c27_9 + t_r24_c27_10;
  assign t_r24_c27_12 = t_r24_c27_11 + p_25_28;
  assign out_24_27 = t_r24_c27_12 >> 4;

  assign t_r24_c28_0 = p_23_28 << 1;
  assign t_r24_c28_1 = p_24_27 << 1;
  assign t_r24_c28_2 = p_24_28 << 2;
  assign t_r24_c28_3 = p_24_29 << 1;
  assign t_r24_c28_4 = p_25_28 << 1;
  assign t_r24_c28_5 = t_r24_c28_0 + p_23_27;
  assign t_r24_c28_6 = t_r24_c28_1 + p_23_29;
  assign t_r24_c28_7 = t_r24_c28_2 + t_r24_c28_3;
  assign t_r24_c28_8 = t_r24_c28_4 + p_25_27;
  assign t_r24_c28_9 = t_r24_c28_5 + t_r24_c28_6;
  assign t_r24_c28_10 = t_r24_c28_7 + t_r24_c28_8;
  assign t_r24_c28_11 = t_r24_c28_9 + t_r24_c28_10;
  assign t_r24_c28_12 = t_r24_c28_11 + p_25_29;
  assign out_24_28 = t_r24_c28_12 >> 4;

  assign t_r24_c29_0 = p_23_29 << 1;
  assign t_r24_c29_1 = p_24_28 << 1;
  assign t_r24_c29_2 = p_24_29 << 2;
  assign t_r24_c29_3 = p_24_30 << 1;
  assign t_r24_c29_4 = p_25_29 << 1;
  assign t_r24_c29_5 = t_r24_c29_0 + p_23_28;
  assign t_r24_c29_6 = t_r24_c29_1 + p_23_30;
  assign t_r24_c29_7 = t_r24_c29_2 + t_r24_c29_3;
  assign t_r24_c29_8 = t_r24_c29_4 + p_25_28;
  assign t_r24_c29_9 = t_r24_c29_5 + t_r24_c29_6;
  assign t_r24_c29_10 = t_r24_c29_7 + t_r24_c29_8;
  assign t_r24_c29_11 = t_r24_c29_9 + t_r24_c29_10;
  assign t_r24_c29_12 = t_r24_c29_11 + p_25_30;
  assign out_24_29 = t_r24_c29_12 >> 4;

  assign t_r24_c30_0 = p_23_30 << 1;
  assign t_r24_c30_1 = p_24_29 << 1;
  assign t_r24_c30_2 = p_24_30 << 2;
  assign t_r24_c30_3 = p_24_31 << 1;
  assign t_r24_c30_4 = p_25_30 << 1;
  assign t_r24_c30_5 = t_r24_c30_0 + p_23_29;
  assign t_r24_c30_6 = t_r24_c30_1 + p_23_31;
  assign t_r24_c30_7 = t_r24_c30_2 + t_r24_c30_3;
  assign t_r24_c30_8 = t_r24_c30_4 + p_25_29;
  assign t_r24_c30_9 = t_r24_c30_5 + t_r24_c30_6;
  assign t_r24_c30_10 = t_r24_c30_7 + t_r24_c30_8;
  assign t_r24_c30_11 = t_r24_c30_9 + t_r24_c30_10;
  assign t_r24_c30_12 = t_r24_c30_11 + p_25_31;
  assign out_24_30 = t_r24_c30_12 >> 4;

  assign t_r24_c31_0 = p_23_31 << 1;
  assign t_r24_c31_1 = p_24_30 << 1;
  assign t_r24_c31_2 = p_24_31 << 2;
  assign t_r24_c31_3 = p_24_32 << 1;
  assign t_r24_c31_4 = p_25_31 << 1;
  assign t_r24_c31_5 = t_r24_c31_0 + p_23_30;
  assign t_r24_c31_6 = t_r24_c31_1 + p_23_32;
  assign t_r24_c31_7 = t_r24_c31_2 + t_r24_c31_3;
  assign t_r24_c31_8 = t_r24_c31_4 + p_25_30;
  assign t_r24_c31_9 = t_r24_c31_5 + t_r24_c31_6;
  assign t_r24_c31_10 = t_r24_c31_7 + t_r24_c31_8;
  assign t_r24_c31_11 = t_r24_c31_9 + t_r24_c31_10;
  assign t_r24_c31_12 = t_r24_c31_11 + p_25_32;
  assign out_24_31 = t_r24_c31_12 >> 4;

  assign t_r24_c32_0 = p_23_32 << 1;
  assign t_r24_c32_1 = p_24_31 << 1;
  assign t_r24_c32_2 = p_24_32 << 2;
  assign t_r24_c32_3 = p_24_33 << 1;
  assign t_r24_c32_4 = p_25_32 << 1;
  assign t_r24_c32_5 = t_r24_c32_0 + p_23_31;
  assign t_r24_c32_6 = t_r24_c32_1 + p_23_33;
  assign t_r24_c32_7 = t_r24_c32_2 + t_r24_c32_3;
  assign t_r24_c32_8 = t_r24_c32_4 + p_25_31;
  assign t_r24_c32_9 = t_r24_c32_5 + t_r24_c32_6;
  assign t_r24_c32_10 = t_r24_c32_7 + t_r24_c32_8;
  assign t_r24_c32_11 = t_r24_c32_9 + t_r24_c32_10;
  assign t_r24_c32_12 = t_r24_c32_11 + p_25_33;
  assign out_24_32 = t_r24_c32_12 >> 4;

  assign t_r24_c33_0 = p_23_33 << 1;
  assign t_r24_c33_1 = p_24_32 << 1;
  assign t_r24_c33_2 = p_24_33 << 2;
  assign t_r24_c33_3 = p_24_34 << 1;
  assign t_r24_c33_4 = p_25_33 << 1;
  assign t_r24_c33_5 = t_r24_c33_0 + p_23_32;
  assign t_r24_c33_6 = t_r24_c33_1 + p_23_34;
  assign t_r24_c33_7 = t_r24_c33_2 + t_r24_c33_3;
  assign t_r24_c33_8 = t_r24_c33_4 + p_25_32;
  assign t_r24_c33_9 = t_r24_c33_5 + t_r24_c33_6;
  assign t_r24_c33_10 = t_r24_c33_7 + t_r24_c33_8;
  assign t_r24_c33_11 = t_r24_c33_9 + t_r24_c33_10;
  assign t_r24_c33_12 = t_r24_c33_11 + p_25_34;
  assign out_24_33 = t_r24_c33_12 >> 4;

  assign t_r24_c34_0 = p_23_34 << 1;
  assign t_r24_c34_1 = p_24_33 << 1;
  assign t_r24_c34_2 = p_24_34 << 2;
  assign t_r24_c34_3 = p_24_35 << 1;
  assign t_r24_c34_4 = p_25_34 << 1;
  assign t_r24_c34_5 = t_r24_c34_0 + p_23_33;
  assign t_r24_c34_6 = t_r24_c34_1 + p_23_35;
  assign t_r24_c34_7 = t_r24_c34_2 + t_r24_c34_3;
  assign t_r24_c34_8 = t_r24_c34_4 + p_25_33;
  assign t_r24_c34_9 = t_r24_c34_5 + t_r24_c34_6;
  assign t_r24_c34_10 = t_r24_c34_7 + t_r24_c34_8;
  assign t_r24_c34_11 = t_r24_c34_9 + t_r24_c34_10;
  assign t_r24_c34_12 = t_r24_c34_11 + p_25_35;
  assign out_24_34 = t_r24_c34_12 >> 4;

  assign t_r24_c35_0 = p_23_35 << 1;
  assign t_r24_c35_1 = p_24_34 << 1;
  assign t_r24_c35_2 = p_24_35 << 2;
  assign t_r24_c35_3 = p_24_36 << 1;
  assign t_r24_c35_4 = p_25_35 << 1;
  assign t_r24_c35_5 = t_r24_c35_0 + p_23_34;
  assign t_r24_c35_6 = t_r24_c35_1 + p_23_36;
  assign t_r24_c35_7 = t_r24_c35_2 + t_r24_c35_3;
  assign t_r24_c35_8 = t_r24_c35_4 + p_25_34;
  assign t_r24_c35_9 = t_r24_c35_5 + t_r24_c35_6;
  assign t_r24_c35_10 = t_r24_c35_7 + t_r24_c35_8;
  assign t_r24_c35_11 = t_r24_c35_9 + t_r24_c35_10;
  assign t_r24_c35_12 = t_r24_c35_11 + p_25_36;
  assign out_24_35 = t_r24_c35_12 >> 4;

  assign t_r24_c36_0 = p_23_36 << 1;
  assign t_r24_c36_1 = p_24_35 << 1;
  assign t_r24_c36_2 = p_24_36 << 2;
  assign t_r24_c36_3 = p_24_37 << 1;
  assign t_r24_c36_4 = p_25_36 << 1;
  assign t_r24_c36_5 = t_r24_c36_0 + p_23_35;
  assign t_r24_c36_6 = t_r24_c36_1 + p_23_37;
  assign t_r24_c36_7 = t_r24_c36_2 + t_r24_c36_3;
  assign t_r24_c36_8 = t_r24_c36_4 + p_25_35;
  assign t_r24_c36_9 = t_r24_c36_5 + t_r24_c36_6;
  assign t_r24_c36_10 = t_r24_c36_7 + t_r24_c36_8;
  assign t_r24_c36_11 = t_r24_c36_9 + t_r24_c36_10;
  assign t_r24_c36_12 = t_r24_c36_11 + p_25_37;
  assign out_24_36 = t_r24_c36_12 >> 4;

  assign t_r24_c37_0 = p_23_37 << 1;
  assign t_r24_c37_1 = p_24_36 << 1;
  assign t_r24_c37_2 = p_24_37 << 2;
  assign t_r24_c37_3 = p_24_38 << 1;
  assign t_r24_c37_4 = p_25_37 << 1;
  assign t_r24_c37_5 = t_r24_c37_0 + p_23_36;
  assign t_r24_c37_6 = t_r24_c37_1 + p_23_38;
  assign t_r24_c37_7 = t_r24_c37_2 + t_r24_c37_3;
  assign t_r24_c37_8 = t_r24_c37_4 + p_25_36;
  assign t_r24_c37_9 = t_r24_c37_5 + t_r24_c37_6;
  assign t_r24_c37_10 = t_r24_c37_7 + t_r24_c37_8;
  assign t_r24_c37_11 = t_r24_c37_9 + t_r24_c37_10;
  assign t_r24_c37_12 = t_r24_c37_11 + p_25_38;
  assign out_24_37 = t_r24_c37_12 >> 4;

  assign t_r24_c38_0 = p_23_38 << 1;
  assign t_r24_c38_1 = p_24_37 << 1;
  assign t_r24_c38_2 = p_24_38 << 2;
  assign t_r24_c38_3 = p_24_39 << 1;
  assign t_r24_c38_4 = p_25_38 << 1;
  assign t_r24_c38_5 = t_r24_c38_0 + p_23_37;
  assign t_r24_c38_6 = t_r24_c38_1 + p_23_39;
  assign t_r24_c38_7 = t_r24_c38_2 + t_r24_c38_3;
  assign t_r24_c38_8 = t_r24_c38_4 + p_25_37;
  assign t_r24_c38_9 = t_r24_c38_5 + t_r24_c38_6;
  assign t_r24_c38_10 = t_r24_c38_7 + t_r24_c38_8;
  assign t_r24_c38_11 = t_r24_c38_9 + t_r24_c38_10;
  assign t_r24_c38_12 = t_r24_c38_11 + p_25_39;
  assign out_24_38 = t_r24_c38_12 >> 4;

  assign t_r24_c39_0 = p_23_39 << 1;
  assign t_r24_c39_1 = p_24_38 << 1;
  assign t_r24_c39_2 = p_24_39 << 2;
  assign t_r24_c39_3 = p_24_40 << 1;
  assign t_r24_c39_4 = p_25_39 << 1;
  assign t_r24_c39_5 = t_r24_c39_0 + p_23_38;
  assign t_r24_c39_6 = t_r24_c39_1 + p_23_40;
  assign t_r24_c39_7 = t_r24_c39_2 + t_r24_c39_3;
  assign t_r24_c39_8 = t_r24_c39_4 + p_25_38;
  assign t_r24_c39_9 = t_r24_c39_5 + t_r24_c39_6;
  assign t_r24_c39_10 = t_r24_c39_7 + t_r24_c39_8;
  assign t_r24_c39_11 = t_r24_c39_9 + t_r24_c39_10;
  assign t_r24_c39_12 = t_r24_c39_11 + p_25_40;
  assign out_24_39 = t_r24_c39_12 >> 4;

  assign t_r24_c40_0 = p_23_40 << 1;
  assign t_r24_c40_1 = p_24_39 << 1;
  assign t_r24_c40_2 = p_24_40 << 2;
  assign t_r24_c40_3 = p_24_41 << 1;
  assign t_r24_c40_4 = p_25_40 << 1;
  assign t_r24_c40_5 = t_r24_c40_0 + p_23_39;
  assign t_r24_c40_6 = t_r24_c40_1 + p_23_41;
  assign t_r24_c40_7 = t_r24_c40_2 + t_r24_c40_3;
  assign t_r24_c40_8 = t_r24_c40_4 + p_25_39;
  assign t_r24_c40_9 = t_r24_c40_5 + t_r24_c40_6;
  assign t_r24_c40_10 = t_r24_c40_7 + t_r24_c40_8;
  assign t_r24_c40_11 = t_r24_c40_9 + t_r24_c40_10;
  assign t_r24_c40_12 = t_r24_c40_11 + p_25_41;
  assign out_24_40 = t_r24_c40_12 >> 4;

  assign t_r24_c41_0 = p_23_41 << 1;
  assign t_r24_c41_1 = p_24_40 << 1;
  assign t_r24_c41_2 = p_24_41 << 2;
  assign t_r24_c41_3 = p_24_42 << 1;
  assign t_r24_c41_4 = p_25_41 << 1;
  assign t_r24_c41_5 = t_r24_c41_0 + p_23_40;
  assign t_r24_c41_6 = t_r24_c41_1 + p_23_42;
  assign t_r24_c41_7 = t_r24_c41_2 + t_r24_c41_3;
  assign t_r24_c41_8 = t_r24_c41_4 + p_25_40;
  assign t_r24_c41_9 = t_r24_c41_5 + t_r24_c41_6;
  assign t_r24_c41_10 = t_r24_c41_7 + t_r24_c41_8;
  assign t_r24_c41_11 = t_r24_c41_9 + t_r24_c41_10;
  assign t_r24_c41_12 = t_r24_c41_11 + p_25_42;
  assign out_24_41 = t_r24_c41_12 >> 4;

  assign t_r24_c42_0 = p_23_42 << 1;
  assign t_r24_c42_1 = p_24_41 << 1;
  assign t_r24_c42_2 = p_24_42 << 2;
  assign t_r24_c42_3 = p_24_43 << 1;
  assign t_r24_c42_4 = p_25_42 << 1;
  assign t_r24_c42_5 = t_r24_c42_0 + p_23_41;
  assign t_r24_c42_6 = t_r24_c42_1 + p_23_43;
  assign t_r24_c42_7 = t_r24_c42_2 + t_r24_c42_3;
  assign t_r24_c42_8 = t_r24_c42_4 + p_25_41;
  assign t_r24_c42_9 = t_r24_c42_5 + t_r24_c42_6;
  assign t_r24_c42_10 = t_r24_c42_7 + t_r24_c42_8;
  assign t_r24_c42_11 = t_r24_c42_9 + t_r24_c42_10;
  assign t_r24_c42_12 = t_r24_c42_11 + p_25_43;
  assign out_24_42 = t_r24_c42_12 >> 4;

  assign t_r24_c43_0 = p_23_43 << 1;
  assign t_r24_c43_1 = p_24_42 << 1;
  assign t_r24_c43_2 = p_24_43 << 2;
  assign t_r24_c43_3 = p_24_44 << 1;
  assign t_r24_c43_4 = p_25_43 << 1;
  assign t_r24_c43_5 = t_r24_c43_0 + p_23_42;
  assign t_r24_c43_6 = t_r24_c43_1 + p_23_44;
  assign t_r24_c43_7 = t_r24_c43_2 + t_r24_c43_3;
  assign t_r24_c43_8 = t_r24_c43_4 + p_25_42;
  assign t_r24_c43_9 = t_r24_c43_5 + t_r24_c43_6;
  assign t_r24_c43_10 = t_r24_c43_7 + t_r24_c43_8;
  assign t_r24_c43_11 = t_r24_c43_9 + t_r24_c43_10;
  assign t_r24_c43_12 = t_r24_c43_11 + p_25_44;
  assign out_24_43 = t_r24_c43_12 >> 4;

  assign t_r24_c44_0 = p_23_44 << 1;
  assign t_r24_c44_1 = p_24_43 << 1;
  assign t_r24_c44_2 = p_24_44 << 2;
  assign t_r24_c44_3 = p_24_45 << 1;
  assign t_r24_c44_4 = p_25_44 << 1;
  assign t_r24_c44_5 = t_r24_c44_0 + p_23_43;
  assign t_r24_c44_6 = t_r24_c44_1 + p_23_45;
  assign t_r24_c44_7 = t_r24_c44_2 + t_r24_c44_3;
  assign t_r24_c44_8 = t_r24_c44_4 + p_25_43;
  assign t_r24_c44_9 = t_r24_c44_5 + t_r24_c44_6;
  assign t_r24_c44_10 = t_r24_c44_7 + t_r24_c44_8;
  assign t_r24_c44_11 = t_r24_c44_9 + t_r24_c44_10;
  assign t_r24_c44_12 = t_r24_c44_11 + p_25_45;
  assign out_24_44 = t_r24_c44_12 >> 4;

  assign t_r24_c45_0 = p_23_45 << 1;
  assign t_r24_c45_1 = p_24_44 << 1;
  assign t_r24_c45_2 = p_24_45 << 2;
  assign t_r24_c45_3 = p_24_46 << 1;
  assign t_r24_c45_4 = p_25_45 << 1;
  assign t_r24_c45_5 = t_r24_c45_0 + p_23_44;
  assign t_r24_c45_6 = t_r24_c45_1 + p_23_46;
  assign t_r24_c45_7 = t_r24_c45_2 + t_r24_c45_3;
  assign t_r24_c45_8 = t_r24_c45_4 + p_25_44;
  assign t_r24_c45_9 = t_r24_c45_5 + t_r24_c45_6;
  assign t_r24_c45_10 = t_r24_c45_7 + t_r24_c45_8;
  assign t_r24_c45_11 = t_r24_c45_9 + t_r24_c45_10;
  assign t_r24_c45_12 = t_r24_c45_11 + p_25_46;
  assign out_24_45 = t_r24_c45_12 >> 4;

  assign t_r24_c46_0 = p_23_46 << 1;
  assign t_r24_c46_1 = p_24_45 << 1;
  assign t_r24_c46_2 = p_24_46 << 2;
  assign t_r24_c46_3 = p_24_47 << 1;
  assign t_r24_c46_4 = p_25_46 << 1;
  assign t_r24_c46_5 = t_r24_c46_0 + p_23_45;
  assign t_r24_c46_6 = t_r24_c46_1 + p_23_47;
  assign t_r24_c46_7 = t_r24_c46_2 + t_r24_c46_3;
  assign t_r24_c46_8 = t_r24_c46_4 + p_25_45;
  assign t_r24_c46_9 = t_r24_c46_5 + t_r24_c46_6;
  assign t_r24_c46_10 = t_r24_c46_7 + t_r24_c46_8;
  assign t_r24_c46_11 = t_r24_c46_9 + t_r24_c46_10;
  assign t_r24_c46_12 = t_r24_c46_11 + p_25_47;
  assign out_24_46 = t_r24_c46_12 >> 4;

  assign t_r24_c47_0 = p_23_47 << 1;
  assign t_r24_c47_1 = p_24_46 << 1;
  assign t_r24_c47_2 = p_24_47 << 2;
  assign t_r24_c47_3 = p_24_48 << 1;
  assign t_r24_c47_4 = p_25_47 << 1;
  assign t_r24_c47_5 = t_r24_c47_0 + p_23_46;
  assign t_r24_c47_6 = t_r24_c47_1 + p_23_48;
  assign t_r24_c47_7 = t_r24_c47_2 + t_r24_c47_3;
  assign t_r24_c47_8 = t_r24_c47_4 + p_25_46;
  assign t_r24_c47_9 = t_r24_c47_5 + t_r24_c47_6;
  assign t_r24_c47_10 = t_r24_c47_7 + t_r24_c47_8;
  assign t_r24_c47_11 = t_r24_c47_9 + t_r24_c47_10;
  assign t_r24_c47_12 = t_r24_c47_11 + p_25_48;
  assign out_24_47 = t_r24_c47_12 >> 4;

  assign t_r24_c48_0 = p_23_48 << 1;
  assign t_r24_c48_1 = p_24_47 << 1;
  assign t_r24_c48_2 = p_24_48 << 2;
  assign t_r24_c48_3 = p_24_49 << 1;
  assign t_r24_c48_4 = p_25_48 << 1;
  assign t_r24_c48_5 = t_r24_c48_0 + p_23_47;
  assign t_r24_c48_6 = t_r24_c48_1 + p_23_49;
  assign t_r24_c48_7 = t_r24_c48_2 + t_r24_c48_3;
  assign t_r24_c48_8 = t_r24_c48_4 + p_25_47;
  assign t_r24_c48_9 = t_r24_c48_5 + t_r24_c48_6;
  assign t_r24_c48_10 = t_r24_c48_7 + t_r24_c48_8;
  assign t_r24_c48_11 = t_r24_c48_9 + t_r24_c48_10;
  assign t_r24_c48_12 = t_r24_c48_11 + p_25_49;
  assign out_24_48 = t_r24_c48_12 >> 4;

  assign t_r24_c49_0 = p_23_49 << 1;
  assign t_r24_c49_1 = p_24_48 << 1;
  assign t_r24_c49_2 = p_24_49 << 2;
  assign t_r24_c49_3 = p_24_50 << 1;
  assign t_r24_c49_4 = p_25_49 << 1;
  assign t_r24_c49_5 = t_r24_c49_0 + p_23_48;
  assign t_r24_c49_6 = t_r24_c49_1 + p_23_50;
  assign t_r24_c49_7 = t_r24_c49_2 + t_r24_c49_3;
  assign t_r24_c49_8 = t_r24_c49_4 + p_25_48;
  assign t_r24_c49_9 = t_r24_c49_5 + t_r24_c49_6;
  assign t_r24_c49_10 = t_r24_c49_7 + t_r24_c49_8;
  assign t_r24_c49_11 = t_r24_c49_9 + t_r24_c49_10;
  assign t_r24_c49_12 = t_r24_c49_11 + p_25_50;
  assign out_24_49 = t_r24_c49_12 >> 4;

  assign t_r24_c50_0 = p_23_50 << 1;
  assign t_r24_c50_1 = p_24_49 << 1;
  assign t_r24_c50_2 = p_24_50 << 2;
  assign t_r24_c50_3 = p_24_51 << 1;
  assign t_r24_c50_4 = p_25_50 << 1;
  assign t_r24_c50_5 = t_r24_c50_0 + p_23_49;
  assign t_r24_c50_6 = t_r24_c50_1 + p_23_51;
  assign t_r24_c50_7 = t_r24_c50_2 + t_r24_c50_3;
  assign t_r24_c50_8 = t_r24_c50_4 + p_25_49;
  assign t_r24_c50_9 = t_r24_c50_5 + t_r24_c50_6;
  assign t_r24_c50_10 = t_r24_c50_7 + t_r24_c50_8;
  assign t_r24_c50_11 = t_r24_c50_9 + t_r24_c50_10;
  assign t_r24_c50_12 = t_r24_c50_11 + p_25_51;
  assign out_24_50 = t_r24_c50_12 >> 4;

  assign t_r24_c51_0 = p_23_51 << 1;
  assign t_r24_c51_1 = p_24_50 << 1;
  assign t_r24_c51_2 = p_24_51 << 2;
  assign t_r24_c51_3 = p_24_52 << 1;
  assign t_r24_c51_4 = p_25_51 << 1;
  assign t_r24_c51_5 = t_r24_c51_0 + p_23_50;
  assign t_r24_c51_6 = t_r24_c51_1 + p_23_52;
  assign t_r24_c51_7 = t_r24_c51_2 + t_r24_c51_3;
  assign t_r24_c51_8 = t_r24_c51_4 + p_25_50;
  assign t_r24_c51_9 = t_r24_c51_5 + t_r24_c51_6;
  assign t_r24_c51_10 = t_r24_c51_7 + t_r24_c51_8;
  assign t_r24_c51_11 = t_r24_c51_9 + t_r24_c51_10;
  assign t_r24_c51_12 = t_r24_c51_11 + p_25_52;
  assign out_24_51 = t_r24_c51_12 >> 4;

  assign t_r24_c52_0 = p_23_52 << 1;
  assign t_r24_c52_1 = p_24_51 << 1;
  assign t_r24_c52_2 = p_24_52 << 2;
  assign t_r24_c52_3 = p_24_53 << 1;
  assign t_r24_c52_4 = p_25_52 << 1;
  assign t_r24_c52_5 = t_r24_c52_0 + p_23_51;
  assign t_r24_c52_6 = t_r24_c52_1 + p_23_53;
  assign t_r24_c52_7 = t_r24_c52_2 + t_r24_c52_3;
  assign t_r24_c52_8 = t_r24_c52_4 + p_25_51;
  assign t_r24_c52_9 = t_r24_c52_5 + t_r24_c52_6;
  assign t_r24_c52_10 = t_r24_c52_7 + t_r24_c52_8;
  assign t_r24_c52_11 = t_r24_c52_9 + t_r24_c52_10;
  assign t_r24_c52_12 = t_r24_c52_11 + p_25_53;
  assign out_24_52 = t_r24_c52_12 >> 4;

  assign t_r24_c53_0 = p_23_53 << 1;
  assign t_r24_c53_1 = p_24_52 << 1;
  assign t_r24_c53_2 = p_24_53 << 2;
  assign t_r24_c53_3 = p_24_54 << 1;
  assign t_r24_c53_4 = p_25_53 << 1;
  assign t_r24_c53_5 = t_r24_c53_0 + p_23_52;
  assign t_r24_c53_6 = t_r24_c53_1 + p_23_54;
  assign t_r24_c53_7 = t_r24_c53_2 + t_r24_c53_3;
  assign t_r24_c53_8 = t_r24_c53_4 + p_25_52;
  assign t_r24_c53_9 = t_r24_c53_5 + t_r24_c53_6;
  assign t_r24_c53_10 = t_r24_c53_7 + t_r24_c53_8;
  assign t_r24_c53_11 = t_r24_c53_9 + t_r24_c53_10;
  assign t_r24_c53_12 = t_r24_c53_11 + p_25_54;
  assign out_24_53 = t_r24_c53_12 >> 4;

  assign t_r24_c54_0 = p_23_54 << 1;
  assign t_r24_c54_1 = p_24_53 << 1;
  assign t_r24_c54_2 = p_24_54 << 2;
  assign t_r24_c54_3 = p_24_55 << 1;
  assign t_r24_c54_4 = p_25_54 << 1;
  assign t_r24_c54_5 = t_r24_c54_0 + p_23_53;
  assign t_r24_c54_6 = t_r24_c54_1 + p_23_55;
  assign t_r24_c54_7 = t_r24_c54_2 + t_r24_c54_3;
  assign t_r24_c54_8 = t_r24_c54_4 + p_25_53;
  assign t_r24_c54_9 = t_r24_c54_5 + t_r24_c54_6;
  assign t_r24_c54_10 = t_r24_c54_7 + t_r24_c54_8;
  assign t_r24_c54_11 = t_r24_c54_9 + t_r24_c54_10;
  assign t_r24_c54_12 = t_r24_c54_11 + p_25_55;
  assign out_24_54 = t_r24_c54_12 >> 4;

  assign t_r24_c55_0 = p_23_55 << 1;
  assign t_r24_c55_1 = p_24_54 << 1;
  assign t_r24_c55_2 = p_24_55 << 2;
  assign t_r24_c55_3 = p_24_56 << 1;
  assign t_r24_c55_4 = p_25_55 << 1;
  assign t_r24_c55_5 = t_r24_c55_0 + p_23_54;
  assign t_r24_c55_6 = t_r24_c55_1 + p_23_56;
  assign t_r24_c55_7 = t_r24_c55_2 + t_r24_c55_3;
  assign t_r24_c55_8 = t_r24_c55_4 + p_25_54;
  assign t_r24_c55_9 = t_r24_c55_5 + t_r24_c55_6;
  assign t_r24_c55_10 = t_r24_c55_7 + t_r24_c55_8;
  assign t_r24_c55_11 = t_r24_c55_9 + t_r24_c55_10;
  assign t_r24_c55_12 = t_r24_c55_11 + p_25_56;
  assign out_24_55 = t_r24_c55_12 >> 4;

  assign t_r24_c56_0 = p_23_56 << 1;
  assign t_r24_c56_1 = p_24_55 << 1;
  assign t_r24_c56_2 = p_24_56 << 2;
  assign t_r24_c56_3 = p_24_57 << 1;
  assign t_r24_c56_4 = p_25_56 << 1;
  assign t_r24_c56_5 = t_r24_c56_0 + p_23_55;
  assign t_r24_c56_6 = t_r24_c56_1 + p_23_57;
  assign t_r24_c56_7 = t_r24_c56_2 + t_r24_c56_3;
  assign t_r24_c56_8 = t_r24_c56_4 + p_25_55;
  assign t_r24_c56_9 = t_r24_c56_5 + t_r24_c56_6;
  assign t_r24_c56_10 = t_r24_c56_7 + t_r24_c56_8;
  assign t_r24_c56_11 = t_r24_c56_9 + t_r24_c56_10;
  assign t_r24_c56_12 = t_r24_c56_11 + p_25_57;
  assign out_24_56 = t_r24_c56_12 >> 4;

  assign t_r24_c57_0 = p_23_57 << 1;
  assign t_r24_c57_1 = p_24_56 << 1;
  assign t_r24_c57_2 = p_24_57 << 2;
  assign t_r24_c57_3 = p_24_58 << 1;
  assign t_r24_c57_4 = p_25_57 << 1;
  assign t_r24_c57_5 = t_r24_c57_0 + p_23_56;
  assign t_r24_c57_6 = t_r24_c57_1 + p_23_58;
  assign t_r24_c57_7 = t_r24_c57_2 + t_r24_c57_3;
  assign t_r24_c57_8 = t_r24_c57_4 + p_25_56;
  assign t_r24_c57_9 = t_r24_c57_5 + t_r24_c57_6;
  assign t_r24_c57_10 = t_r24_c57_7 + t_r24_c57_8;
  assign t_r24_c57_11 = t_r24_c57_9 + t_r24_c57_10;
  assign t_r24_c57_12 = t_r24_c57_11 + p_25_58;
  assign out_24_57 = t_r24_c57_12 >> 4;

  assign t_r24_c58_0 = p_23_58 << 1;
  assign t_r24_c58_1 = p_24_57 << 1;
  assign t_r24_c58_2 = p_24_58 << 2;
  assign t_r24_c58_3 = p_24_59 << 1;
  assign t_r24_c58_4 = p_25_58 << 1;
  assign t_r24_c58_5 = t_r24_c58_0 + p_23_57;
  assign t_r24_c58_6 = t_r24_c58_1 + p_23_59;
  assign t_r24_c58_7 = t_r24_c58_2 + t_r24_c58_3;
  assign t_r24_c58_8 = t_r24_c58_4 + p_25_57;
  assign t_r24_c58_9 = t_r24_c58_5 + t_r24_c58_6;
  assign t_r24_c58_10 = t_r24_c58_7 + t_r24_c58_8;
  assign t_r24_c58_11 = t_r24_c58_9 + t_r24_c58_10;
  assign t_r24_c58_12 = t_r24_c58_11 + p_25_59;
  assign out_24_58 = t_r24_c58_12 >> 4;

  assign t_r24_c59_0 = p_23_59 << 1;
  assign t_r24_c59_1 = p_24_58 << 1;
  assign t_r24_c59_2 = p_24_59 << 2;
  assign t_r24_c59_3 = p_24_60 << 1;
  assign t_r24_c59_4 = p_25_59 << 1;
  assign t_r24_c59_5 = t_r24_c59_0 + p_23_58;
  assign t_r24_c59_6 = t_r24_c59_1 + p_23_60;
  assign t_r24_c59_7 = t_r24_c59_2 + t_r24_c59_3;
  assign t_r24_c59_8 = t_r24_c59_4 + p_25_58;
  assign t_r24_c59_9 = t_r24_c59_5 + t_r24_c59_6;
  assign t_r24_c59_10 = t_r24_c59_7 + t_r24_c59_8;
  assign t_r24_c59_11 = t_r24_c59_9 + t_r24_c59_10;
  assign t_r24_c59_12 = t_r24_c59_11 + p_25_60;
  assign out_24_59 = t_r24_c59_12 >> 4;

  assign t_r24_c60_0 = p_23_60 << 1;
  assign t_r24_c60_1 = p_24_59 << 1;
  assign t_r24_c60_2 = p_24_60 << 2;
  assign t_r24_c60_3 = p_24_61 << 1;
  assign t_r24_c60_4 = p_25_60 << 1;
  assign t_r24_c60_5 = t_r24_c60_0 + p_23_59;
  assign t_r24_c60_6 = t_r24_c60_1 + p_23_61;
  assign t_r24_c60_7 = t_r24_c60_2 + t_r24_c60_3;
  assign t_r24_c60_8 = t_r24_c60_4 + p_25_59;
  assign t_r24_c60_9 = t_r24_c60_5 + t_r24_c60_6;
  assign t_r24_c60_10 = t_r24_c60_7 + t_r24_c60_8;
  assign t_r24_c60_11 = t_r24_c60_9 + t_r24_c60_10;
  assign t_r24_c60_12 = t_r24_c60_11 + p_25_61;
  assign out_24_60 = t_r24_c60_12 >> 4;

  assign t_r24_c61_0 = p_23_61 << 1;
  assign t_r24_c61_1 = p_24_60 << 1;
  assign t_r24_c61_2 = p_24_61 << 2;
  assign t_r24_c61_3 = p_24_62 << 1;
  assign t_r24_c61_4 = p_25_61 << 1;
  assign t_r24_c61_5 = t_r24_c61_0 + p_23_60;
  assign t_r24_c61_6 = t_r24_c61_1 + p_23_62;
  assign t_r24_c61_7 = t_r24_c61_2 + t_r24_c61_3;
  assign t_r24_c61_8 = t_r24_c61_4 + p_25_60;
  assign t_r24_c61_9 = t_r24_c61_5 + t_r24_c61_6;
  assign t_r24_c61_10 = t_r24_c61_7 + t_r24_c61_8;
  assign t_r24_c61_11 = t_r24_c61_9 + t_r24_c61_10;
  assign t_r24_c61_12 = t_r24_c61_11 + p_25_62;
  assign out_24_61 = t_r24_c61_12 >> 4;

  assign t_r24_c62_0 = p_23_62 << 1;
  assign t_r24_c62_1 = p_24_61 << 1;
  assign t_r24_c62_2 = p_24_62 << 2;
  assign t_r24_c62_3 = p_24_63 << 1;
  assign t_r24_c62_4 = p_25_62 << 1;
  assign t_r24_c62_5 = t_r24_c62_0 + p_23_61;
  assign t_r24_c62_6 = t_r24_c62_1 + p_23_63;
  assign t_r24_c62_7 = t_r24_c62_2 + t_r24_c62_3;
  assign t_r24_c62_8 = t_r24_c62_4 + p_25_61;
  assign t_r24_c62_9 = t_r24_c62_5 + t_r24_c62_6;
  assign t_r24_c62_10 = t_r24_c62_7 + t_r24_c62_8;
  assign t_r24_c62_11 = t_r24_c62_9 + t_r24_c62_10;
  assign t_r24_c62_12 = t_r24_c62_11 + p_25_63;
  assign out_24_62 = t_r24_c62_12 >> 4;

  assign t_r24_c63_0 = p_23_63 << 1;
  assign t_r24_c63_1 = p_24_62 << 1;
  assign t_r24_c63_2 = p_24_63 << 2;
  assign t_r24_c63_3 = p_24_64 << 1;
  assign t_r24_c63_4 = p_25_63 << 1;
  assign t_r24_c63_5 = t_r24_c63_0 + p_23_62;
  assign t_r24_c63_6 = t_r24_c63_1 + p_23_64;
  assign t_r24_c63_7 = t_r24_c63_2 + t_r24_c63_3;
  assign t_r24_c63_8 = t_r24_c63_4 + p_25_62;
  assign t_r24_c63_9 = t_r24_c63_5 + t_r24_c63_6;
  assign t_r24_c63_10 = t_r24_c63_7 + t_r24_c63_8;
  assign t_r24_c63_11 = t_r24_c63_9 + t_r24_c63_10;
  assign t_r24_c63_12 = t_r24_c63_11 + p_25_64;
  assign out_24_63 = t_r24_c63_12 >> 4;

  assign t_r24_c64_0 = p_23_64 << 1;
  assign t_r24_c64_1 = p_24_63 << 1;
  assign t_r24_c64_2 = p_24_64 << 2;
  assign t_r24_c64_3 = p_24_65 << 1;
  assign t_r24_c64_4 = p_25_64 << 1;
  assign t_r24_c64_5 = t_r24_c64_0 + p_23_63;
  assign t_r24_c64_6 = t_r24_c64_1 + p_23_65;
  assign t_r24_c64_7 = t_r24_c64_2 + t_r24_c64_3;
  assign t_r24_c64_8 = t_r24_c64_4 + p_25_63;
  assign t_r24_c64_9 = t_r24_c64_5 + t_r24_c64_6;
  assign t_r24_c64_10 = t_r24_c64_7 + t_r24_c64_8;
  assign t_r24_c64_11 = t_r24_c64_9 + t_r24_c64_10;
  assign t_r24_c64_12 = t_r24_c64_11 + p_25_65;
  assign out_24_64 = t_r24_c64_12 >> 4;

  assign t_r25_c1_0 = p_24_1 << 1;
  assign t_r25_c1_1 = p_25_0 << 1;
  assign t_r25_c1_2 = p_25_1 << 2;
  assign t_r25_c1_3 = p_25_2 << 1;
  assign t_r25_c1_4 = p_26_1 << 1;
  assign t_r25_c1_5 = t_r25_c1_0 + p_24_0;
  assign t_r25_c1_6 = t_r25_c1_1 + p_24_2;
  assign t_r25_c1_7 = t_r25_c1_2 + t_r25_c1_3;
  assign t_r25_c1_8 = t_r25_c1_4 + p_26_0;
  assign t_r25_c1_9 = t_r25_c1_5 + t_r25_c1_6;
  assign t_r25_c1_10 = t_r25_c1_7 + t_r25_c1_8;
  assign t_r25_c1_11 = t_r25_c1_9 + t_r25_c1_10;
  assign t_r25_c1_12 = t_r25_c1_11 + p_26_2;
  assign out_25_1 = t_r25_c1_12 >> 4;

  assign t_r25_c2_0 = p_24_2 << 1;
  assign t_r25_c2_1 = p_25_1 << 1;
  assign t_r25_c2_2 = p_25_2 << 2;
  assign t_r25_c2_3 = p_25_3 << 1;
  assign t_r25_c2_4 = p_26_2 << 1;
  assign t_r25_c2_5 = t_r25_c2_0 + p_24_1;
  assign t_r25_c2_6 = t_r25_c2_1 + p_24_3;
  assign t_r25_c2_7 = t_r25_c2_2 + t_r25_c2_3;
  assign t_r25_c2_8 = t_r25_c2_4 + p_26_1;
  assign t_r25_c2_9 = t_r25_c2_5 + t_r25_c2_6;
  assign t_r25_c2_10 = t_r25_c2_7 + t_r25_c2_8;
  assign t_r25_c2_11 = t_r25_c2_9 + t_r25_c2_10;
  assign t_r25_c2_12 = t_r25_c2_11 + p_26_3;
  assign out_25_2 = t_r25_c2_12 >> 4;

  assign t_r25_c3_0 = p_24_3 << 1;
  assign t_r25_c3_1 = p_25_2 << 1;
  assign t_r25_c3_2 = p_25_3 << 2;
  assign t_r25_c3_3 = p_25_4 << 1;
  assign t_r25_c3_4 = p_26_3 << 1;
  assign t_r25_c3_5 = t_r25_c3_0 + p_24_2;
  assign t_r25_c3_6 = t_r25_c3_1 + p_24_4;
  assign t_r25_c3_7 = t_r25_c3_2 + t_r25_c3_3;
  assign t_r25_c3_8 = t_r25_c3_4 + p_26_2;
  assign t_r25_c3_9 = t_r25_c3_5 + t_r25_c3_6;
  assign t_r25_c3_10 = t_r25_c3_7 + t_r25_c3_8;
  assign t_r25_c3_11 = t_r25_c3_9 + t_r25_c3_10;
  assign t_r25_c3_12 = t_r25_c3_11 + p_26_4;
  assign out_25_3 = t_r25_c3_12 >> 4;

  assign t_r25_c4_0 = p_24_4 << 1;
  assign t_r25_c4_1 = p_25_3 << 1;
  assign t_r25_c4_2 = p_25_4 << 2;
  assign t_r25_c4_3 = p_25_5 << 1;
  assign t_r25_c4_4 = p_26_4 << 1;
  assign t_r25_c4_5 = t_r25_c4_0 + p_24_3;
  assign t_r25_c4_6 = t_r25_c4_1 + p_24_5;
  assign t_r25_c4_7 = t_r25_c4_2 + t_r25_c4_3;
  assign t_r25_c4_8 = t_r25_c4_4 + p_26_3;
  assign t_r25_c4_9 = t_r25_c4_5 + t_r25_c4_6;
  assign t_r25_c4_10 = t_r25_c4_7 + t_r25_c4_8;
  assign t_r25_c4_11 = t_r25_c4_9 + t_r25_c4_10;
  assign t_r25_c4_12 = t_r25_c4_11 + p_26_5;
  assign out_25_4 = t_r25_c4_12 >> 4;

  assign t_r25_c5_0 = p_24_5 << 1;
  assign t_r25_c5_1 = p_25_4 << 1;
  assign t_r25_c5_2 = p_25_5 << 2;
  assign t_r25_c5_3 = p_25_6 << 1;
  assign t_r25_c5_4 = p_26_5 << 1;
  assign t_r25_c5_5 = t_r25_c5_0 + p_24_4;
  assign t_r25_c5_6 = t_r25_c5_1 + p_24_6;
  assign t_r25_c5_7 = t_r25_c5_2 + t_r25_c5_3;
  assign t_r25_c5_8 = t_r25_c5_4 + p_26_4;
  assign t_r25_c5_9 = t_r25_c5_5 + t_r25_c5_6;
  assign t_r25_c5_10 = t_r25_c5_7 + t_r25_c5_8;
  assign t_r25_c5_11 = t_r25_c5_9 + t_r25_c5_10;
  assign t_r25_c5_12 = t_r25_c5_11 + p_26_6;
  assign out_25_5 = t_r25_c5_12 >> 4;

  assign t_r25_c6_0 = p_24_6 << 1;
  assign t_r25_c6_1 = p_25_5 << 1;
  assign t_r25_c6_2 = p_25_6 << 2;
  assign t_r25_c6_3 = p_25_7 << 1;
  assign t_r25_c6_4 = p_26_6 << 1;
  assign t_r25_c6_5 = t_r25_c6_0 + p_24_5;
  assign t_r25_c6_6 = t_r25_c6_1 + p_24_7;
  assign t_r25_c6_7 = t_r25_c6_2 + t_r25_c6_3;
  assign t_r25_c6_8 = t_r25_c6_4 + p_26_5;
  assign t_r25_c6_9 = t_r25_c6_5 + t_r25_c6_6;
  assign t_r25_c6_10 = t_r25_c6_7 + t_r25_c6_8;
  assign t_r25_c6_11 = t_r25_c6_9 + t_r25_c6_10;
  assign t_r25_c6_12 = t_r25_c6_11 + p_26_7;
  assign out_25_6 = t_r25_c6_12 >> 4;

  assign t_r25_c7_0 = p_24_7 << 1;
  assign t_r25_c7_1 = p_25_6 << 1;
  assign t_r25_c7_2 = p_25_7 << 2;
  assign t_r25_c7_3 = p_25_8 << 1;
  assign t_r25_c7_4 = p_26_7 << 1;
  assign t_r25_c7_5 = t_r25_c7_0 + p_24_6;
  assign t_r25_c7_6 = t_r25_c7_1 + p_24_8;
  assign t_r25_c7_7 = t_r25_c7_2 + t_r25_c7_3;
  assign t_r25_c7_8 = t_r25_c7_4 + p_26_6;
  assign t_r25_c7_9 = t_r25_c7_5 + t_r25_c7_6;
  assign t_r25_c7_10 = t_r25_c7_7 + t_r25_c7_8;
  assign t_r25_c7_11 = t_r25_c7_9 + t_r25_c7_10;
  assign t_r25_c7_12 = t_r25_c7_11 + p_26_8;
  assign out_25_7 = t_r25_c7_12 >> 4;

  assign t_r25_c8_0 = p_24_8 << 1;
  assign t_r25_c8_1 = p_25_7 << 1;
  assign t_r25_c8_2 = p_25_8 << 2;
  assign t_r25_c8_3 = p_25_9 << 1;
  assign t_r25_c8_4 = p_26_8 << 1;
  assign t_r25_c8_5 = t_r25_c8_0 + p_24_7;
  assign t_r25_c8_6 = t_r25_c8_1 + p_24_9;
  assign t_r25_c8_7 = t_r25_c8_2 + t_r25_c8_3;
  assign t_r25_c8_8 = t_r25_c8_4 + p_26_7;
  assign t_r25_c8_9 = t_r25_c8_5 + t_r25_c8_6;
  assign t_r25_c8_10 = t_r25_c8_7 + t_r25_c8_8;
  assign t_r25_c8_11 = t_r25_c8_9 + t_r25_c8_10;
  assign t_r25_c8_12 = t_r25_c8_11 + p_26_9;
  assign out_25_8 = t_r25_c8_12 >> 4;

  assign t_r25_c9_0 = p_24_9 << 1;
  assign t_r25_c9_1 = p_25_8 << 1;
  assign t_r25_c9_2 = p_25_9 << 2;
  assign t_r25_c9_3 = p_25_10 << 1;
  assign t_r25_c9_4 = p_26_9 << 1;
  assign t_r25_c9_5 = t_r25_c9_0 + p_24_8;
  assign t_r25_c9_6 = t_r25_c9_1 + p_24_10;
  assign t_r25_c9_7 = t_r25_c9_2 + t_r25_c9_3;
  assign t_r25_c9_8 = t_r25_c9_4 + p_26_8;
  assign t_r25_c9_9 = t_r25_c9_5 + t_r25_c9_6;
  assign t_r25_c9_10 = t_r25_c9_7 + t_r25_c9_8;
  assign t_r25_c9_11 = t_r25_c9_9 + t_r25_c9_10;
  assign t_r25_c9_12 = t_r25_c9_11 + p_26_10;
  assign out_25_9 = t_r25_c9_12 >> 4;

  assign t_r25_c10_0 = p_24_10 << 1;
  assign t_r25_c10_1 = p_25_9 << 1;
  assign t_r25_c10_2 = p_25_10 << 2;
  assign t_r25_c10_3 = p_25_11 << 1;
  assign t_r25_c10_4 = p_26_10 << 1;
  assign t_r25_c10_5 = t_r25_c10_0 + p_24_9;
  assign t_r25_c10_6 = t_r25_c10_1 + p_24_11;
  assign t_r25_c10_7 = t_r25_c10_2 + t_r25_c10_3;
  assign t_r25_c10_8 = t_r25_c10_4 + p_26_9;
  assign t_r25_c10_9 = t_r25_c10_5 + t_r25_c10_6;
  assign t_r25_c10_10 = t_r25_c10_7 + t_r25_c10_8;
  assign t_r25_c10_11 = t_r25_c10_9 + t_r25_c10_10;
  assign t_r25_c10_12 = t_r25_c10_11 + p_26_11;
  assign out_25_10 = t_r25_c10_12 >> 4;

  assign t_r25_c11_0 = p_24_11 << 1;
  assign t_r25_c11_1 = p_25_10 << 1;
  assign t_r25_c11_2 = p_25_11 << 2;
  assign t_r25_c11_3 = p_25_12 << 1;
  assign t_r25_c11_4 = p_26_11 << 1;
  assign t_r25_c11_5 = t_r25_c11_0 + p_24_10;
  assign t_r25_c11_6 = t_r25_c11_1 + p_24_12;
  assign t_r25_c11_7 = t_r25_c11_2 + t_r25_c11_3;
  assign t_r25_c11_8 = t_r25_c11_4 + p_26_10;
  assign t_r25_c11_9 = t_r25_c11_5 + t_r25_c11_6;
  assign t_r25_c11_10 = t_r25_c11_7 + t_r25_c11_8;
  assign t_r25_c11_11 = t_r25_c11_9 + t_r25_c11_10;
  assign t_r25_c11_12 = t_r25_c11_11 + p_26_12;
  assign out_25_11 = t_r25_c11_12 >> 4;

  assign t_r25_c12_0 = p_24_12 << 1;
  assign t_r25_c12_1 = p_25_11 << 1;
  assign t_r25_c12_2 = p_25_12 << 2;
  assign t_r25_c12_3 = p_25_13 << 1;
  assign t_r25_c12_4 = p_26_12 << 1;
  assign t_r25_c12_5 = t_r25_c12_0 + p_24_11;
  assign t_r25_c12_6 = t_r25_c12_1 + p_24_13;
  assign t_r25_c12_7 = t_r25_c12_2 + t_r25_c12_3;
  assign t_r25_c12_8 = t_r25_c12_4 + p_26_11;
  assign t_r25_c12_9 = t_r25_c12_5 + t_r25_c12_6;
  assign t_r25_c12_10 = t_r25_c12_7 + t_r25_c12_8;
  assign t_r25_c12_11 = t_r25_c12_9 + t_r25_c12_10;
  assign t_r25_c12_12 = t_r25_c12_11 + p_26_13;
  assign out_25_12 = t_r25_c12_12 >> 4;

  assign t_r25_c13_0 = p_24_13 << 1;
  assign t_r25_c13_1 = p_25_12 << 1;
  assign t_r25_c13_2 = p_25_13 << 2;
  assign t_r25_c13_3 = p_25_14 << 1;
  assign t_r25_c13_4 = p_26_13 << 1;
  assign t_r25_c13_5 = t_r25_c13_0 + p_24_12;
  assign t_r25_c13_6 = t_r25_c13_1 + p_24_14;
  assign t_r25_c13_7 = t_r25_c13_2 + t_r25_c13_3;
  assign t_r25_c13_8 = t_r25_c13_4 + p_26_12;
  assign t_r25_c13_9 = t_r25_c13_5 + t_r25_c13_6;
  assign t_r25_c13_10 = t_r25_c13_7 + t_r25_c13_8;
  assign t_r25_c13_11 = t_r25_c13_9 + t_r25_c13_10;
  assign t_r25_c13_12 = t_r25_c13_11 + p_26_14;
  assign out_25_13 = t_r25_c13_12 >> 4;

  assign t_r25_c14_0 = p_24_14 << 1;
  assign t_r25_c14_1 = p_25_13 << 1;
  assign t_r25_c14_2 = p_25_14 << 2;
  assign t_r25_c14_3 = p_25_15 << 1;
  assign t_r25_c14_4 = p_26_14 << 1;
  assign t_r25_c14_5 = t_r25_c14_0 + p_24_13;
  assign t_r25_c14_6 = t_r25_c14_1 + p_24_15;
  assign t_r25_c14_7 = t_r25_c14_2 + t_r25_c14_3;
  assign t_r25_c14_8 = t_r25_c14_4 + p_26_13;
  assign t_r25_c14_9 = t_r25_c14_5 + t_r25_c14_6;
  assign t_r25_c14_10 = t_r25_c14_7 + t_r25_c14_8;
  assign t_r25_c14_11 = t_r25_c14_9 + t_r25_c14_10;
  assign t_r25_c14_12 = t_r25_c14_11 + p_26_15;
  assign out_25_14 = t_r25_c14_12 >> 4;

  assign t_r25_c15_0 = p_24_15 << 1;
  assign t_r25_c15_1 = p_25_14 << 1;
  assign t_r25_c15_2 = p_25_15 << 2;
  assign t_r25_c15_3 = p_25_16 << 1;
  assign t_r25_c15_4 = p_26_15 << 1;
  assign t_r25_c15_5 = t_r25_c15_0 + p_24_14;
  assign t_r25_c15_6 = t_r25_c15_1 + p_24_16;
  assign t_r25_c15_7 = t_r25_c15_2 + t_r25_c15_3;
  assign t_r25_c15_8 = t_r25_c15_4 + p_26_14;
  assign t_r25_c15_9 = t_r25_c15_5 + t_r25_c15_6;
  assign t_r25_c15_10 = t_r25_c15_7 + t_r25_c15_8;
  assign t_r25_c15_11 = t_r25_c15_9 + t_r25_c15_10;
  assign t_r25_c15_12 = t_r25_c15_11 + p_26_16;
  assign out_25_15 = t_r25_c15_12 >> 4;

  assign t_r25_c16_0 = p_24_16 << 1;
  assign t_r25_c16_1 = p_25_15 << 1;
  assign t_r25_c16_2 = p_25_16 << 2;
  assign t_r25_c16_3 = p_25_17 << 1;
  assign t_r25_c16_4 = p_26_16 << 1;
  assign t_r25_c16_5 = t_r25_c16_0 + p_24_15;
  assign t_r25_c16_6 = t_r25_c16_1 + p_24_17;
  assign t_r25_c16_7 = t_r25_c16_2 + t_r25_c16_3;
  assign t_r25_c16_8 = t_r25_c16_4 + p_26_15;
  assign t_r25_c16_9 = t_r25_c16_5 + t_r25_c16_6;
  assign t_r25_c16_10 = t_r25_c16_7 + t_r25_c16_8;
  assign t_r25_c16_11 = t_r25_c16_9 + t_r25_c16_10;
  assign t_r25_c16_12 = t_r25_c16_11 + p_26_17;
  assign out_25_16 = t_r25_c16_12 >> 4;

  assign t_r25_c17_0 = p_24_17 << 1;
  assign t_r25_c17_1 = p_25_16 << 1;
  assign t_r25_c17_2 = p_25_17 << 2;
  assign t_r25_c17_3 = p_25_18 << 1;
  assign t_r25_c17_4 = p_26_17 << 1;
  assign t_r25_c17_5 = t_r25_c17_0 + p_24_16;
  assign t_r25_c17_6 = t_r25_c17_1 + p_24_18;
  assign t_r25_c17_7 = t_r25_c17_2 + t_r25_c17_3;
  assign t_r25_c17_8 = t_r25_c17_4 + p_26_16;
  assign t_r25_c17_9 = t_r25_c17_5 + t_r25_c17_6;
  assign t_r25_c17_10 = t_r25_c17_7 + t_r25_c17_8;
  assign t_r25_c17_11 = t_r25_c17_9 + t_r25_c17_10;
  assign t_r25_c17_12 = t_r25_c17_11 + p_26_18;
  assign out_25_17 = t_r25_c17_12 >> 4;

  assign t_r25_c18_0 = p_24_18 << 1;
  assign t_r25_c18_1 = p_25_17 << 1;
  assign t_r25_c18_2 = p_25_18 << 2;
  assign t_r25_c18_3 = p_25_19 << 1;
  assign t_r25_c18_4 = p_26_18 << 1;
  assign t_r25_c18_5 = t_r25_c18_0 + p_24_17;
  assign t_r25_c18_6 = t_r25_c18_1 + p_24_19;
  assign t_r25_c18_7 = t_r25_c18_2 + t_r25_c18_3;
  assign t_r25_c18_8 = t_r25_c18_4 + p_26_17;
  assign t_r25_c18_9 = t_r25_c18_5 + t_r25_c18_6;
  assign t_r25_c18_10 = t_r25_c18_7 + t_r25_c18_8;
  assign t_r25_c18_11 = t_r25_c18_9 + t_r25_c18_10;
  assign t_r25_c18_12 = t_r25_c18_11 + p_26_19;
  assign out_25_18 = t_r25_c18_12 >> 4;

  assign t_r25_c19_0 = p_24_19 << 1;
  assign t_r25_c19_1 = p_25_18 << 1;
  assign t_r25_c19_2 = p_25_19 << 2;
  assign t_r25_c19_3 = p_25_20 << 1;
  assign t_r25_c19_4 = p_26_19 << 1;
  assign t_r25_c19_5 = t_r25_c19_0 + p_24_18;
  assign t_r25_c19_6 = t_r25_c19_1 + p_24_20;
  assign t_r25_c19_7 = t_r25_c19_2 + t_r25_c19_3;
  assign t_r25_c19_8 = t_r25_c19_4 + p_26_18;
  assign t_r25_c19_9 = t_r25_c19_5 + t_r25_c19_6;
  assign t_r25_c19_10 = t_r25_c19_7 + t_r25_c19_8;
  assign t_r25_c19_11 = t_r25_c19_9 + t_r25_c19_10;
  assign t_r25_c19_12 = t_r25_c19_11 + p_26_20;
  assign out_25_19 = t_r25_c19_12 >> 4;

  assign t_r25_c20_0 = p_24_20 << 1;
  assign t_r25_c20_1 = p_25_19 << 1;
  assign t_r25_c20_2 = p_25_20 << 2;
  assign t_r25_c20_3 = p_25_21 << 1;
  assign t_r25_c20_4 = p_26_20 << 1;
  assign t_r25_c20_5 = t_r25_c20_0 + p_24_19;
  assign t_r25_c20_6 = t_r25_c20_1 + p_24_21;
  assign t_r25_c20_7 = t_r25_c20_2 + t_r25_c20_3;
  assign t_r25_c20_8 = t_r25_c20_4 + p_26_19;
  assign t_r25_c20_9 = t_r25_c20_5 + t_r25_c20_6;
  assign t_r25_c20_10 = t_r25_c20_7 + t_r25_c20_8;
  assign t_r25_c20_11 = t_r25_c20_9 + t_r25_c20_10;
  assign t_r25_c20_12 = t_r25_c20_11 + p_26_21;
  assign out_25_20 = t_r25_c20_12 >> 4;

  assign t_r25_c21_0 = p_24_21 << 1;
  assign t_r25_c21_1 = p_25_20 << 1;
  assign t_r25_c21_2 = p_25_21 << 2;
  assign t_r25_c21_3 = p_25_22 << 1;
  assign t_r25_c21_4 = p_26_21 << 1;
  assign t_r25_c21_5 = t_r25_c21_0 + p_24_20;
  assign t_r25_c21_6 = t_r25_c21_1 + p_24_22;
  assign t_r25_c21_7 = t_r25_c21_2 + t_r25_c21_3;
  assign t_r25_c21_8 = t_r25_c21_4 + p_26_20;
  assign t_r25_c21_9 = t_r25_c21_5 + t_r25_c21_6;
  assign t_r25_c21_10 = t_r25_c21_7 + t_r25_c21_8;
  assign t_r25_c21_11 = t_r25_c21_9 + t_r25_c21_10;
  assign t_r25_c21_12 = t_r25_c21_11 + p_26_22;
  assign out_25_21 = t_r25_c21_12 >> 4;

  assign t_r25_c22_0 = p_24_22 << 1;
  assign t_r25_c22_1 = p_25_21 << 1;
  assign t_r25_c22_2 = p_25_22 << 2;
  assign t_r25_c22_3 = p_25_23 << 1;
  assign t_r25_c22_4 = p_26_22 << 1;
  assign t_r25_c22_5 = t_r25_c22_0 + p_24_21;
  assign t_r25_c22_6 = t_r25_c22_1 + p_24_23;
  assign t_r25_c22_7 = t_r25_c22_2 + t_r25_c22_3;
  assign t_r25_c22_8 = t_r25_c22_4 + p_26_21;
  assign t_r25_c22_9 = t_r25_c22_5 + t_r25_c22_6;
  assign t_r25_c22_10 = t_r25_c22_7 + t_r25_c22_8;
  assign t_r25_c22_11 = t_r25_c22_9 + t_r25_c22_10;
  assign t_r25_c22_12 = t_r25_c22_11 + p_26_23;
  assign out_25_22 = t_r25_c22_12 >> 4;

  assign t_r25_c23_0 = p_24_23 << 1;
  assign t_r25_c23_1 = p_25_22 << 1;
  assign t_r25_c23_2 = p_25_23 << 2;
  assign t_r25_c23_3 = p_25_24 << 1;
  assign t_r25_c23_4 = p_26_23 << 1;
  assign t_r25_c23_5 = t_r25_c23_0 + p_24_22;
  assign t_r25_c23_6 = t_r25_c23_1 + p_24_24;
  assign t_r25_c23_7 = t_r25_c23_2 + t_r25_c23_3;
  assign t_r25_c23_8 = t_r25_c23_4 + p_26_22;
  assign t_r25_c23_9 = t_r25_c23_5 + t_r25_c23_6;
  assign t_r25_c23_10 = t_r25_c23_7 + t_r25_c23_8;
  assign t_r25_c23_11 = t_r25_c23_9 + t_r25_c23_10;
  assign t_r25_c23_12 = t_r25_c23_11 + p_26_24;
  assign out_25_23 = t_r25_c23_12 >> 4;

  assign t_r25_c24_0 = p_24_24 << 1;
  assign t_r25_c24_1 = p_25_23 << 1;
  assign t_r25_c24_2 = p_25_24 << 2;
  assign t_r25_c24_3 = p_25_25 << 1;
  assign t_r25_c24_4 = p_26_24 << 1;
  assign t_r25_c24_5 = t_r25_c24_0 + p_24_23;
  assign t_r25_c24_6 = t_r25_c24_1 + p_24_25;
  assign t_r25_c24_7 = t_r25_c24_2 + t_r25_c24_3;
  assign t_r25_c24_8 = t_r25_c24_4 + p_26_23;
  assign t_r25_c24_9 = t_r25_c24_5 + t_r25_c24_6;
  assign t_r25_c24_10 = t_r25_c24_7 + t_r25_c24_8;
  assign t_r25_c24_11 = t_r25_c24_9 + t_r25_c24_10;
  assign t_r25_c24_12 = t_r25_c24_11 + p_26_25;
  assign out_25_24 = t_r25_c24_12 >> 4;

  assign t_r25_c25_0 = p_24_25 << 1;
  assign t_r25_c25_1 = p_25_24 << 1;
  assign t_r25_c25_2 = p_25_25 << 2;
  assign t_r25_c25_3 = p_25_26 << 1;
  assign t_r25_c25_4 = p_26_25 << 1;
  assign t_r25_c25_5 = t_r25_c25_0 + p_24_24;
  assign t_r25_c25_6 = t_r25_c25_1 + p_24_26;
  assign t_r25_c25_7 = t_r25_c25_2 + t_r25_c25_3;
  assign t_r25_c25_8 = t_r25_c25_4 + p_26_24;
  assign t_r25_c25_9 = t_r25_c25_5 + t_r25_c25_6;
  assign t_r25_c25_10 = t_r25_c25_7 + t_r25_c25_8;
  assign t_r25_c25_11 = t_r25_c25_9 + t_r25_c25_10;
  assign t_r25_c25_12 = t_r25_c25_11 + p_26_26;
  assign out_25_25 = t_r25_c25_12 >> 4;

  assign t_r25_c26_0 = p_24_26 << 1;
  assign t_r25_c26_1 = p_25_25 << 1;
  assign t_r25_c26_2 = p_25_26 << 2;
  assign t_r25_c26_3 = p_25_27 << 1;
  assign t_r25_c26_4 = p_26_26 << 1;
  assign t_r25_c26_5 = t_r25_c26_0 + p_24_25;
  assign t_r25_c26_6 = t_r25_c26_1 + p_24_27;
  assign t_r25_c26_7 = t_r25_c26_2 + t_r25_c26_3;
  assign t_r25_c26_8 = t_r25_c26_4 + p_26_25;
  assign t_r25_c26_9 = t_r25_c26_5 + t_r25_c26_6;
  assign t_r25_c26_10 = t_r25_c26_7 + t_r25_c26_8;
  assign t_r25_c26_11 = t_r25_c26_9 + t_r25_c26_10;
  assign t_r25_c26_12 = t_r25_c26_11 + p_26_27;
  assign out_25_26 = t_r25_c26_12 >> 4;

  assign t_r25_c27_0 = p_24_27 << 1;
  assign t_r25_c27_1 = p_25_26 << 1;
  assign t_r25_c27_2 = p_25_27 << 2;
  assign t_r25_c27_3 = p_25_28 << 1;
  assign t_r25_c27_4 = p_26_27 << 1;
  assign t_r25_c27_5 = t_r25_c27_0 + p_24_26;
  assign t_r25_c27_6 = t_r25_c27_1 + p_24_28;
  assign t_r25_c27_7 = t_r25_c27_2 + t_r25_c27_3;
  assign t_r25_c27_8 = t_r25_c27_4 + p_26_26;
  assign t_r25_c27_9 = t_r25_c27_5 + t_r25_c27_6;
  assign t_r25_c27_10 = t_r25_c27_7 + t_r25_c27_8;
  assign t_r25_c27_11 = t_r25_c27_9 + t_r25_c27_10;
  assign t_r25_c27_12 = t_r25_c27_11 + p_26_28;
  assign out_25_27 = t_r25_c27_12 >> 4;

  assign t_r25_c28_0 = p_24_28 << 1;
  assign t_r25_c28_1 = p_25_27 << 1;
  assign t_r25_c28_2 = p_25_28 << 2;
  assign t_r25_c28_3 = p_25_29 << 1;
  assign t_r25_c28_4 = p_26_28 << 1;
  assign t_r25_c28_5 = t_r25_c28_0 + p_24_27;
  assign t_r25_c28_6 = t_r25_c28_1 + p_24_29;
  assign t_r25_c28_7 = t_r25_c28_2 + t_r25_c28_3;
  assign t_r25_c28_8 = t_r25_c28_4 + p_26_27;
  assign t_r25_c28_9 = t_r25_c28_5 + t_r25_c28_6;
  assign t_r25_c28_10 = t_r25_c28_7 + t_r25_c28_8;
  assign t_r25_c28_11 = t_r25_c28_9 + t_r25_c28_10;
  assign t_r25_c28_12 = t_r25_c28_11 + p_26_29;
  assign out_25_28 = t_r25_c28_12 >> 4;

  assign t_r25_c29_0 = p_24_29 << 1;
  assign t_r25_c29_1 = p_25_28 << 1;
  assign t_r25_c29_2 = p_25_29 << 2;
  assign t_r25_c29_3 = p_25_30 << 1;
  assign t_r25_c29_4 = p_26_29 << 1;
  assign t_r25_c29_5 = t_r25_c29_0 + p_24_28;
  assign t_r25_c29_6 = t_r25_c29_1 + p_24_30;
  assign t_r25_c29_7 = t_r25_c29_2 + t_r25_c29_3;
  assign t_r25_c29_8 = t_r25_c29_4 + p_26_28;
  assign t_r25_c29_9 = t_r25_c29_5 + t_r25_c29_6;
  assign t_r25_c29_10 = t_r25_c29_7 + t_r25_c29_8;
  assign t_r25_c29_11 = t_r25_c29_9 + t_r25_c29_10;
  assign t_r25_c29_12 = t_r25_c29_11 + p_26_30;
  assign out_25_29 = t_r25_c29_12 >> 4;

  assign t_r25_c30_0 = p_24_30 << 1;
  assign t_r25_c30_1 = p_25_29 << 1;
  assign t_r25_c30_2 = p_25_30 << 2;
  assign t_r25_c30_3 = p_25_31 << 1;
  assign t_r25_c30_4 = p_26_30 << 1;
  assign t_r25_c30_5 = t_r25_c30_0 + p_24_29;
  assign t_r25_c30_6 = t_r25_c30_1 + p_24_31;
  assign t_r25_c30_7 = t_r25_c30_2 + t_r25_c30_3;
  assign t_r25_c30_8 = t_r25_c30_4 + p_26_29;
  assign t_r25_c30_9 = t_r25_c30_5 + t_r25_c30_6;
  assign t_r25_c30_10 = t_r25_c30_7 + t_r25_c30_8;
  assign t_r25_c30_11 = t_r25_c30_9 + t_r25_c30_10;
  assign t_r25_c30_12 = t_r25_c30_11 + p_26_31;
  assign out_25_30 = t_r25_c30_12 >> 4;

  assign t_r25_c31_0 = p_24_31 << 1;
  assign t_r25_c31_1 = p_25_30 << 1;
  assign t_r25_c31_2 = p_25_31 << 2;
  assign t_r25_c31_3 = p_25_32 << 1;
  assign t_r25_c31_4 = p_26_31 << 1;
  assign t_r25_c31_5 = t_r25_c31_0 + p_24_30;
  assign t_r25_c31_6 = t_r25_c31_1 + p_24_32;
  assign t_r25_c31_7 = t_r25_c31_2 + t_r25_c31_3;
  assign t_r25_c31_8 = t_r25_c31_4 + p_26_30;
  assign t_r25_c31_9 = t_r25_c31_5 + t_r25_c31_6;
  assign t_r25_c31_10 = t_r25_c31_7 + t_r25_c31_8;
  assign t_r25_c31_11 = t_r25_c31_9 + t_r25_c31_10;
  assign t_r25_c31_12 = t_r25_c31_11 + p_26_32;
  assign out_25_31 = t_r25_c31_12 >> 4;

  assign t_r25_c32_0 = p_24_32 << 1;
  assign t_r25_c32_1 = p_25_31 << 1;
  assign t_r25_c32_2 = p_25_32 << 2;
  assign t_r25_c32_3 = p_25_33 << 1;
  assign t_r25_c32_4 = p_26_32 << 1;
  assign t_r25_c32_5 = t_r25_c32_0 + p_24_31;
  assign t_r25_c32_6 = t_r25_c32_1 + p_24_33;
  assign t_r25_c32_7 = t_r25_c32_2 + t_r25_c32_3;
  assign t_r25_c32_8 = t_r25_c32_4 + p_26_31;
  assign t_r25_c32_9 = t_r25_c32_5 + t_r25_c32_6;
  assign t_r25_c32_10 = t_r25_c32_7 + t_r25_c32_8;
  assign t_r25_c32_11 = t_r25_c32_9 + t_r25_c32_10;
  assign t_r25_c32_12 = t_r25_c32_11 + p_26_33;
  assign out_25_32 = t_r25_c32_12 >> 4;

  assign t_r25_c33_0 = p_24_33 << 1;
  assign t_r25_c33_1 = p_25_32 << 1;
  assign t_r25_c33_2 = p_25_33 << 2;
  assign t_r25_c33_3 = p_25_34 << 1;
  assign t_r25_c33_4 = p_26_33 << 1;
  assign t_r25_c33_5 = t_r25_c33_0 + p_24_32;
  assign t_r25_c33_6 = t_r25_c33_1 + p_24_34;
  assign t_r25_c33_7 = t_r25_c33_2 + t_r25_c33_3;
  assign t_r25_c33_8 = t_r25_c33_4 + p_26_32;
  assign t_r25_c33_9 = t_r25_c33_5 + t_r25_c33_6;
  assign t_r25_c33_10 = t_r25_c33_7 + t_r25_c33_8;
  assign t_r25_c33_11 = t_r25_c33_9 + t_r25_c33_10;
  assign t_r25_c33_12 = t_r25_c33_11 + p_26_34;
  assign out_25_33 = t_r25_c33_12 >> 4;

  assign t_r25_c34_0 = p_24_34 << 1;
  assign t_r25_c34_1 = p_25_33 << 1;
  assign t_r25_c34_2 = p_25_34 << 2;
  assign t_r25_c34_3 = p_25_35 << 1;
  assign t_r25_c34_4 = p_26_34 << 1;
  assign t_r25_c34_5 = t_r25_c34_0 + p_24_33;
  assign t_r25_c34_6 = t_r25_c34_1 + p_24_35;
  assign t_r25_c34_7 = t_r25_c34_2 + t_r25_c34_3;
  assign t_r25_c34_8 = t_r25_c34_4 + p_26_33;
  assign t_r25_c34_9 = t_r25_c34_5 + t_r25_c34_6;
  assign t_r25_c34_10 = t_r25_c34_7 + t_r25_c34_8;
  assign t_r25_c34_11 = t_r25_c34_9 + t_r25_c34_10;
  assign t_r25_c34_12 = t_r25_c34_11 + p_26_35;
  assign out_25_34 = t_r25_c34_12 >> 4;

  assign t_r25_c35_0 = p_24_35 << 1;
  assign t_r25_c35_1 = p_25_34 << 1;
  assign t_r25_c35_2 = p_25_35 << 2;
  assign t_r25_c35_3 = p_25_36 << 1;
  assign t_r25_c35_4 = p_26_35 << 1;
  assign t_r25_c35_5 = t_r25_c35_0 + p_24_34;
  assign t_r25_c35_6 = t_r25_c35_1 + p_24_36;
  assign t_r25_c35_7 = t_r25_c35_2 + t_r25_c35_3;
  assign t_r25_c35_8 = t_r25_c35_4 + p_26_34;
  assign t_r25_c35_9 = t_r25_c35_5 + t_r25_c35_6;
  assign t_r25_c35_10 = t_r25_c35_7 + t_r25_c35_8;
  assign t_r25_c35_11 = t_r25_c35_9 + t_r25_c35_10;
  assign t_r25_c35_12 = t_r25_c35_11 + p_26_36;
  assign out_25_35 = t_r25_c35_12 >> 4;

  assign t_r25_c36_0 = p_24_36 << 1;
  assign t_r25_c36_1 = p_25_35 << 1;
  assign t_r25_c36_2 = p_25_36 << 2;
  assign t_r25_c36_3 = p_25_37 << 1;
  assign t_r25_c36_4 = p_26_36 << 1;
  assign t_r25_c36_5 = t_r25_c36_0 + p_24_35;
  assign t_r25_c36_6 = t_r25_c36_1 + p_24_37;
  assign t_r25_c36_7 = t_r25_c36_2 + t_r25_c36_3;
  assign t_r25_c36_8 = t_r25_c36_4 + p_26_35;
  assign t_r25_c36_9 = t_r25_c36_5 + t_r25_c36_6;
  assign t_r25_c36_10 = t_r25_c36_7 + t_r25_c36_8;
  assign t_r25_c36_11 = t_r25_c36_9 + t_r25_c36_10;
  assign t_r25_c36_12 = t_r25_c36_11 + p_26_37;
  assign out_25_36 = t_r25_c36_12 >> 4;

  assign t_r25_c37_0 = p_24_37 << 1;
  assign t_r25_c37_1 = p_25_36 << 1;
  assign t_r25_c37_2 = p_25_37 << 2;
  assign t_r25_c37_3 = p_25_38 << 1;
  assign t_r25_c37_4 = p_26_37 << 1;
  assign t_r25_c37_5 = t_r25_c37_0 + p_24_36;
  assign t_r25_c37_6 = t_r25_c37_1 + p_24_38;
  assign t_r25_c37_7 = t_r25_c37_2 + t_r25_c37_3;
  assign t_r25_c37_8 = t_r25_c37_4 + p_26_36;
  assign t_r25_c37_9 = t_r25_c37_5 + t_r25_c37_6;
  assign t_r25_c37_10 = t_r25_c37_7 + t_r25_c37_8;
  assign t_r25_c37_11 = t_r25_c37_9 + t_r25_c37_10;
  assign t_r25_c37_12 = t_r25_c37_11 + p_26_38;
  assign out_25_37 = t_r25_c37_12 >> 4;

  assign t_r25_c38_0 = p_24_38 << 1;
  assign t_r25_c38_1 = p_25_37 << 1;
  assign t_r25_c38_2 = p_25_38 << 2;
  assign t_r25_c38_3 = p_25_39 << 1;
  assign t_r25_c38_4 = p_26_38 << 1;
  assign t_r25_c38_5 = t_r25_c38_0 + p_24_37;
  assign t_r25_c38_6 = t_r25_c38_1 + p_24_39;
  assign t_r25_c38_7 = t_r25_c38_2 + t_r25_c38_3;
  assign t_r25_c38_8 = t_r25_c38_4 + p_26_37;
  assign t_r25_c38_9 = t_r25_c38_5 + t_r25_c38_6;
  assign t_r25_c38_10 = t_r25_c38_7 + t_r25_c38_8;
  assign t_r25_c38_11 = t_r25_c38_9 + t_r25_c38_10;
  assign t_r25_c38_12 = t_r25_c38_11 + p_26_39;
  assign out_25_38 = t_r25_c38_12 >> 4;

  assign t_r25_c39_0 = p_24_39 << 1;
  assign t_r25_c39_1 = p_25_38 << 1;
  assign t_r25_c39_2 = p_25_39 << 2;
  assign t_r25_c39_3 = p_25_40 << 1;
  assign t_r25_c39_4 = p_26_39 << 1;
  assign t_r25_c39_5 = t_r25_c39_0 + p_24_38;
  assign t_r25_c39_6 = t_r25_c39_1 + p_24_40;
  assign t_r25_c39_7 = t_r25_c39_2 + t_r25_c39_3;
  assign t_r25_c39_8 = t_r25_c39_4 + p_26_38;
  assign t_r25_c39_9 = t_r25_c39_5 + t_r25_c39_6;
  assign t_r25_c39_10 = t_r25_c39_7 + t_r25_c39_8;
  assign t_r25_c39_11 = t_r25_c39_9 + t_r25_c39_10;
  assign t_r25_c39_12 = t_r25_c39_11 + p_26_40;
  assign out_25_39 = t_r25_c39_12 >> 4;

  assign t_r25_c40_0 = p_24_40 << 1;
  assign t_r25_c40_1 = p_25_39 << 1;
  assign t_r25_c40_2 = p_25_40 << 2;
  assign t_r25_c40_3 = p_25_41 << 1;
  assign t_r25_c40_4 = p_26_40 << 1;
  assign t_r25_c40_5 = t_r25_c40_0 + p_24_39;
  assign t_r25_c40_6 = t_r25_c40_1 + p_24_41;
  assign t_r25_c40_7 = t_r25_c40_2 + t_r25_c40_3;
  assign t_r25_c40_8 = t_r25_c40_4 + p_26_39;
  assign t_r25_c40_9 = t_r25_c40_5 + t_r25_c40_6;
  assign t_r25_c40_10 = t_r25_c40_7 + t_r25_c40_8;
  assign t_r25_c40_11 = t_r25_c40_9 + t_r25_c40_10;
  assign t_r25_c40_12 = t_r25_c40_11 + p_26_41;
  assign out_25_40 = t_r25_c40_12 >> 4;

  assign t_r25_c41_0 = p_24_41 << 1;
  assign t_r25_c41_1 = p_25_40 << 1;
  assign t_r25_c41_2 = p_25_41 << 2;
  assign t_r25_c41_3 = p_25_42 << 1;
  assign t_r25_c41_4 = p_26_41 << 1;
  assign t_r25_c41_5 = t_r25_c41_0 + p_24_40;
  assign t_r25_c41_6 = t_r25_c41_1 + p_24_42;
  assign t_r25_c41_7 = t_r25_c41_2 + t_r25_c41_3;
  assign t_r25_c41_8 = t_r25_c41_4 + p_26_40;
  assign t_r25_c41_9 = t_r25_c41_5 + t_r25_c41_6;
  assign t_r25_c41_10 = t_r25_c41_7 + t_r25_c41_8;
  assign t_r25_c41_11 = t_r25_c41_9 + t_r25_c41_10;
  assign t_r25_c41_12 = t_r25_c41_11 + p_26_42;
  assign out_25_41 = t_r25_c41_12 >> 4;

  assign t_r25_c42_0 = p_24_42 << 1;
  assign t_r25_c42_1 = p_25_41 << 1;
  assign t_r25_c42_2 = p_25_42 << 2;
  assign t_r25_c42_3 = p_25_43 << 1;
  assign t_r25_c42_4 = p_26_42 << 1;
  assign t_r25_c42_5 = t_r25_c42_0 + p_24_41;
  assign t_r25_c42_6 = t_r25_c42_1 + p_24_43;
  assign t_r25_c42_7 = t_r25_c42_2 + t_r25_c42_3;
  assign t_r25_c42_8 = t_r25_c42_4 + p_26_41;
  assign t_r25_c42_9 = t_r25_c42_5 + t_r25_c42_6;
  assign t_r25_c42_10 = t_r25_c42_7 + t_r25_c42_8;
  assign t_r25_c42_11 = t_r25_c42_9 + t_r25_c42_10;
  assign t_r25_c42_12 = t_r25_c42_11 + p_26_43;
  assign out_25_42 = t_r25_c42_12 >> 4;

  assign t_r25_c43_0 = p_24_43 << 1;
  assign t_r25_c43_1 = p_25_42 << 1;
  assign t_r25_c43_2 = p_25_43 << 2;
  assign t_r25_c43_3 = p_25_44 << 1;
  assign t_r25_c43_4 = p_26_43 << 1;
  assign t_r25_c43_5 = t_r25_c43_0 + p_24_42;
  assign t_r25_c43_6 = t_r25_c43_1 + p_24_44;
  assign t_r25_c43_7 = t_r25_c43_2 + t_r25_c43_3;
  assign t_r25_c43_8 = t_r25_c43_4 + p_26_42;
  assign t_r25_c43_9 = t_r25_c43_5 + t_r25_c43_6;
  assign t_r25_c43_10 = t_r25_c43_7 + t_r25_c43_8;
  assign t_r25_c43_11 = t_r25_c43_9 + t_r25_c43_10;
  assign t_r25_c43_12 = t_r25_c43_11 + p_26_44;
  assign out_25_43 = t_r25_c43_12 >> 4;

  assign t_r25_c44_0 = p_24_44 << 1;
  assign t_r25_c44_1 = p_25_43 << 1;
  assign t_r25_c44_2 = p_25_44 << 2;
  assign t_r25_c44_3 = p_25_45 << 1;
  assign t_r25_c44_4 = p_26_44 << 1;
  assign t_r25_c44_5 = t_r25_c44_0 + p_24_43;
  assign t_r25_c44_6 = t_r25_c44_1 + p_24_45;
  assign t_r25_c44_7 = t_r25_c44_2 + t_r25_c44_3;
  assign t_r25_c44_8 = t_r25_c44_4 + p_26_43;
  assign t_r25_c44_9 = t_r25_c44_5 + t_r25_c44_6;
  assign t_r25_c44_10 = t_r25_c44_7 + t_r25_c44_8;
  assign t_r25_c44_11 = t_r25_c44_9 + t_r25_c44_10;
  assign t_r25_c44_12 = t_r25_c44_11 + p_26_45;
  assign out_25_44 = t_r25_c44_12 >> 4;

  assign t_r25_c45_0 = p_24_45 << 1;
  assign t_r25_c45_1 = p_25_44 << 1;
  assign t_r25_c45_2 = p_25_45 << 2;
  assign t_r25_c45_3 = p_25_46 << 1;
  assign t_r25_c45_4 = p_26_45 << 1;
  assign t_r25_c45_5 = t_r25_c45_0 + p_24_44;
  assign t_r25_c45_6 = t_r25_c45_1 + p_24_46;
  assign t_r25_c45_7 = t_r25_c45_2 + t_r25_c45_3;
  assign t_r25_c45_8 = t_r25_c45_4 + p_26_44;
  assign t_r25_c45_9 = t_r25_c45_5 + t_r25_c45_6;
  assign t_r25_c45_10 = t_r25_c45_7 + t_r25_c45_8;
  assign t_r25_c45_11 = t_r25_c45_9 + t_r25_c45_10;
  assign t_r25_c45_12 = t_r25_c45_11 + p_26_46;
  assign out_25_45 = t_r25_c45_12 >> 4;

  assign t_r25_c46_0 = p_24_46 << 1;
  assign t_r25_c46_1 = p_25_45 << 1;
  assign t_r25_c46_2 = p_25_46 << 2;
  assign t_r25_c46_3 = p_25_47 << 1;
  assign t_r25_c46_4 = p_26_46 << 1;
  assign t_r25_c46_5 = t_r25_c46_0 + p_24_45;
  assign t_r25_c46_6 = t_r25_c46_1 + p_24_47;
  assign t_r25_c46_7 = t_r25_c46_2 + t_r25_c46_3;
  assign t_r25_c46_8 = t_r25_c46_4 + p_26_45;
  assign t_r25_c46_9 = t_r25_c46_5 + t_r25_c46_6;
  assign t_r25_c46_10 = t_r25_c46_7 + t_r25_c46_8;
  assign t_r25_c46_11 = t_r25_c46_9 + t_r25_c46_10;
  assign t_r25_c46_12 = t_r25_c46_11 + p_26_47;
  assign out_25_46 = t_r25_c46_12 >> 4;

  assign t_r25_c47_0 = p_24_47 << 1;
  assign t_r25_c47_1 = p_25_46 << 1;
  assign t_r25_c47_2 = p_25_47 << 2;
  assign t_r25_c47_3 = p_25_48 << 1;
  assign t_r25_c47_4 = p_26_47 << 1;
  assign t_r25_c47_5 = t_r25_c47_0 + p_24_46;
  assign t_r25_c47_6 = t_r25_c47_1 + p_24_48;
  assign t_r25_c47_7 = t_r25_c47_2 + t_r25_c47_3;
  assign t_r25_c47_8 = t_r25_c47_4 + p_26_46;
  assign t_r25_c47_9 = t_r25_c47_5 + t_r25_c47_6;
  assign t_r25_c47_10 = t_r25_c47_7 + t_r25_c47_8;
  assign t_r25_c47_11 = t_r25_c47_9 + t_r25_c47_10;
  assign t_r25_c47_12 = t_r25_c47_11 + p_26_48;
  assign out_25_47 = t_r25_c47_12 >> 4;

  assign t_r25_c48_0 = p_24_48 << 1;
  assign t_r25_c48_1 = p_25_47 << 1;
  assign t_r25_c48_2 = p_25_48 << 2;
  assign t_r25_c48_3 = p_25_49 << 1;
  assign t_r25_c48_4 = p_26_48 << 1;
  assign t_r25_c48_5 = t_r25_c48_0 + p_24_47;
  assign t_r25_c48_6 = t_r25_c48_1 + p_24_49;
  assign t_r25_c48_7 = t_r25_c48_2 + t_r25_c48_3;
  assign t_r25_c48_8 = t_r25_c48_4 + p_26_47;
  assign t_r25_c48_9 = t_r25_c48_5 + t_r25_c48_6;
  assign t_r25_c48_10 = t_r25_c48_7 + t_r25_c48_8;
  assign t_r25_c48_11 = t_r25_c48_9 + t_r25_c48_10;
  assign t_r25_c48_12 = t_r25_c48_11 + p_26_49;
  assign out_25_48 = t_r25_c48_12 >> 4;

  assign t_r25_c49_0 = p_24_49 << 1;
  assign t_r25_c49_1 = p_25_48 << 1;
  assign t_r25_c49_2 = p_25_49 << 2;
  assign t_r25_c49_3 = p_25_50 << 1;
  assign t_r25_c49_4 = p_26_49 << 1;
  assign t_r25_c49_5 = t_r25_c49_0 + p_24_48;
  assign t_r25_c49_6 = t_r25_c49_1 + p_24_50;
  assign t_r25_c49_7 = t_r25_c49_2 + t_r25_c49_3;
  assign t_r25_c49_8 = t_r25_c49_4 + p_26_48;
  assign t_r25_c49_9 = t_r25_c49_5 + t_r25_c49_6;
  assign t_r25_c49_10 = t_r25_c49_7 + t_r25_c49_8;
  assign t_r25_c49_11 = t_r25_c49_9 + t_r25_c49_10;
  assign t_r25_c49_12 = t_r25_c49_11 + p_26_50;
  assign out_25_49 = t_r25_c49_12 >> 4;

  assign t_r25_c50_0 = p_24_50 << 1;
  assign t_r25_c50_1 = p_25_49 << 1;
  assign t_r25_c50_2 = p_25_50 << 2;
  assign t_r25_c50_3 = p_25_51 << 1;
  assign t_r25_c50_4 = p_26_50 << 1;
  assign t_r25_c50_5 = t_r25_c50_0 + p_24_49;
  assign t_r25_c50_6 = t_r25_c50_1 + p_24_51;
  assign t_r25_c50_7 = t_r25_c50_2 + t_r25_c50_3;
  assign t_r25_c50_8 = t_r25_c50_4 + p_26_49;
  assign t_r25_c50_9 = t_r25_c50_5 + t_r25_c50_6;
  assign t_r25_c50_10 = t_r25_c50_7 + t_r25_c50_8;
  assign t_r25_c50_11 = t_r25_c50_9 + t_r25_c50_10;
  assign t_r25_c50_12 = t_r25_c50_11 + p_26_51;
  assign out_25_50 = t_r25_c50_12 >> 4;

  assign t_r25_c51_0 = p_24_51 << 1;
  assign t_r25_c51_1 = p_25_50 << 1;
  assign t_r25_c51_2 = p_25_51 << 2;
  assign t_r25_c51_3 = p_25_52 << 1;
  assign t_r25_c51_4 = p_26_51 << 1;
  assign t_r25_c51_5 = t_r25_c51_0 + p_24_50;
  assign t_r25_c51_6 = t_r25_c51_1 + p_24_52;
  assign t_r25_c51_7 = t_r25_c51_2 + t_r25_c51_3;
  assign t_r25_c51_8 = t_r25_c51_4 + p_26_50;
  assign t_r25_c51_9 = t_r25_c51_5 + t_r25_c51_6;
  assign t_r25_c51_10 = t_r25_c51_7 + t_r25_c51_8;
  assign t_r25_c51_11 = t_r25_c51_9 + t_r25_c51_10;
  assign t_r25_c51_12 = t_r25_c51_11 + p_26_52;
  assign out_25_51 = t_r25_c51_12 >> 4;

  assign t_r25_c52_0 = p_24_52 << 1;
  assign t_r25_c52_1 = p_25_51 << 1;
  assign t_r25_c52_2 = p_25_52 << 2;
  assign t_r25_c52_3 = p_25_53 << 1;
  assign t_r25_c52_4 = p_26_52 << 1;
  assign t_r25_c52_5 = t_r25_c52_0 + p_24_51;
  assign t_r25_c52_6 = t_r25_c52_1 + p_24_53;
  assign t_r25_c52_7 = t_r25_c52_2 + t_r25_c52_3;
  assign t_r25_c52_8 = t_r25_c52_4 + p_26_51;
  assign t_r25_c52_9 = t_r25_c52_5 + t_r25_c52_6;
  assign t_r25_c52_10 = t_r25_c52_7 + t_r25_c52_8;
  assign t_r25_c52_11 = t_r25_c52_9 + t_r25_c52_10;
  assign t_r25_c52_12 = t_r25_c52_11 + p_26_53;
  assign out_25_52 = t_r25_c52_12 >> 4;

  assign t_r25_c53_0 = p_24_53 << 1;
  assign t_r25_c53_1 = p_25_52 << 1;
  assign t_r25_c53_2 = p_25_53 << 2;
  assign t_r25_c53_3 = p_25_54 << 1;
  assign t_r25_c53_4 = p_26_53 << 1;
  assign t_r25_c53_5 = t_r25_c53_0 + p_24_52;
  assign t_r25_c53_6 = t_r25_c53_1 + p_24_54;
  assign t_r25_c53_7 = t_r25_c53_2 + t_r25_c53_3;
  assign t_r25_c53_8 = t_r25_c53_4 + p_26_52;
  assign t_r25_c53_9 = t_r25_c53_5 + t_r25_c53_6;
  assign t_r25_c53_10 = t_r25_c53_7 + t_r25_c53_8;
  assign t_r25_c53_11 = t_r25_c53_9 + t_r25_c53_10;
  assign t_r25_c53_12 = t_r25_c53_11 + p_26_54;
  assign out_25_53 = t_r25_c53_12 >> 4;

  assign t_r25_c54_0 = p_24_54 << 1;
  assign t_r25_c54_1 = p_25_53 << 1;
  assign t_r25_c54_2 = p_25_54 << 2;
  assign t_r25_c54_3 = p_25_55 << 1;
  assign t_r25_c54_4 = p_26_54 << 1;
  assign t_r25_c54_5 = t_r25_c54_0 + p_24_53;
  assign t_r25_c54_6 = t_r25_c54_1 + p_24_55;
  assign t_r25_c54_7 = t_r25_c54_2 + t_r25_c54_3;
  assign t_r25_c54_8 = t_r25_c54_4 + p_26_53;
  assign t_r25_c54_9 = t_r25_c54_5 + t_r25_c54_6;
  assign t_r25_c54_10 = t_r25_c54_7 + t_r25_c54_8;
  assign t_r25_c54_11 = t_r25_c54_9 + t_r25_c54_10;
  assign t_r25_c54_12 = t_r25_c54_11 + p_26_55;
  assign out_25_54 = t_r25_c54_12 >> 4;

  assign t_r25_c55_0 = p_24_55 << 1;
  assign t_r25_c55_1 = p_25_54 << 1;
  assign t_r25_c55_2 = p_25_55 << 2;
  assign t_r25_c55_3 = p_25_56 << 1;
  assign t_r25_c55_4 = p_26_55 << 1;
  assign t_r25_c55_5 = t_r25_c55_0 + p_24_54;
  assign t_r25_c55_6 = t_r25_c55_1 + p_24_56;
  assign t_r25_c55_7 = t_r25_c55_2 + t_r25_c55_3;
  assign t_r25_c55_8 = t_r25_c55_4 + p_26_54;
  assign t_r25_c55_9 = t_r25_c55_5 + t_r25_c55_6;
  assign t_r25_c55_10 = t_r25_c55_7 + t_r25_c55_8;
  assign t_r25_c55_11 = t_r25_c55_9 + t_r25_c55_10;
  assign t_r25_c55_12 = t_r25_c55_11 + p_26_56;
  assign out_25_55 = t_r25_c55_12 >> 4;

  assign t_r25_c56_0 = p_24_56 << 1;
  assign t_r25_c56_1 = p_25_55 << 1;
  assign t_r25_c56_2 = p_25_56 << 2;
  assign t_r25_c56_3 = p_25_57 << 1;
  assign t_r25_c56_4 = p_26_56 << 1;
  assign t_r25_c56_5 = t_r25_c56_0 + p_24_55;
  assign t_r25_c56_6 = t_r25_c56_1 + p_24_57;
  assign t_r25_c56_7 = t_r25_c56_2 + t_r25_c56_3;
  assign t_r25_c56_8 = t_r25_c56_4 + p_26_55;
  assign t_r25_c56_9 = t_r25_c56_5 + t_r25_c56_6;
  assign t_r25_c56_10 = t_r25_c56_7 + t_r25_c56_8;
  assign t_r25_c56_11 = t_r25_c56_9 + t_r25_c56_10;
  assign t_r25_c56_12 = t_r25_c56_11 + p_26_57;
  assign out_25_56 = t_r25_c56_12 >> 4;

  assign t_r25_c57_0 = p_24_57 << 1;
  assign t_r25_c57_1 = p_25_56 << 1;
  assign t_r25_c57_2 = p_25_57 << 2;
  assign t_r25_c57_3 = p_25_58 << 1;
  assign t_r25_c57_4 = p_26_57 << 1;
  assign t_r25_c57_5 = t_r25_c57_0 + p_24_56;
  assign t_r25_c57_6 = t_r25_c57_1 + p_24_58;
  assign t_r25_c57_7 = t_r25_c57_2 + t_r25_c57_3;
  assign t_r25_c57_8 = t_r25_c57_4 + p_26_56;
  assign t_r25_c57_9 = t_r25_c57_5 + t_r25_c57_6;
  assign t_r25_c57_10 = t_r25_c57_7 + t_r25_c57_8;
  assign t_r25_c57_11 = t_r25_c57_9 + t_r25_c57_10;
  assign t_r25_c57_12 = t_r25_c57_11 + p_26_58;
  assign out_25_57 = t_r25_c57_12 >> 4;

  assign t_r25_c58_0 = p_24_58 << 1;
  assign t_r25_c58_1 = p_25_57 << 1;
  assign t_r25_c58_2 = p_25_58 << 2;
  assign t_r25_c58_3 = p_25_59 << 1;
  assign t_r25_c58_4 = p_26_58 << 1;
  assign t_r25_c58_5 = t_r25_c58_0 + p_24_57;
  assign t_r25_c58_6 = t_r25_c58_1 + p_24_59;
  assign t_r25_c58_7 = t_r25_c58_2 + t_r25_c58_3;
  assign t_r25_c58_8 = t_r25_c58_4 + p_26_57;
  assign t_r25_c58_9 = t_r25_c58_5 + t_r25_c58_6;
  assign t_r25_c58_10 = t_r25_c58_7 + t_r25_c58_8;
  assign t_r25_c58_11 = t_r25_c58_9 + t_r25_c58_10;
  assign t_r25_c58_12 = t_r25_c58_11 + p_26_59;
  assign out_25_58 = t_r25_c58_12 >> 4;

  assign t_r25_c59_0 = p_24_59 << 1;
  assign t_r25_c59_1 = p_25_58 << 1;
  assign t_r25_c59_2 = p_25_59 << 2;
  assign t_r25_c59_3 = p_25_60 << 1;
  assign t_r25_c59_4 = p_26_59 << 1;
  assign t_r25_c59_5 = t_r25_c59_0 + p_24_58;
  assign t_r25_c59_6 = t_r25_c59_1 + p_24_60;
  assign t_r25_c59_7 = t_r25_c59_2 + t_r25_c59_3;
  assign t_r25_c59_8 = t_r25_c59_4 + p_26_58;
  assign t_r25_c59_9 = t_r25_c59_5 + t_r25_c59_6;
  assign t_r25_c59_10 = t_r25_c59_7 + t_r25_c59_8;
  assign t_r25_c59_11 = t_r25_c59_9 + t_r25_c59_10;
  assign t_r25_c59_12 = t_r25_c59_11 + p_26_60;
  assign out_25_59 = t_r25_c59_12 >> 4;

  assign t_r25_c60_0 = p_24_60 << 1;
  assign t_r25_c60_1 = p_25_59 << 1;
  assign t_r25_c60_2 = p_25_60 << 2;
  assign t_r25_c60_3 = p_25_61 << 1;
  assign t_r25_c60_4 = p_26_60 << 1;
  assign t_r25_c60_5 = t_r25_c60_0 + p_24_59;
  assign t_r25_c60_6 = t_r25_c60_1 + p_24_61;
  assign t_r25_c60_7 = t_r25_c60_2 + t_r25_c60_3;
  assign t_r25_c60_8 = t_r25_c60_4 + p_26_59;
  assign t_r25_c60_9 = t_r25_c60_5 + t_r25_c60_6;
  assign t_r25_c60_10 = t_r25_c60_7 + t_r25_c60_8;
  assign t_r25_c60_11 = t_r25_c60_9 + t_r25_c60_10;
  assign t_r25_c60_12 = t_r25_c60_11 + p_26_61;
  assign out_25_60 = t_r25_c60_12 >> 4;

  assign t_r25_c61_0 = p_24_61 << 1;
  assign t_r25_c61_1 = p_25_60 << 1;
  assign t_r25_c61_2 = p_25_61 << 2;
  assign t_r25_c61_3 = p_25_62 << 1;
  assign t_r25_c61_4 = p_26_61 << 1;
  assign t_r25_c61_5 = t_r25_c61_0 + p_24_60;
  assign t_r25_c61_6 = t_r25_c61_1 + p_24_62;
  assign t_r25_c61_7 = t_r25_c61_2 + t_r25_c61_3;
  assign t_r25_c61_8 = t_r25_c61_4 + p_26_60;
  assign t_r25_c61_9 = t_r25_c61_5 + t_r25_c61_6;
  assign t_r25_c61_10 = t_r25_c61_7 + t_r25_c61_8;
  assign t_r25_c61_11 = t_r25_c61_9 + t_r25_c61_10;
  assign t_r25_c61_12 = t_r25_c61_11 + p_26_62;
  assign out_25_61 = t_r25_c61_12 >> 4;

  assign t_r25_c62_0 = p_24_62 << 1;
  assign t_r25_c62_1 = p_25_61 << 1;
  assign t_r25_c62_2 = p_25_62 << 2;
  assign t_r25_c62_3 = p_25_63 << 1;
  assign t_r25_c62_4 = p_26_62 << 1;
  assign t_r25_c62_5 = t_r25_c62_0 + p_24_61;
  assign t_r25_c62_6 = t_r25_c62_1 + p_24_63;
  assign t_r25_c62_7 = t_r25_c62_2 + t_r25_c62_3;
  assign t_r25_c62_8 = t_r25_c62_4 + p_26_61;
  assign t_r25_c62_9 = t_r25_c62_5 + t_r25_c62_6;
  assign t_r25_c62_10 = t_r25_c62_7 + t_r25_c62_8;
  assign t_r25_c62_11 = t_r25_c62_9 + t_r25_c62_10;
  assign t_r25_c62_12 = t_r25_c62_11 + p_26_63;
  assign out_25_62 = t_r25_c62_12 >> 4;

  assign t_r25_c63_0 = p_24_63 << 1;
  assign t_r25_c63_1 = p_25_62 << 1;
  assign t_r25_c63_2 = p_25_63 << 2;
  assign t_r25_c63_3 = p_25_64 << 1;
  assign t_r25_c63_4 = p_26_63 << 1;
  assign t_r25_c63_5 = t_r25_c63_0 + p_24_62;
  assign t_r25_c63_6 = t_r25_c63_1 + p_24_64;
  assign t_r25_c63_7 = t_r25_c63_2 + t_r25_c63_3;
  assign t_r25_c63_8 = t_r25_c63_4 + p_26_62;
  assign t_r25_c63_9 = t_r25_c63_5 + t_r25_c63_6;
  assign t_r25_c63_10 = t_r25_c63_7 + t_r25_c63_8;
  assign t_r25_c63_11 = t_r25_c63_9 + t_r25_c63_10;
  assign t_r25_c63_12 = t_r25_c63_11 + p_26_64;
  assign out_25_63 = t_r25_c63_12 >> 4;

  assign t_r25_c64_0 = p_24_64 << 1;
  assign t_r25_c64_1 = p_25_63 << 1;
  assign t_r25_c64_2 = p_25_64 << 2;
  assign t_r25_c64_3 = p_25_65 << 1;
  assign t_r25_c64_4 = p_26_64 << 1;
  assign t_r25_c64_5 = t_r25_c64_0 + p_24_63;
  assign t_r25_c64_6 = t_r25_c64_1 + p_24_65;
  assign t_r25_c64_7 = t_r25_c64_2 + t_r25_c64_3;
  assign t_r25_c64_8 = t_r25_c64_4 + p_26_63;
  assign t_r25_c64_9 = t_r25_c64_5 + t_r25_c64_6;
  assign t_r25_c64_10 = t_r25_c64_7 + t_r25_c64_8;
  assign t_r25_c64_11 = t_r25_c64_9 + t_r25_c64_10;
  assign t_r25_c64_12 = t_r25_c64_11 + p_26_65;
  assign out_25_64 = t_r25_c64_12 >> 4;

  assign t_r26_c1_0 = p_25_1 << 1;
  assign t_r26_c1_1 = p_26_0 << 1;
  assign t_r26_c1_2 = p_26_1 << 2;
  assign t_r26_c1_3 = p_26_2 << 1;
  assign t_r26_c1_4 = p_27_1 << 1;
  assign t_r26_c1_5 = t_r26_c1_0 + p_25_0;
  assign t_r26_c1_6 = t_r26_c1_1 + p_25_2;
  assign t_r26_c1_7 = t_r26_c1_2 + t_r26_c1_3;
  assign t_r26_c1_8 = t_r26_c1_4 + p_27_0;
  assign t_r26_c1_9 = t_r26_c1_5 + t_r26_c1_6;
  assign t_r26_c1_10 = t_r26_c1_7 + t_r26_c1_8;
  assign t_r26_c1_11 = t_r26_c1_9 + t_r26_c1_10;
  assign t_r26_c1_12 = t_r26_c1_11 + p_27_2;
  assign out_26_1 = t_r26_c1_12 >> 4;

  assign t_r26_c2_0 = p_25_2 << 1;
  assign t_r26_c2_1 = p_26_1 << 1;
  assign t_r26_c2_2 = p_26_2 << 2;
  assign t_r26_c2_3 = p_26_3 << 1;
  assign t_r26_c2_4 = p_27_2 << 1;
  assign t_r26_c2_5 = t_r26_c2_0 + p_25_1;
  assign t_r26_c2_6 = t_r26_c2_1 + p_25_3;
  assign t_r26_c2_7 = t_r26_c2_2 + t_r26_c2_3;
  assign t_r26_c2_8 = t_r26_c2_4 + p_27_1;
  assign t_r26_c2_9 = t_r26_c2_5 + t_r26_c2_6;
  assign t_r26_c2_10 = t_r26_c2_7 + t_r26_c2_8;
  assign t_r26_c2_11 = t_r26_c2_9 + t_r26_c2_10;
  assign t_r26_c2_12 = t_r26_c2_11 + p_27_3;
  assign out_26_2 = t_r26_c2_12 >> 4;

  assign t_r26_c3_0 = p_25_3 << 1;
  assign t_r26_c3_1 = p_26_2 << 1;
  assign t_r26_c3_2 = p_26_3 << 2;
  assign t_r26_c3_3 = p_26_4 << 1;
  assign t_r26_c3_4 = p_27_3 << 1;
  assign t_r26_c3_5 = t_r26_c3_0 + p_25_2;
  assign t_r26_c3_6 = t_r26_c3_1 + p_25_4;
  assign t_r26_c3_7 = t_r26_c3_2 + t_r26_c3_3;
  assign t_r26_c3_8 = t_r26_c3_4 + p_27_2;
  assign t_r26_c3_9 = t_r26_c3_5 + t_r26_c3_6;
  assign t_r26_c3_10 = t_r26_c3_7 + t_r26_c3_8;
  assign t_r26_c3_11 = t_r26_c3_9 + t_r26_c3_10;
  assign t_r26_c3_12 = t_r26_c3_11 + p_27_4;
  assign out_26_3 = t_r26_c3_12 >> 4;

  assign t_r26_c4_0 = p_25_4 << 1;
  assign t_r26_c4_1 = p_26_3 << 1;
  assign t_r26_c4_2 = p_26_4 << 2;
  assign t_r26_c4_3 = p_26_5 << 1;
  assign t_r26_c4_4 = p_27_4 << 1;
  assign t_r26_c4_5 = t_r26_c4_0 + p_25_3;
  assign t_r26_c4_6 = t_r26_c4_1 + p_25_5;
  assign t_r26_c4_7 = t_r26_c4_2 + t_r26_c4_3;
  assign t_r26_c4_8 = t_r26_c4_4 + p_27_3;
  assign t_r26_c4_9 = t_r26_c4_5 + t_r26_c4_6;
  assign t_r26_c4_10 = t_r26_c4_7 + t_r26_c4_8;
  assign t_r26_c4_11 = t_r26_c4_9 + t_r26_c4_10;
  assign t_r26_c4_12 = t_r26_c4_11 + p_27_5;
  assign out_26_4 = t_r26_c4_12 >> 4;

  assign t_r26_c5_0 = p_25_5 << 1;
  assign t_r26_c5_1 = p_26_4 << 1;
  assign t_r26_c5_2 = p_26_5 << 2;
  assign t_r26_c5_3 = p_26_6 << 1;
  assign t_r26_c5_4 = p_27_5 << 1;
  assign t_r26_c5_5 = t_r26_c5_0 + p_25_4;
  assign t_r26_c5_6 = t_r26_c5_1 + p_25_6;
  assign t_r26_c5_7 = t_r26_c5_2 + t_r26_c5_3;
  assign t_r26_c5_8 = t_r26_c5_4 + p_27_4;
  assign t_r26_c5_9 = t_r26_c5_5 + t_r26_c5_6;
  assign t_r26_c5_10 = t_r26_c5_7 + t_r26_c5_8;
  assign t_r26_c5_11 = t_r26_c5_9 + t_r26_c5_10;
  assign t_r26_c5_12 = t_r26_c5_11 + p_27_6;
  assign out_26_5 = t_r26_c5_12 >> 4;

  assign t_r26_c6_0 = p_25_6 << 1;
  assign t_r26_c6_1 = p_26_5 << 1;
  assign t_r26_c6_2 = p_26_6 << 2;
  assign t_r26_c6_3 = p_26_7 << 1;
  assign t_r26_c6_4 = p_27_6 << 1;
  assign t_r26_c6_5 = t_r26_c6_0 + p_25_5;
  assign t_r26_c6_6 = t_r26_c6_1 + p_25_7;
  assign t_r26_c6_7 = t_r26_c6_2 + t_r26_c6_3;
  assign t_r26_c6_8 = t_r26_c6_4 + p_27_5;
  assign t_r26_c6_9 = t_r26_c6_5 + t_r26_c6_6;
  assign t_r26_c6_10 = t_r26_c6_7 + t_r26_c6_8;
  assign t_r26_c6_11 = t_r26_c6_9 + t_r26_c6_10;
  assign t_r26_c6_12 = t_r26_c6_11 + p_27_7;
  assign out_26_6 = t_r26_c6_12 >> 4;

  assign t_r26_c7_0 = p_25_7 << 1;
  assign t_r26_c7_1 = p_26_6 << 1;
  assign t_r26_c7_2 = p_26_7 << 2;
  assign t_r26_c7_3 = p_26_8 << 1;
  assign t_r26_c7_4 = p_27_7 << 1;
  assign t_r26_c7_5 = t_r26_c7_0 + p_25_6;
  assign t_r26_c7_6 = t_r26_c7_1 + p_25_8;
  assign t_r26_c7_7 = t_r26_c7_2 + t_r26_c7_3;
  assign t_r26_c7_8 = t_r26_c7_4 + p_27_6;
  assign t_r26_c7_9 = t_r26_c7_5 + t_r26_c7_6;
  assign t_r26_c7_10 = t_r26_c7_7 + t_r26_c7_8;
  assign t_r26_c7_11 = t_r26_c7_9 + t_r26_c7_10;
  assign t_r26_c7_12 = t_r26_c7_11 + p_27_8;
  assign out_26_7 = t_r26_c7_12 >> 4;

  assign t_r26_c8_0 = p_25_8 << 1;
  assign t_r26_c8_1 = p_26_7 << 1;
  assign t_r26_c8_2 = p_26_8 << 2;
  assign t_r26_c8_3 = p_26_9 << 1;
  assign t_r26_c8_4 = p_27_8 << 1;
  assign t_r26_c8_5 = t_r26_c8_0 + p_25_7;
  assign t_r26_c8_6 = t_r26_c8_1 + p_25_9;
  assign t_r26_c8_7 = t_r26_c8_2 + t_r26_c8_3;
  assign t_r26_c8_8 = t_r26_c8_4 + p_27_7;
  assign t_r26_c8_9 = t_r26_c8_5 + t_r26_c8_6;
  assign t_r26_c8_10 = t_r26_c8_7 + t_r26_c8_8;
  assign t_r26_c8_11 = t_r26_c8_9 + t_r26_c8_10;
  assign t_r26_c8_12 = t_r26_c8_11 + p_27_9;
  assign out_26_8 = t_r26_c8_12 >> 4;

  assign t_r26_c9_0 = p_25_9 << 1;
  assign t_r26_c9_1 = p_26_8 << 1;
  assign t_r26_c9_2 = p_26_9 << 2;
  assign t_r26_c9_3 = p_26_10 << 1;
  assign t_r26_c9_4 = p_27_9 << 1;
  assign t_r26_c9_5 = t_r26_c9_0 + p_25_8;
  assign t_r26_c9_6 = t_r26_c9_1 + p_25_10;
  assign t_r26_c9_7 = t_r26_c9_2 + t_r26_c9_3;
  assign t_r26_c9_8 = t_r26_c9_4 + p_27_8;
  assign t_r26_c9_9 = t_r26_c9_5 + t_r26_c9_6;
  assign t_r26_c9_10 = t_r26_c9_7 + t_r26_c9_8;
  assign t_r26_c9_11 = t_r26_c9_9 + t_r26_c9_10;
  assign t_r26_c9_12 = t_r26_c9_11 + p_27_10;
  assign out_26_9 = t_r26_c9_12 >> 4;

  assign t_r26_c10_0 = p_25_10 << 1;
  assign t_r26_c10_1 = p_26_9 << 1;
  assign t_r26_c10_2 = p_26_10 << 2;
  assign t_r26_c10_3 = p_26_11 << 1;
  assign t_r26_c10_4 = p_27_10 << 1;
  assign t_r26_c10_5 = t_r26_c10_0 + p_25_9;
  assign t_r26_c10_6 = t_r26_c10_1 + p_25_11;
  assign t_r26_c10_7 = t_r26_c10_2 + t_r26_c10_3;
  assign t_r26_c10_8 = t_r26_c10_4 + p_27_9;
  assign t_r26_c10_9 = t_r26_c10_5 + t_r26_c10_6;
  assign t_r26_c10_10 = t_r26_c10_7 + t_r26_c10_8;
  assign t_r26_c10_11 = t_r26_c10_9 + t_r26_c10_10;
  assign t_r26_c10_12 = t_r26_c10_11 + p_27_11;
  assign out_26_10 = t_r26_c10_12 >> 4;

  assign t_r26_c11_0 = p_25_11 << 1;
  assign t_r26_c11_1 = p_26_10 << 1;
  assign t_r26_c11_2 = p_26_11 << 2;
  assign t_r26_c11_3 = p_26_12 << 1;
  assign t_r26_c11_4 = p_27_11 << 1;
  assign t_r26_c11_5 = t_r26_c11_0 + p_25_10;
  assign t_r26_c11_6 = t_r26_c11_1 + p_25_12;
  assign t_r26_c11_7 = t_r26_c11_2 + t_r26_c11_3;
  assign t_r26_c11_8 = t_r26_c11_4 + p_27_10;
  assign t_r26_c11_9 = t_r26_c11_5 + t_r26_c11_6;
  assign t_r26_c11_10 = t_r26_c11_7 + t_r26_c11_8;
  assign t_r26_c11_11 = t_r26_c11_9 + t_r26_c11_10;
  assign t_r26_c11_12 = t_r26_c11_11 + p_27_12;
  assign out_26_11 = t_r26_c11_12 >> 4;

  assign t_r26_c12_0 = p_25_12 << 1;
  assign t_r26_c12_1 = p_26_11 << 1;
  assign t_r26_c12_2 = p_26_12 << 2;
  assign t_r26_c12_3 = p_26_13 << 1;
  assign t_r26_c12_4 = p_27_12 << 1;
  assign t_r26_c12_5 = t_r26_c12_0 + p_25_11;
  assign t_r26_c12_6 = t_r26_c12_1 + p_25_13;
  assign t_r26_c12_7 = t_r26_c12_2 + t_r26_c12_3;
  assign t_r26_c12_8 = t_r26_c12_4 + p_27_11;
  assign t_r26_c12_9 = t_r26_c12_5 + t_r26_c12_6;
  assign t_r26_c12_10 = t_r26_c12_7 + t_r26_c12_8;
  assign t_r26_c12_11 = t_r26_c12_9 + t_r26_c12_10;
  assign t_r26_c12_12 = t_r26_c12_11 + p_27_13;
  assign out_26_12 = t_r26_c12_12 >> 4;

  assign t_r26_c13_0 = p_25_13 << 1;
  assign t_r26_c13_1 = p_26_12 << 1;
  assign t_r26_c13_2 = p_26_13 << 2;
  assign t_r26_c13_3 = p_26_14 << 1;
  assign t_r26_c13_4 = p_27_13 << 1;
  assign t_r26_c13_5 = t_r26_c13_0 + p_25_12;
  assign t_r26_c13_6 = t_r26_c13_1 + p_25_14;
  assign t_r26_c13_7 = t_r26_c13_2 + t_r26_c13_3;
  assign t_r26_c13_8 = t_r26_c13_4 + p_27_12;
  assign t_r26_c13_9 = t_r26_c13_5 + t_r26_c13_6;
  assign t_r26_c13_10 = t_r26_c13_7 + t_r26_c13_8;
  assign t_r26_c13_11 = t_r26_c13_9 + t_r26_c13_10;
  assign t_r26_c13_12 = t_r26_c13_11 + p_27_14;
  assign out_26_13 = t_r26_c13_12 >> 4;

  assign t_r26_c14_0 = p_25_14 << 1;
  assign t_r26_c14_1 = p_26_13 << 1;
  assign t_r26_c14_2 = p_26_14 << 2;
  assign t_r26_c14_3 = p_26_15 << 1;
  assign t_r26_c14_4 = p_27_14 << 1;
  assign t_r26_c14_5 = t_r26_c14_0 + p_25_13;
  assign t_r26_c14_6 = t_r26_c14_1 + p_25_15;
  assign t_r26_c14_7 = t_r26_c14_2 + t_r26_c14_3;
  assign t_r26_c14_8 = t_r26_c14_4 + p_27_13;
  assign t_r26_c14_9 = t_r26_c14_5 + t_r26_c14_6;
  assign t_r26_c14_10 = t_r26_c14_7 + t_r26_c14_8;
  assign t_r26_c14_11 = t_r26_c14_9 + t_r26_c14_10;
  assign t_r26_c14_12 = t_r26_c14_11 + p_27_15;
  assign out_26_14 = t_r26_c14_12 >> 4;

  assign t_r26_c15_0 = p_25_15 << 1;
  assign t_r26_c15_1 = p_26_14 << 1;
  assign t_r26_c15_2 = p_26_15 << 2;
  assign t_r26_c15_3 = p_26_16 << 1;
  assign t_r26_c15_4 = p_27_15 << 1;
  assign t_r26_c15_5 = t_r26_c15_0 + p_25_14;
  assign t_r26_c15_6 = t_r26_c15_1 + p_25_16;
  assign t_r26_c15_7 = t_r26_c15_2 + t_r26_c15_3;
  assign t_r26_c15_8 = t_r26_c15_4 + p_27_14;
  assign t_r26_c15_9 = t_r26_c15_5 + t_r26_c15_6;
  assign t_r26_c15_10 = t_r26_c15_7 + t_r26_c15_8;
  assign t_r26_c15_11 = t_r26_c15_9 + t_r26_c15_10;
  assign t_r26_c15_12 = t_r26_c15_11 + p_27_16;
  assign out_26_15 = t_r26_c15_12 >> 4;

  assign t_r26_c16_0 = p_25_16 << 1;
  assign t_r26_c16_1 = p_26_15 << 1;
  assign t_r26_c16_2 = p_26_16 << 2;
  assign t_r26_c16_3 = p_26_17 << 1;
  assign t_r26_c16_4 = p_27_16 << 1;
  assign t_r26_c16_5 = t_r26_c16_0 + p_25_15;
  assign t_r26_c16_6 = t_r26_c16_1 + p_25_17;
  assign t_r26_c16_7 = t_r26_c16_2 + t_r26_c16_3;
  assign t_r26_c16_8 = t_r26_c16_4 + p_27_15;
  assign t_r26_c16_9 = t_r26_c16_5 + t_r26_c16_6;
  assign t_r26_c16_10 = t_r26_c16_7 + t_r26_c16_8;
  assign t_r26_c16_11 = t_r26_c16_9 + t_r26_c16_10;
  assign t_r26_c16_12 = t_r26_c16_11 + p_27_17;
  assign out_26_16 = t_r26_c16_12 >> 4;

  assign t_r26_c17_0 = p_25_17 << 1;
  assign t_r26_c17_1 = p_26_16 << 1;
  assign t_r26_c17_2 = p_26_17 << 2;
  assign t_r26_c17_3 = p_26_18 << 1;
  assign t_r26_c17_4 = p_27_17 << 1;
  assign t_r26_c17_5 = t_r26_c17_0 + p_25_16;
  assign t_r26_c17_6 = t_r26_c17_1 + p_25_18;
  assign t_r26_c17_7 = t_r26_c17_2 + t_r26_c17_3;
  assign t_r26_c17_8 = t_r26_c17_4 + p_27_16;
  assign t_r26_c17_9 = t_r26_c17_5 + t_r26_c17_6;
  assign t_r26_c17_10 = t_r26_c17_7 + t_r26_c17_8;
  assign t_r26_c17_11 = t_r26_c17_9 + t_r26_c17_10;
  assign t_r26_c17_12 = t_r26_c17_11 + p_27_18;
  assign out_26_17 = t_r26_c17_12 >> 4;

  assign t_r26_c18_0 = p_25_18 << 1;
  assign t_r26_c18_1 = p_26_17 << 1;
  assign t_r26_c18_2 = p_26_18 << 2;
  assign t_r26_c18_3 = p_26_19 << 1;
  assign t_r26_c18_4 = p_27_18 << 1;
  assign t_r26_c18_5 = t_r26_c18_0 + p_25_17;
  assign t_r26_c18_6 = t_r26_c18_1 + p_25_19;
  assign t_r26_c18_7 = t_r26_c18_2 + t_r26_c18_3;
  assign t_r26_c18_8 = t_r26_c18_4 + p_27_17;
  assign t_r26_c18_9 = t_r26_c18_5 + t_r26_c18_6;
  assign t_r26_c18_10 = t_r26_c18_7 + t_r26_c18_8;
  assign t_r26_c18_11 = t_r26_c18_9 + t_r26_c18_10;
  assign t_r26_c18_12 = t_r26_c18_11 + p_27_19;
  assign out_26_18 = t_r26_c18_12 >> 4;

  assign t_r26_c19_0 = p_25_19 << 1;
  assign t_r26_c19_1 = p_26_18 << 1;
  assign t_r26_c19_2 = p_26_19 << 2;
  assign t_r26_c19_3 = p_26_20 << 1;
  assign t_r26_c19_4 = p_27_19 << 1;
  assign t_r26_c19_5 = t_r26_c19_0 + p_25_18;
  assign t_r26_c19_6 = t_r26_c19_1 + p_25_20;
  assign t_r26_c19_7 = t_r26_c19_2 + t_r26_c19_3;
  assign t_r26_c19_8 = t_r26_c19_4 + p_27_18;
  assign t_r26_c19_9 = t_r26_c19_5 + t_r26_c19_6;
  assign t_r26_c19_10 = t_r26_c19_7 + t_r26_c19_8;
  assign t_r26_c19_11 = t_r26_c19_9 + t_r26_c19_10;
  assign t_r26_c19_12 = t_r26_c19_11 + p_27_20;
  assign out_26_19 = t_r26_c19_12 >> 4;

  assign t_r26_c20_0 = p_25_20 << 1;
  assign t_r26_c20_1 = p_26_19 << 1;
  assign t_r26_c20_2 = p_26_20 << 2;
  assign t_r26_c20_3 = p_26_21 << 1;
  assign t_r26_c20_4 = p_27_20 << 1;
  assign t_r26_c20_5 = t_r26_c20_0 + p_25_19;
  assign t_r26_c20_6 = t_r26_c20_1 + p_25_21;
  assign t_r26_c20_7 = t_r26_c20_2 + t_r26_c20_3;
  assign t_r26_c20_8 = t_r26_c20_4 + p_27_19;
  assign t_r26_c20_9 = t_r26_c20_5 + t_r26_c20_6;
  assign t_r26_c20_10 = t_r26_c20_7 + t_r26_c20_8;
  assign t_r26_c20_11 = t_r26_c20_9 + t_r26_c20_10;
  assign t_r26_c20_12 = t_r26_c20_11 + p_27_21;
  assign out_26_20 = t_r26_c20_12 >> 4;

  assign t_r26_c21_0 = p_25_21 << 1;
  assign t_r26_c21_1 = p_26_20 << 1;
  assign t_r26_c21_2 = p_26_21 << 2;
  assign t_r26_c21_3 = p_26_22 << 1;
  assign t_r26_c21_4 = p_27_21 << 1;
  assign t_r26_c21_5 = t_r26_c21_0 + p_25_20;
  assign t_r26_c21_6 = t_r26_c21_1 + p_25_22;
  assign t_r26_c21_7 = t_r26_c21_2 + t_r26_c21_3;
  assign t_r26_c21_8 = t_r26_c21_4 + p_27_20;
  assign t_r26_c21_9 = t_r26_c21_5 + t_r26_c21_6;
  assign t_r26_c21_10 = t_r26_c21_7 + t_r26_c21_8;
  assign t_r26_c21_11 = t_r26_c21_9 + t_r26_c21_10;
  assign t_r26_c21_12 = t_r26_c21_11 + p_27_22;
  assign out_26_21 = t_r26_c21_12 >> 4;

  assign t_r26_c22_0 = p_25_22 << 1;
  assign t_r26_c22_1 = p_26_21 << 1;
  assign t_r26_c22_2 = p_26_22 << 2;
  assign t_r26_c22_3 = p_26_23 << 1;
  assign t_r26_c22_4 = p_27_22 << 1;
  assign t_r26_c22_5 = t_r26_c22_0 + p_25_21;
  assign t_r26_c22_6 = t_r26_c22_1 + p_25_23;
  assign t_r26_c22_7 = t_r26_c22_2 + t_r26_c22_3;
  assign t_r26_c22_8 = t_r26_c22_4 + p_27_21;
  assign t_r26_c22_9 = t_r26_c22_5 + t_r26_c22_6;
  assign t_r26_c22_10 = t_r26_c22_7 + t_r26_c22_8;
  assign t_r26_c22_11 = t_r26_c22_9 + t_r26_c22_10;
  assign t_r26_c22_12 = t_r26_c22_11 + p_27_23;
  assign out_26_22 = t_r26_c22_12 >> 4;

  assign t_r26_c23_0 = p_25_23 << 1;
  assign t_r26_c23_1 = p_26_22 << 1;
  assign t_r26_c23_2 = p_26_23 << 2;
  assign t_r26_c23_3 = p_26_24 << 1;
  assign t_r26_c23_4 = p_27_23 << 1;
  assign t_r26_c23_5 = t_r26_c23_0 + p_25_22;
  assign t_r26_c23_6 = t_r26_c23_1 + p_25_24;
  assign t_r26_c23_7 = t_r26_c23_2 + t_r26_c23_3;
  assign t_r26_c23_8 = t_r26_c23_4 + p_27_22;
  assign t_r26_c23_9 = t_r26_c23_5 + t_r26_c23_6;
  assign t_r26_c23_10 = t_r26_c23_7 + t_r26_c23_8;
  assign t_r26_c23_11 = t_r26_c23_9 + t_r26_c23_10;
  assign t_r26_c23_12 = t_r26_c23_11 + p_27_24;
  assign out_26_23 = t_r26_c23_12 >> 4;

  assign t_r26_c24_0 = p_25_24 << 1;
  assign t_r26_c24_1 = p_26_23 << 1;
  assign t_r26_c24_2 = p_26_24 << 2;
  assign t_r26_c24_3 = p_26_25 << 1;
  assign t_r26_c24_4 = p_27_24 << 1;
  assign t_r26_c24_5 = t_r26_c24_0 + p_25_23;
  assign t_r26_c24_6 = t_r26_c24_1 + p_25_25;
  assign t_r26_c24_7 = t_r26_c24_2 + t_r26_c24_3;
  assign t_r26_c24_8 = t_r26_c24_4 + p_27_23;
  assign t_r26_c24_9 = t_r26_c24_5 + t_r26_c24_6;
  assign t_r26_c24_10 = t_r26_c24_7 + t_r26_c24_8;
  assign t_r26_c24_11 = t_r26_c24_9 + t_r26_c24_10;
  assign t_r26_c24_12 = t_r26_c24_11 + p_27_25;
  assign out_26_24 = t_r26_c24_12 >> 4;

  assign t_r26_c25_0 = p_25_25 << 1;
  assign t_r26_c25_1 = p_26_24 << 1;
  assign t_r26_c25_2 = p_26_25 << 2;
  assign t_r26_c25_3 = p_26_26 << 1;
  assign t_r26_c25_4 = p_27_25 << 1;
  assign t_r26_c25_5 = t_r26_c25_0 + p_25_24;
  assign t_r26_c25_6 = t_r26_c25_1 + p_25_26;
  assign t_r26_c25_7 = t_r26_c25_2 + t_r26_c25_3;
  assign t_r26_c25_8 = t_r26_c25_4 + p_27_24;
  assign t_r26_c25_9 = t_r26_c25_5 + t_r26_c25_6;
  assign t_r26_c25_10 = t_r26_c25_7 + t_r26_c25_8;
  assign t_r26_c25_11 = t_r26_c25_9 + t_r26_c25_10;
  assign t_r26_c25_12 = t_r26_c25_11 + p_27_26;
  assign out_26_25 = t_r26_c25_12 >> 4;

  assign t_r26_c26_0 = p_25_26 << 1;
  assign t_r26_c26_1 = p_26_25 << 1;
  assign t_r26_c26_2 = p_26_26 << 2;
  assign t_r26_c26_3 = p_26_27 << 1;
  assign t_r26_c26_4 = p_27_26 << 1;
  assign t_r26_c26_5 = t_r26_c26_0 + p_25_25;
  assign t_r26_c26_6 = t_r26_c26_1 + p_25_27;
  assign t_r26_c26_7 = t_r26_c26_2 + t_r26_c26_3;
  assign t_r26_c26_8 = t_r26_c26_4 + p_27_25;
  assign t_r26_c26_9 = t_r26_c26_5 + t_r26_c26_6;
  assign t_r26_c26_10 = t_r26_c26_7 + t_r26_c26_8;
  assign t_r26_c26_11 = t_r26_c26_9 + t_r26_c26_10;
  assign t_r26_c26_12 = t_r26_c26_11 + p_27_27;
  assign out_26_26 = t_r26_c26_12 >> 4;

  assign t_r26_c27_0 = p_25_27 << 1;
  assign t_r26_c27_1 = p_26_26 << 1;
  assign t_r26_c27_2 = p_26_27 << 2;
  assign t_r26_c27_3 = p_26_28 << 1;
  assign t_r26_c27_4 = p_27_27 << 1;
  assign t_r26_c27_5 = t_r26_c27_0 + p_25_26;
  assign t_r26_c27_6 = t_r26_c27_1 + p_25_28;
  assign t_r26_c27_7 = t_r26_c27_2 + t_r26_c27_3;
  assign t_r26_c27_8 = t_r26_c27_4 + p_27_26;
  assign t_r26_c27_9 = t_r26_c27_5 + t_r26_c27_6;
  assign t_r26_c27_10 = t_r26_c27_7 + t_r26_c27_8;
  assign t_r26_c27_11 = t_r26_c27_9 + t_r26_c27_10;
  assign t_r26_c27_12 = t_r26_c27_11 + p_27_28;
  assign out_26_27 = t_r26_c27_12 >> 4;

  assign t_r26_c28_0 = p_25_28 << 1;
  assign t_r26_c28_1 = p_26_27 << 1;
  assign t_r26_c28_2 = p_26_28 << 2;
  assign t_r26_c28_3 = p_26_29 << 1;
  assign t_r26_c28_4 = p_27_28 << 1;
  assign t_r26_c28_5 = t_r26_c28_0 + p_25_27;
  assign t_r26_c28_6 = t_r26_c28_1 + p_25_29;
  assign t_r26_c28_7 = t_r26_c28_2 + t_r26_c28_3;
  assign t_r26_c28_8 = t_r26_c28_4 + p_27_27;
  assign t_r26_c28_9 = t_r26_c28_5 + t_r26_c28_6;
  assign t_r26_c28_10 = t_r26_c28_7 + t_r26_c28_8;
  assign t_r26_c28_11 = t_r26_c28_9 + t_r26_c28_10;
  assign t_r26_c28_12 = t_r26_c28_11 + p_27_29;
  assign out_26_28 = t_r26_c28_12 >> 4;

  assign t_r26_c29_0 = p_25_29 << 1;
  assign t_r26_c29_1 = p_26_28 << 1;
  assign t_r26_c29_2 = p_26_29 << 2;
  assign t_r26_c29_3 = p_26_30 << 1;
  assign t_r26_c29_4 = p_27_29 << 1;
  assign t_r26_c29_5 = t_r26_c29_0 + p_25_28;
  assign t_r26_c29_6 = t_r26_c29_1 + p_25_30;
  assign t_r26_c29_7 = t_r26_c29_2 + t_r26_c29_3;
  assign t_r26_c29_8 = t_r26_c29_4 + p_27_28;
  assign t_r26_c29_9 = t_r26_c29_5 + t_r26_c29_6;
  assign t_r26_c29_10 = t_r26_c29_7 + t_r26_c29_8;
  assign t_r26_c29_11 = t_r26_c29_9 + t_r26_c29_10;
  assign t_r26_c29_12 = t_r26_c29_11 + p_27_30;
  assign out_26_29 = t_r26_c29_12 >> 4;

  assign t_r26_c30_0 = p_25_30 << 1;
  assign t_r26_c30_1 = p_26_29 << 1;
  assign t_r26_c30_2 = p_26_30 << 2;
  assign t_r26_c30_3 = p_26_31 << 1;
  assign t_r26_c30_4 = p_27_30 << 1;
  assign t_r26_c30_5 = t_r26_c30_0 + p_25_29;
  assign t_r26_c30_6 = t_r26_c30_1 + p_25_31;
  assign t_r26_c30_7 = t_r26_c30_2 + t_r26_c30_3;
  assign t_r26_c30_8 = t_r26_c30_4 + p_27_29;
  assign t_r26_c30_9 = t_r26_c30_5 + t_r26_c30_6;
  assign t_r26_c30_10 = t_r26_c30_7 + t_r26_c30_8;
  assign t_r26_c30_11 = t_r26_c30_9 + t_r26_c30_10;
  assign t_r26_c30_12 = t_r26_c30_11 + p_27_31;
  assign out_26_30 = t_r26_c30_12 >> 4;

  assign t_r26_c31_0 = p_25_31 << 1;
  assign t_r26_c31_1 = p_26_30 << 1;
  assign t_r26_c31_2 = p_26_31 << 2;
  assign t_r26_c31_3 = p_26_32 << 1;
  assign t_r26_c31_4 = p_27_31 << 1;
  assign t_r26_c31_5 = t_r26_c31_0 + p_25_30;
  assign t_r26_c31_6 = t_r26_c31_1 + p_25_32;
  assign t_r26_c31_7 = t_r26_c31_2 + t_r26_c31_3;
  assign t_r26_c31_8 = t_r26_c31_4 + p_27_30;
  assign t_r26_c31_9 = t_r26_c31_5 + t_r26_c31_6;
  assign t_r26_c31_10 = t_r26_c31_7 + t_r26_c31_8;
  assign t_r26_c31_11 = t_r26_c31_9 + t_r26_c31_10;
  assign t_r26_c31_12 = t_r26_c31_11 + p_27_32;
  assign out_26_31 = t_r26_c31_12 >> 4;

  assign t_r26_c32_0 = p_25_32 << 1;
  assign t_r26_c32_1 = p_26_31 << 1;
  assign t_r26_c32_2 = p_26_32 << 2;
  assign t_r26_c32_3 = p_26_33 << 1;
  assign t_r26_c32_4 = p_27_32 << 1;
  assign t_r26_c32_5 = t_r26_c32_0 + p_25_31;
  assign t_r26_c32_6 = t_r26_c32_1 + p_25_33;
  assign t_r26_c32_7 = t_r26_c32_2 + t_r26_c32_3;
  assign t_r26_c32_8 = t_r26_c32_4 + p_27_31;
  assign t_r26_c32_9 = t_r26_c32_5 + t_r26_c32_6;
  assign t_r26_c32_10 = t_r26_c32_7 + t_r26_c32_8;
  assign t_r26_c32_11 = t_r26_c32_9 + t_r26_c32_10;
  assign t_r26_c32_12 = t_r26_c32_11 + p_27_33;
  assign out_26_32 = t_r26_c32_12 >> 4;

  assign t_r26_c33_0 = p_25_33 << 1;
  assign t_r26_c33_1 = p_26_32 << 1;
  assign t_r26_c33_2 = p_26_33 << 2;
  assign t_r26_c33_3 = p_26_34 << 1;
  assign t_r26_c33_4 = p_27_33 << 1;
  assign t_r26_c33_5 = t_r26_c33_0 + p_25_32;
  assign t_r26_c33_6 = t_r26_c33_1 + p_25_34;
  assign t_r26_c33_7 = t_r26_c33_2 + t_r26_c33_3;
  assign t_r26_c33_8 = t_r26_c33_4 + p_27_32;
  assign t_r26_c33_9 = t_r26_c33_5 + t_r26_c33_6;
  assign t_r26_c33_10 = t_r26_c33_7 + t_r26_c33_8;
  assign t_r26_c33_11 = t_r26_c33_9 + t_r26_c33_10;
  assign t_r26_c33_12 = t_r26_c33_11 + p_27_34;
  assign out_26_33 = t_r26_c33_12 >> 4;

  assign t_r26_c34_0 = p_25_34 << 1;
  assign t_r26_c34_1 = p_26_33 << 1;
  assign t_r26_c34_2 = p_26_34 << 2;
  assign t_r26_c34_3 = p_26_35 << 1;
  assign t_r26_c34_4 = p_27_34 << 1;
  assign t_r26_c34_5 = t_r26_c34_0 + p_25_33;
  assign t_r26_c34_6 = t_r26_c34_1 + p_25_35;
  assign t_r26_c34_7 = t_r26_c34_2 + t_r26_c34_3;
  assign t_r26_c34_8 = t_r26_c34_4 + p_27_33;
  assign t_r26_c34_9 = t_r26_c34_5 + t_r26_c34_6;
  assign t_r26_c34_10 = t_r26_c34_7 + t_r26_c34_8;
  assign t_r26_c34_11 = t_r26_c34_9 + t_r26_c34_10;
  assign t_r26_c34_12 = t_r26_c34_11 + p_27_35;
  assign out_26_34 = t_r26_c34_12 >> 4;

  assign t_r26_c35_0 = p_25_35 << 1;
  assign t_r26_c35_1 = p_26_34 << 1;
  assign t_r26_c35_2 = p_26_35 << 2;
  assign t_r26_c35_3 = p_26_36 << 1;
  assign t_r26_c35_4 = p_27_35 << 1;
  assign t_r26_c35_5 = t_r26_c35_0 + p_25_34;
  assign t_r26_c35_6 = t_r26_c35_1 + p_25_36;
  assign t_r26_c35_7 = t_r26_c35_2 + t_r26_c35_3;
  assign t_r26_c35_8 = t_r26_c35_4 + p_27_34;
  assign t_r26_c35_9 = t_r26_c35_5 + t_r26_c35_6;
  assign t_r26_c35_10 = t_r26_c35_7 + t_r26_c35_8;
  assign t_r26_c35_11 = t_r26_c35_9 + t_r26_c35_10;
  assign t_r26_c35_12 = t_r26_c35_11 + p_27_36;
  assign out_26_35 = t_r26_c35_12 >> 4;

  assign t_r26_c36_0 = p_25_36 << 1;
  assign t_r26_c36_1 = p_26_35 << 1;
  assign t_r26_c36_2 = p_26_36 << 2;
  assign t_r26_c36_3 = p_26_37 << 1;
  assign t_r26_c36_4 = p_27_36 << 1;
  assign t_r26_c36_5 = t_r26_c36_0 + p_25_35;
  assign t_r26_c36_6 = t_r26_c36_1 + p_25_37;
  assign t_r26_c36_7 = t_r26_c36_2 + t_r26_c36_3;
  assign t_r26_c36_8 = t_r26_c36_4 + p_27_35;
  assign t_r26_c36_9 = t_r26_c36_5 + t_r26_c36_6;
  assign t_r26_c36_10 = t_r26_c36_7 + t_r26_c36_8;
  assign t_r26_c36_11 = t_r26_c36_9 + t_r26_c36_10;
  assign t_r26_c36_12 = t_r26_c36_11 + p_27_37;
  assign out_26_36 = t_r26_c36_12 >> 4;

  assign t_r26_c37_0 = p_25_37 << 1;
  assign t_r26_c37_1 = p_26_36 << 1;
  assign t_r26_c37_2 = p_26_37 << 2;
  assign t_r26_c37_3 = p_26_38 << 1;
  assign t_r26_c37_4 = p_27_37 << 1;
  assign t_r26_c37_5 = t_r26_c37_0 + p_25_36;
  assign t_r26_c37_6 = t_r26_c37_1 + p_25_38;
  assign t_r26_c37_7 = t_r26_c37_2 + t_r26_c37_3;
  assign t_r26_c37_8 = t_r26_c37_4 + p_27_36;
  assign t_r26_c37_9 = t_r26_c37_5 + t_r26_c37_6;
  assign t_r26_c37_10 = t_r26_c37_7 + t_r26_c37_8;
  assign t_r26_c37_11 = t_r26_c37_9 + t_r26_c37_10;
  assign t_r26_c37_12 = t_r26_c37_11 + p_27_38;
  assign out_26_37 = t_r26_c37_12 >> 4;

  assign t_r26_c38_0 = p_25_38 << 1;
  assign t_r26_c38_1 = p_26_37 << 1;
  assign t_r26_c38_2 = p_26_38 << 2;
  assign t_r26_c38_3 = p_26_39 << 1;
  assign t_r26_c38_4 = p_27_38 << 1;
  assign t_r26_c38_5 = t_r26_c38_0 + p_25_37;
  assign t_r26_c38_6 = t_r26_c38_1 + p_25_39;
  assign t_r26_c38_7 = t_r26_c38_2 + t_r26_c38_3;
  assign t_r26_c38_8 = t_r26_c38_4 + p_27_37;
  assign t_r26_c38_9 = t_r26_c38_5 + t_r26_c38_6;
  assign t_r26_c38_10 = t_r26_c38_7 + t_r26_c38_8;
  assign t_r26_c38_11 = t_r26_c38_9 + t_r26_c38_10;
  assign t_r26_c38_12 = t_r26_c38_11 + p_27_39;
  assign out_26_38 = t_r26_c38_12 >> 4;

  assign t_r26_c39_0 = p_25_39 << 1;
  assign t_r26_c39_1 = p_26_38 << 1;
  assign t_r26_c39_2 = p_26_39 << 2;
  assign t_r26_c39_3 = p_26_40 << 1;
  assign t_r26_c39_4 = p_27_39 << 1;
  assign t_r26_c39_5 = t_r26_c39_0 + p_25_38;
  assign t_r26_c39_6 = t_r26_c39_1 + p_25_40;
  assign t_r26_c39_7 = t_r26_c39_2 + t_r26_c39_3;
  assign t_r26_c39_8 = t_r26_c39_4 + p_27_38;
  assign t_r26_c39_9 = t_r26_c39_5 + t_r26_c39_6;
  assign t_r26_c39_10 = t_r26_c39_7 + t_r26_c39_8;
  assign t_r26_c39_11 = t_r26_c39_9 + t_r26_c39_10;
  assign t_r26_c39_12 = t_r26_c39_11 + p_27_40;
  assign out_26_39 = t_r26_c39_12 >> 4;

  assign t_r26_c40_0 = p_25_40 << 1;
  assign t_r26_c40_1 = p_26_39 << 1;
  assign t_r26_c40_2 = p_26_40 << 2;
  assign t_r26_c40_3 = p_26_41 << 1;
  assign t_r26_c40_4 = p_27_40 << 1;
  assign t_r26_c40_5 = t_r26_c40_0 + p_25_39;
  assign t_r26_c40_6 = t_r26_c40_1 + p_25_41;
  assign t_r26_c40_7 = t_r26_c40_2 + t_r26_c40_3;
  assign t_r26_c40_8 = t_r26_c40_4 + p_27_39;
  assign t_r26_c40_9 = t_r26_c40_5 + t_r26_c40_6;
  assign t_r26_c40_10 = t_r26_c40_7 + t_r26_c40_8;
  assign t_r26_c40_11 = t_r26_c40_9 + t_r26_c40_10;
  assign t_r26_c40_12 = t_r26_c40_11 + p_27_41;
  assign out_26_40 = t_r26_c40_12 >> 4;

  assign t_r26_c41_0 = p_25_41 << 1;
  assign t_r26_c41_1 = p_26_40 << 1;
  assign t_r26_c41_2 = p_26_41 << 2;
  assign t_r26_c41_3 = p_26_42 << 1;
  assign t_r26_c41_4 = p_27_41 << 1;
  assign t_r26_c41_5 = t_r26_c41_0 + p_25_40;
  assign t_r26_c41_6 = t_r26_c41_1 + p_25_42;
  assign t_r26_c41_7 = t_r26_c41_2 + t_r26_c41_3;
  assign t_r26_c41_8 = t_r26_c41_4 + p_27_40;
  assign t_r26_c41_9 = t_r26_c41_5 + t_r26_c41_6;
  assign t_r26_c41_10 = t_r26_c41_7 + t_r26_c41_8;
  assign t_r26_c41_11 = t_r26_c41_9 + t_r26_c41_10;
  assign t_r26_c41_12 = t_r26_c41_11 + p_27_42;
  assign out_26_41 = t_r26_c41_12 >> 4;

  assign t_r26_c42_0 = p_25_42 << 1;
  assign t_r26_c42_1 = p_26_41 << 1;
  assign t_r26_c42_2 = p_26_42 << 2;
  assign t_r26_c42_3 = p_26_43 << 1;
  assign t_r26_c42_4 = p_27_42 << 1;
  assign t_r26_c42_5 = t_r26_c42_0 + p_25_41;
  assign t_r26_c42_6 = t_r26_c42_1 + p_25_43;
  assign t_r26_c42_7 = t_r26_c42_2 + t_r26_c42_3;
  assign t_r26_c42_8 = t_r26_c42_4 + p_27_41;
  assign t_r26_c42_9 = t_r26_c42_5 + t_r26_c42_6;
  assign t_r26_c42_10 = t_r26_c42_7 + t_r26_c42_8;
  assign t_r26_c42_11 = t_r26_c42_9 + t_r26_c42_10;
  assign t_r26_c42_12 = t_r26_c42_11 + p_27_43;
  assign out_26_42 = t_r26_c42_12 >> 4;

  assign t_r26_c43_0 = p_25_43 << 1;
  assign t_r26_c43_1 = p_26_42 << 1;
  assign t_r26_c43_2 = p_26_43 << 2;
  assign t_r26_c43_3 = p_26_44 << 1;
  assign t_r26_c43_4 = p_27_43 << 1;
  assign t_r26_c43_5 = t_r26_c43_0 + p_25_42;
  assign t_r26_c43_6 = t_r26_c43_1 + p_25_44;
  assign t_r26_c43_7 = t_r26_c43_2 + t_r26_c43_3;
  assign t_r26_c43_8 = t_r26_c43_4 + p_27_42;
  assign t_r26_c43_9 = t_r26_c43_5 + t_r26_c43_6;
  assign t_r26_c43_10 = t_r26_c43_7 + t_r26_c43_8;
  assign t_r26_c43_11 = t_r26_c43_9 + t_r26_c43_10;
  assign t_r26_c43_12 = t_r26_c43_11 + p_27_44;
  assign out_26_43 = t_r26_c43_12 >> 4;

  assign t_r26_c44_0 = p_25_44 << 1;
  assign t_r26_c44_1 = p_26_43 << 1;
  assign t_r26_c44_2 = p_26_44 << 2;
  assign t_r26_c44_3 = p_26_45 << 1;
  assign t_r26_c44_4 = p_27_44 << 1;
  assign t_r26_c44_5 = t_r26_c44_0 + p_25_43;
  assign t_r26_c44_6 = t_r26_c44_1 + p_25_45;
  assign t_r26_c44_7 = t_r26_c44_2 + t_r26_c44_3;
  assign t_r26_c44_8 = t_r26_c44_4 + p_27_43;
  assign t_r26_c44_9 = t_r26_c44_5 + t_r26_c44_6;
  assign t_r26_c44_10 = t_r26_c44_7 + t_r26_c44_8;
  assign t_r26_c44_11 = t_r26_c44_9 + t_r26_c44_10;
  assign t_r26_c44_12 = t_r26_c44_11 + p_27_45;
  assign out_26_44 = t_r26_c44_12 >> 4;

  assign t_r26_c45_0 = p_25_45 << 1;
  assign t_r26_c45_1 = p_26_44 << 1;
  assign t_r26_c45_2 = p_26_45 << 2;
  assign t_r26_c45_3 = p_26_46 << 1;
  assign t_r26_c45_4 = p_27_45 << 1;
  assign t_r26_c45_5 = t_r26_c45_0 + p_25_44;
  assign t_r26_c45_6 = t_r26_c45_1 + p_25_46;
  assign t_r26_c45_7 = t_r26_c45_2 + t_r26_c45_3;
  assign t_r26_c45_8 = t_r26_c45_4 + p_27_44;
  assign t_r26_c45_9 = t_r26_c45_5 + t_r26_c45_6;
  assign t_r26_c45_10 = t_r26_c45_7 + t_r26_c45_8;
  assign t_r26_c45_11 = t_r26_c45_9 + t_r26_c45_10;
  assign t_r26_c45_12 = t_r26_c45_11 + p_27_46;
  assign out_26_45 = t_r26_c45_12 >> 4;

  assign t_r26_c46_0 = p_25_46 << 1;
  assign t_r26_c46_1 = p_26_45 << 1;
  assign t_r26_c46_2 = p_26_46 << 2;
  assign t_r26_c46_3 = p_26_47 << 1;
  assign t_r26_c46_4 = p_27_46 << 1;
  assign t_r26_c46_5 = t_r26_c46_0 + p_25_45;
  assign t_r26_c46_6 = t_r26_c46_1 + p_25_47;
  assign t_r26_c46_7 = t_r26_c46_2 + t_r26_c46_3;
  assign t_r26_c46_8 = t_r26_c46_4 + p_27_45;
  assign t_r26_c46_9 = t_r26_c46_5 + t_r26_c46_6;
  assign t_r26_c46_10 = t_r26_c46_7 + t_r26_c46_8;
  assign t_r26_c46_11 = t_r26_c46_9 + t_r26_c46_10;
  assign t_r26_c46_12 = t_r26_c46_11 + p_27_47;
  assign out_26_46 = t_r26_c46_12 >> 4;

  assign t_r26_c47_0 = p_25_47 << 1;
  assign t_r26_c47_1 = p_26_46 << 1;
  assign t_r26_c47_2 = p_26_47 << 2;
  assign t_r26_c47_3 = p_26_48 << 1;
  assign t_r26_c47_4 = p_27_47 << 1;
  assign t_r26_c47_5 = t_r26_c47_0 + p_25_46;
  assign t_r26_c47_6 = t_r26_c47_1 + p_25_48;
  assign t_r26_c47_7 = t_r26_c47_2 + t_r26_c47_3;
  assign t_r26_c47_8 = t_r26_c47_4 + p_27_46;
  assign t_r26_c47_9 = t_r26_c47_5 + t_r26_c47_6;
  assign t_r26_c47_10 = t_r26_c47_7 + t_r26_c47_8;
  assign t_r26_c47_11 = t_r26_c47_9 + t_r26_c47_10;
  assign t_r26_c47_12 = t_r26_c47_11 + p_27_48;
  assign out_26_47 = t_r26_c47_12 >> 4;

  assign t_r26_c48_0 = p_25_48 << 1;
  assign t_r26_c48_1 = p_26_47 << 1;
  assign t_r26_c48_2 = p_26_48 << 2;
  assign t_r26_c48_3 = p_26_49 << 1;
  assign t_r26_c48_4 = p_27_48 << 1;
  assign t_r26_c48_5 = t_r26_c48_0 + p_25_47;
  assign t_r26_c48_6 = t_r26_c48_1 + p_25_49;
  assign t_r26_c48_7 = t_r26_c48_2 + t_r26_c48_3;
  assign t_r26_c48_8 = t_r26_c48_4 + p_27_47;
  assign t_r26_c48_9 = t_r26_c48_5 + t_r26_c48_6;
  assign t_r26_c48_10 = t_r26_c48_7 + t_r26_c48_8;
  assign t_r26_c48_11 = t_r26_c48_9 + t_r26_c48_10;
  assign t_r26_c48_12 = t_r26_c48_11 + p_27_49;
  assign out_26_48 = t_r26_c48_12 >> 4;

  assign t_r26_c49_0 = p_25_49 << 1;
  assign t_r26_c49_1 = p_26_48 << 1;
  assign t_r26_c49_2 = p_26_49 << 2;
  assign t_r26_c49_3 = p_26_50 << 1;
  assign t_r26_c49_4 = p_27_49 << 1;
  assign t_r26_c49_5 = t_r26_c49_0 + p_25_48;
  assign t_r26_c49_6 = t_r26_c49_1 + p_25_50;
  assign t_r26_c49_7 = t_r26_c49_2 + t_r26_c49_3;
  assign t_r26_c49_8 = t_r26_c49_4 + p_27_48;
  assign t_r26_c49_9 = t_r26_c49_5 + t_r26_c49_6;
  assign t_r26_c49_10 = t_r26_c49_7 + t_r26_c49_8;
  assign t_r26_c49_11 = t_r26_c49_9 + t_r26_c49_10;
  assign t_r26_c49_12 = t_r26_c49_11 + p_27_50;
  assign out_26_49 = t_r26_c49_12 >> 4;

  assign t_r26_c50_0 = p_25_50 << 1;
  assign t_r26_c50_1 = p_26_49 << 1;
  assign t_r26_c50_2 = p_26_50 << 2;
  assign t_r26_c50_3 = p_26_51 << 1;
  assign t_r26_c50_4 = p_27_50 << 1;
  assign t_r26_c50_5 = t_r26_c50_0 + p_25_49;
  assign t_r26_c50_6 = t_r26_c50_1 + p_25_51;
  assign t_r26_c50_7 = t_r26_c50_2 + t_r26_c50_3;
  assign t_r26_c50_8 = t_r26_c50_4 + p_27_49;
  assign t_r26_c50_9 = t_r26_c50_5 + t_r26_c50_6;
  assign t_r26_c50_10 = t_r26_c50_7 + t_r26_c50_8;
  assign t_r26_c50_11 = t_r26_c50_9 + t_r26_c50_10;
  assign t_r26_c50_12 = t_r26_c50_11 + p_27_51;
  assign out_26_50 = t_r26_c50_12 >> 4;

  assign t_r26_c51_0 = p_25_51 << 1;
  assign t_r26_c51_1 = p_26_50 << 1;
  assign t_r26_c51_2 = p_26_51 << 2;
  assign t_r26_c51_3 = p_26_52 << 1;
  assign t_r26_c51_4 = p_27_51 << 1;
  assign t_r26_c51_5 = t_r26_c51_0 + p_25_50;
  assign t_r26_c51_6 = t_r26_c51_1 + p_25_52;
  assign t_r26_c51_7 = t_r26_c51_2 + t_r26_c51_3;
  assign t_r26_c51_8 = t_r26_c51_4 + p_27_50;
  assign t_r26_c51_9 = t_r26_c51_5 + t_r26_c51_6;
  assign t_r26_c51_10 = t_r26_c51_7 + t_r26_c51_8;
  assign t_r26_c51_11 = t_r26_c51_9 + t_r26_c51_10;
  assign t_r26_c51_12 = t_r26_c51_11 + p_27_52;
  assign out_26_51 = t_r26_c51_12 >> 4;

  assign t_r26_c52_0 = p_25_52 << 1;
  assign t_r26_c52_1 = p_26_51 << 1;
  assign t_r26_c52_2 = p_26_52 << 2;
  assign t_r26_c52_3 = p_26_53 << 1;
  assign t_r26_c52_4 = p_27_52 << 1;
  assign t_r26_c52_5 = t_r26_c52_0 + p_25_51;
  assign t_r26_c52_6 = t_r26_c52_1 + p_25_53;
  assign t_r26_c52_7 = t_r26_c52_2 + t_r26_c52_3;
  assign t_r26_c52_8 = t_r26_c52_4 + p_27_51;
  assign t_r26_c52_9 = t_r26_c52_5 + t_r26_c52_6;
  assign t_r26_c52_10 = t_r26_c52_7 + t_r26_c52_8;
  assign t_r26_c52_11 = t_r26_c52_9 + t_r26_c52_10;
  assign t_r26_c52_12 = t_r26_c52_11 + p_27_53;
  assign out_26_52 = t_r26_c52_12 >> 4;

  assign t_r26_c53_0 = p_25_53 << 1;
  assign t_r26_c53_1 = p_26_52 << 1;
  assign t_r26_c53_2 = p_26_53 << 2;
  assign t_r26_c53_3 = p_26_54 << 1;
  assign t_r26_c53_4 = p_27_53 << 1;
  assign t_r26_c53_5 = t_r26_c53_0 + p_25_52;
  assign t_r26_c53_6 = t_r26_c53_1 + p_25_54;
  assign t_r26_c53_7 = t_r26_c53_2 + t_r26_c53_3;
  assign t_r26_c53_8 = t_r26_c53_4 + p_27_52;
  assign t_r26_c53_9 = t_r26_c53_5 + t_r26_c53_6;
  assign t_r26_c53_10 = t_r26_c53_7 + t_r26_c53_8;
  assign t_r26_c53_11 = t_r26_c53_9 + t_r26_c53_10;
  assign t_r26_c53_12 = t_r26_c53_11 + p_27_54;
  assign out_26_53 = t_r26_c53_12 >> 4;

  assign t_r26_c54_0 = p_25_54 << 1;
  assign t_r26_c54_1 = p_26_53 << 1;
  assign t_r26_c54_2 = p_26_54 << 2;
  assign t_r26_c54_3 = p_26_55 << 1;
  assign t_r26_c54_4 = p_27_54 << 1;
  assign t_r26_c54_5 = t_r26_c54_0 + p_25_53;
  assign t_r26_c54_6 = t_r26_c54_1 + p_25_55;
  assign t_r26_c54_7 = t_r26_c54_2 + t_r26_c54_3;
  assign t_r26_c54_8 = t_r26_c54_4 + p_27_53;
  assign t_r26_c54_9 = t_r26_c54_5 + t_r26_c54_6;
  assign t_r26_c54_10 = t_r26_c54_7 + t_r26_c54_8;
  assign t_r26_c54_11 = t_r26_c54_9 + t_r26_c54_10;
  assign t_r26_c54_12 = t_r26_c54_11 + p_27_55;
  assign out_26_54 = t_r26_c54_12 >> 4;

  assign t_r26_c55_0 = p_25_55 << 1;
  assign t_r26_c55_1 = p_26_54 << 1;
  assign t_r26_c55_2 = p_26_55 << 2;
  assign t_r26_c55_3 = p_26_56 << 1;
  assign t_r26_c55_4 = p_27_55 << 1;
  assign t_r26_c55_5 = t_r26_c55_0 + p_25_54;
  assign t_r26_c55_6 = t_r26_c55_1 + p_25_56;
  assign t_r26_c55_7 = t_r26_c55_2 + t_r26_c55_3;
  assign t_r26_c55_8 = t_r26_c55_4 + p_27_54;
  assign t_r26_c55_9 = t_r26_c55_5 + t_r26_c55_6;
  assign t_r26_c55_10 = t_r26_c55_7 + t_r26_c55_8;
  assign t_r26_c55_11 = t_r26_c55_9 + t_r26_c55_10;
  assign t_r26_c55_12 = t_r26_c55_11 + p_27_56;
  assign out_26_55 = t_r26_c55_12 >> 4;

  assign t_r26_c56_0 = p_25_56 << 1;
  assign t_r26_c56_1 = p_26_55 << 1;
  assign t_r26_c56_2 = p_26_56 << 2;
  assign t_r26_c56_3 = p_26_57 << 1;
  assign t_r26_c56_4 = p_27_56 << 1;
  assign t_r26_c56_5 = t_r26_c56_0 + p_25_55;
  assign t_r26_c56_6 = t_r26_c56_1 + p_25_57;
  assign t_r26_c56_7 = t_r26_c56_2 + t_r26_c56_3;
  assign t_r26_c56_8 = t_r26_c56_4 + p_27_55;
  assign t_r26_c56_9 = t_r26_c56_5 + t_r26_c56_6;
  assign t_r26_c56_10 = t_r26_c56_7 + t_r26_c56_8;
  assign t_r26_c56_11 = t_r26_c56_9 + t_r26_c56_10;
  assign t_r26_c56_12 = t_r26_c56_11 + p_27_57;
  assign out_26_56 = t_r26_c56_12 >> 4;

  assign t_r26_c57_0 = p_25_57 << 1;
  assign t_r26_c57_1 = p_26_56 << 1;
  assign t_r26_c57_2 = p_26_57 << 2;
  assign t_r26_c57_3 = p_26_58 << 1;
  assign t_r26_c57_4 = p_27_57 << 1;
  assign t_r26_c57_5 = t_r26_c57_0 + p_25_56;
  assign t_r26_c57_6 = t_r26_c57_1 + p_25_58;
  assign t_r26_c57_7 = t_r26_c57_2 + t_r26_c57_3;
  assign t_r26_c57_8 = t_r26_c57_4 + p_27_56;
  assign t_r26_c57_9 = t_r26_c57_5 + t_r26_c57_6;
  assign t_r26_c57_10 = t_r26_c57_7 + t_r26_c57_8;
  assign t_r26_c57_11 = t_r26_c57_9 + t_r26_c57_10;
  assign t_r26_c57_12 = t_r26_c57_11 + p_27_58;
  assign out_26_57 = t_r26_c57_12 >> 4;

  assign t_r26_c58_0 = p_25_58 << 1;
  assign t_r26_c58_1 = p_26_57 << 1;
  assign t_r26_c58_2 = p_26_58 << 2;
  assign t_r26_c58_3 = p_26_59 << 1;
  assign t_r26_c58_4 = p_27_58 << 1;
  assign t_r26_c58_5 = t_r26_c58_0 + p_25_57;
  assign t_r26_c58_6 = t_r26_c58_1 + p_25_59;
  assign t_r26_c58_7 = t_r26_c58_2 + t_r26_c58_3;
  assign t_r26_c58_8 = t_r26_c58_4 + p_27_57;
  assign t_r26_c58_9 = t_r26_c58_5 + t_r26_c58_6;
  assign t_r26_c58_10 = t_r26_c58_7 + t_r26_c58_8;
  assign t_r26_c58_11 = t_r26_c58_9 + t_r26_c58_10;
  assign t_r26_c58_12 = t_r26_c58_11 + p_27_59;
  assign out_26_58 = t_r26_c58_12 >> 4;

  assign t_r26_c59_0 = p_25_59 << 1;
  assign t_r26_c59_1 = p_26_58 << 1;
  assign t_r26_c59_2 = p_26_59 << 2;
  assign t_r26_c59_3 = p_26_60 << 1;
  assign t_r26_c59_4 = p_27_59 << 1;
  assign t_r26_c59_5 = t_r26_c59_0 + p_25_58;
  assign t_r26_c59_6 = t_r26_c59_1 + p_25_60;
  assign t_r26_c59_7 = t_r26_c59_2 + t_r26_c59_3;
  assign t_r26_c59_8 = t_r26_c59_4 + p_27_58;
  assign t_r26_c59_9 = t_r26_c59_5 + t_r26_c59_6;
  assign t_r26_c59_10 = t_r26_c59_7 + t_r26_c59_8;
  assign t_r26_c59_11 = t_r26_c59_9 + t_r26_c59_10;
  assign t_r26_c59_12 = t_r26_c59_11 + p_27_60;
  assign out_26_59 = t_r26_c59_12 >> 4;

  assign t_r26_c60_0 = p_25_60 << 1;
  assign t_r26_c60_1 = p_26_59 << 1;
  assign t_r26_c60_2 = p_26_60 << 2;
  assign t_r26_c60_3 = p_26_61 << 1;
  assign t_r26_c60_4 = p_27_60 << 1;
  assign t_r26_c60_5 = t_r26_c60_0 + p_25_59;
  assign t_r26_c60_6 = t_r26_c60_1 + p_25_61;
  assign t_r26_c60_7 = t_r26_c60_2 + t_r26_c60_3;
  assign t_r26_c60_8 = t_r26_c60_4 + p_27_59;
  assign t_r26_c60_9 = t_r26_c60_5 + t_r26_c60_6;
  assign t_r26_c60_10 = t_r26_c60_7 + t_r26_c60_8;
  assign t_r26_c60_11 = t_r26_c60_9 + t_r26_c60_10;
  assign t_r26_c60_12 = t_r26_c60_11 + p_27_61;
  assign out_26_60 = t_r26_c60_12 >> 4;

  assign t_r26_c61_0 = p_25_61 << 1;
  assign t_r26_c61_1 = p_26_60 << 1;
  assign t_r26_c61_2 = p_26_61 << 2;
  assign t_r26_c61_3 = p_26_62 << 1;
  assign t_r26_c61_4 = p_27_61 << 1;
  assign t_r26_c61_5 = t_r26_c61_0 + p_25_60;
  assign t_r26_c61_6 = t_r26_c61_1 + p_25_62;
  assign t_r26_c61_7 = t_r26_c61_2 + t_r26_c61_3;
  assign t_r26_c61_8 = t_r26_c61_4 + p_27_60;
  assign t_r26_c61_9 = t_r26_c61_5 + t_r26_c61_6;
  assign t_r26_c61_10 = t_r26_c61_7 + t_r26_c61_8;
  assign t_r26_c61_11 = t_r26_c61_9 + t_r26_c61_10;
  assign t_r26_c61_12 = t_r26_c61_11 + p_27_62;
  assign out_26_61 = t_r26_c61_12 >> 4;

  assign t_r26_c62_0 = p_25_62 << 1;
  assign t_r26_c62_1 = p_26_61 << 1;
  assign t_r26_c62_2 = p_26_62 << 2;
  assign t_r26_c62_3 = p_26_63 << 1;
  assign t_r26_c62_4 = p_27_62 << 1;
  assign t_r26_c62_5 = t_r26_c62_0 + p_25_61;
  assign t_r26_c62_6 = t_r26_c62_1 + p_25_63;
  assign t_r26_c62_7 = t_r26_c62_2 + t_r26_c62_3;
  assign t_r26_c62_8 = t_r26_c62_4 + p_27_61;
  assign t_r26_c62_9 = t_r26_c62_5 + t_r26_c62_6;
  assign t_r26_c62_10 = t_r26_c62_7 + t_r26_c62_8;
  assign t_r26_c62_11 = t_r26_c62_9 + t_r26_c62_10;
  assign t_r26_c62_12 = t_r26_c62_11 + p_27_63;
  assign out_26_62 = t_r26_c62_12 >> 4;

  assign t_r26_c63_0 = p_25_63 << 1;
  assign t_r26_c63_1 = p_26_62 << 1;
  assign t_r26_c63_2 = p_26_63 << 2;
  assign t_r26_c63_3 = p_26_64 << 1;
  assign t_r26_c63_4 = p_27_63 << 1;
  assign t_r26_c63_5 = t_r26_c63_0 + p_25_62;
  assign t_r26_c63_6 = t_r26_c63_1 + p_25_64;
  assign t_r26_c63_7 = t_r26_c63_2 + t_r26_c63_3;
  assign t_r26_c63_8 = t_r26_c63_4 + p_27_62;
  assign t_r26_c63_9 = t_r26_c63_5 + t_r26_c63_6;
  assign t_r26_c63_10 = t_r26_c63_7 + t_r26_c63_8;
  assign t_r26_c63_11 = t_r26_c63_9 + t_r26_c63_10;
  assign t_r26_c63_12 = t_r26_c63_11 + p_27_64;
  assign out_26_63 = t_r26_c63_12 >> 4;

  assign t_r26_c64_0 = p_25_64 << 1;
  assign t_r26_c64_1 = p_26_63 << 1;
  assign t_r26_c64_2 = p_26_64 << 2;
  assign t_r26_c64_3 = p_26_65 << 1;
  assign t_r26_c64_4 = p_27_64 << 1;
  assign t_r26_c64_5 = t_r26_c64_0 + p_25_63;
  assign t_r26_c64_6 = t_r26_c64_1 + p_25_65;
  assign t_r26_c64_7 = t_r26_c64_2 + t_r26_c64_3;
  assign t_r26_c64_8 = t_r26_c64_4 + p_27_63;
  assign t_r26_c64_9 = t_r26_c64_5 + t_r26_c64_6;
  assign t_r26_c64_10 = t_r26_c64_7 + t_r26_c64_8;
  assign t_r26_c64_11 = t_r26_c64_9 + t_r26_c64_10;
  assign t_r26_c64_12 = t_r26_c64_11 + p_27_65;
  assign out_26_64 = t_r26_c64_12 >> 4;

  assign t_r27_c1_0 = p_26_1 << 1;
  assign t_r27_c1_1 = p_27_0 << 1;
  assign t_r27_c1_2 = p_27_1 << 2;
  assign t_r27_c1_3 = p_27_2 << 1;
  assign t_r27_c1_4 = p_28_1 << 1;
  assign t_r27_c1_5 = t_r27_c1_0 + p_26_0;
  assign t_r27_c1_6 = t_r27_c1_1 + p_26_2;
  assign t_r27_c1_7 = t_r27_c1_2 + t_r27_c1_3;
  assign t_r27_c1_8 = t_r27_c1_4 + p_28_0;
  assign t_r27_c1_9 = t_r27_c1_5 + t_r27_c1_6;
  assign t_r27_c1_10 = t_r27_c1_7 + t_r27_c1_8;
  assign t_r27_c1_11 = t_r27_c1_9 + t_r27_c1_10;
  assign t_r27_c1_12 = t_r27_c1_11 + p_28_2;
  assign out_27_1 = t_r27_c1_12 >> 4;

  assign t_r27_c2_0 = p_26_2 << 1;
  assign t_r27_c2_1 = p_27_1 << 1;
  assign t_r27_c2_2 = p_27_2 << 2;
  assign t_r27_c2_3 = p_27_3 << 1;
  assign t_r27_c2_4 = p_28_2 << 1;
  assign t_r27_c2_5 = t_r27_c2_0 + p_26_1;
  assign t_r27_c2_6 = t_r27_c2_1 + p_26_3;
  assign t_r27_c2_7 = t_r27_c2_2 + t_r27_c2_3;
  assign t_r27_c2_8 = t_r27_c2_4 + p_28_1;
  assign t_r27_c2_9 = t_r27_c2_5 + t_r27_c2_6;
  assign t_r27_c2_10 = t_r27_c2_7 + t_r27_c2_8;
  assign t_r27_c2_11 = t_r27_c2_9 + t_r27_c2_10;
  assign t_r27_c2_12 = t_r27_c2_11 + p_28_3;
  assign out_27_2 = t_r27_c2_12 >> 4;

  assign t_r27_c3_0 = p_26_3 << 1;
  assign t_r27_c3_1 = p_27_2 << 1;
  assign t_r27_c3_2 = p_27_3 << 2;
  assign t_r27_c3_3 = p_27_4 << 1;
  assign t_r27_c3_4 = p_28_3 << 1;
  assign t_r27_c3_5 = t_r27_c3_0 + p_26_2;
  assign t_r27_c3_6 = t_r27_c3_1 + p_26_4;
  assign t_r27_c3_7 = t_r27_c3_2 + t_r27_c3_3;
  assign t_r27_c3_8 = t_r27_c3_4 + p_28_2;
  assign t_r27_c3_9 = t_r27_c3_5 + t_r27_c3_6;
  assign t_r27_c3_10 = t_r27_c3_7 + t_r27_c3_8;
  assign t_r27_c3_11 = t_r27_c3_9 + t_r27_c3_10;
  assign t_r27_c3_12 = t_r27_c3_11 + p_28_4;
  assign out_27_3 = t_r27_c3_12 >> 4;

  assign t_r27_c4_0 = p_26_4 << 1;
  assign t_r27_c4_1 = p_27_3 << 1;
  assign t_r27_c4_2 = p_27_4 << 2;
  assign t_r27_c4_3 = p_27_5 << 1;
  assign t_r27_c4_4 = p_28_4 << 1;
  assign t_r27_c4_5 = t_r27_c4_0 + p_26_3;
  assign t_r27_c4_6 = t_r27_c4_1 + p_26_5;
  assign t_r27_c4_7 = t_r27_c4_2 + t_r27_c4_3;
  assign t_r27_c4_8 = t_r27_c4_4 + p_28_3;
  assign t_r27_c4_9 = t_r27_c4_5 + t_r27_c4_6;
  assign t_r27_c4_10 = t_r27_c4_7 + t_r27_c4_8;
  assign t_r27_c4_11 = t_r27_c4_9 + t_r27_c4_10;
  assign t_r27_c4_12 = t_r27_c4_11 + p_28_5;
  assign out_27_4 = t_r27_c4_12 >> 4;

  assign t_r27_c5_0 = p_26_5 << 1;
  assign t_r27_c5_1 = p_27_4 << 1;
  assign t_r27_c5_2 = p_27_5 << 2;
  assign t_r27_c5_3 = p_27_6 << 1;
  assign t_r27_c5_4 = p_28_5 << 1;
  assign t_r27_c5_5 = t_r27_c5_0 + p_26_4;
  assign t_r27_c5_6 = t_r27_c5_1 + p_26_6;
  assign t_r27_c5_7 = t_r27_c5_2 + t_r27_c5_3;
  assign t_r27_c5_8 = t_r27_c5_4 + p_28_4;
  assign t_r27_c5_9 = t_r27_c5_5 + t_r27_c5_6;
  assign t_r27_c5_10 = t_r27_c5_7 + t_r27_c5_8;
  assign t_r27_c5_11 = t_r27_c5_9 + t_r27_c5_10;
  assign t_r27_c5_12 = t_r27_c5_11 + p_28_6;
  assign out_27_5 = t_r27_c5_12 >> 4;

  assign t_r27_c6_0 = p_26_6 << 1;
  assign t_r27_c6_1 = p_27_5 << 1;
  assign t_r27_c6_2 = p_27_6 << 2;
  assign t_r27_c6_3 = p_27_7 << 1;
  assign t_r27_c6_4 = p_28_6 << 1;
  assign t_r27_c6_5 = t_r27_c6_0 + p_26_5;
  assign t_r27_c6_6 = t_r27_c6_1 + p_26_7;
  assign t_r27_c6_7 = t_r27_c6_2 + t_r27_c6_3;
  assign t_r27_c6_8 = t_r27_c6_4 + p_28_5;
  assign t_r27_c6_9 = t_r27_c6_5 + t_r27_c6_6;
  assign t_r27_c6_10 = t_r27_c6_7 + t_r27_c6_8;
  assign t_r27_c6_11 = t_r27_c6_9 + t_r27_c6_10;
  assign t_r27_c6_12 = t_r27_c6_11 + p_28_7;
  assign out_27_6 = t_r27_c6_12 >> 4;

  assign t_r27_c7_0 = p_26_7 << 1;
  assign t_r27_c7_1 = p_27_6 << 1;
  assign t_r27_c7_2 = p_27_7 << 2;
  assign t_r27_c7_3 = p_27_8 << 1;
  assign t_r27_c7_4 = p_28_7 << 1;
  assign t_r27_c7_5 = t_r27_c7_0 + p_26_6;
  assign t_r27_c7_6 = t_r27_c7_1 + p_26_8;
  assign t_r27_c7_7 = t_r27_c7_2 + t_r27_c7_3;
  assign t_r27_c7_8 = t_r27_c7_4 + p_28_6;
  assign t_r27_c7_9 = t_r27_c7_5 + t_r27_c7_6;
  assign t_r27_c7_10 = t_r27_c7_7 + t_r27_c7_8;
  assign t_r27_c7_11 = t_r27_c7_9 + t_r27_c7_10;
  assign t_r27_c7_12 = t_r27_c7_11 + p_28_8;
  assign out_27_7 = t_r27_c7_12 >> 4;

  assign t_r27_c8_0 = p_26_8 << 1;
  assign t_r27_c8_1 = p_27_7 << 1;
  assign t_r27_c8_2 = p_27_8 << 2;
  assign t_r27_c8_3 = p_27_9 << 1;
  assign t_r27_c8_4 = p_28_8 << 1;
  assign t_r27_c8_5 = t_r27_c8_0 + p_26_7;
  assign t_r27_c8_6 = t_r27_c8_1 + p_26_9;
  assign t_r27_c8_7 = t_r27_c8_2 + t_r27_c8_3;
  assign t_r27_c8_8 = t_r27_c8_4 + p_28_7;
  assign t_r27_c8_9 = t_r27_c8_5 + t_r27_c8_6;
  assign t_r27_c8_10 = t_r27_c8_7 + t_r27_c8_8;
  assign t_r27_c8_11 = t_r27_c8_9 + t_r27_c8_10;
  assign t_r27_c8_12 = t_r27_c8_11 + p_28_9;
  assign out_27_8 = t_r27_c8_12 >> 4;

  assign t_r27_c9_0 = p_26_9 << 1;
  assign t_r27_c9_1 = p_27_8 << 1;
  assign t_r27_c9_2 = p_27_9 << 2;
  assign t_r27_c9_3 = p_27_10 << 1;
  assign t_r27_c9_4 = p_28_9 << 1;
  assign t_r27_c9_5 = t_r27_c9_0 + p_26_8;
  assign t_r27_c9_6 = t_r27_c9_1 + p_26_10;
  assign t_r27_c9_7 = t_r27_c9_2 + t_r27_c9_3;
  assign t_r27_c9_8 = t_r27_c9_4 + p_28_8;
  assign t_r27_c9_9 = t_r27_c9_5 + t_r27_c9_6;
  assign t_r27_c9_10 = t_r27_c9_7 + t_r27_c9_8;
  assign t_r27_c9_11 = t_r27_c9_9 + t_r27_c9_10;
  assign t_r27_c9_12 = t_r27_c9_11 + p_28_10;
  assign out_27_9 = t_r27_c9_12 >> 4;

  assign t_r27_c10_0 = p_26_10 << 1;
  assign t_r27_c10_1 = p_27_9 << 1;
  assign t_r27_c10_2 = p_27_10 << 2;
  assign t_r27_c10_3 = p_27_11 << 1;
  assign t_r27_c10_4 = p_28_10 << 1;
  assign t_r27_c10_5 = t_r27_c10_0 + p_26_9;
  assign t_r27_c10_6 = t_r27_c10_1 + p_26_11;
  assign t_r27_c10_7 = t_r27_c10_2 + t_r27_c10_3;
  assign t_r27_c10_8 = t_r27_c10_4 + p_28_9;
  assign t_r27_c10_9 = t_r27_c10_5 + t_r27_c10_6;
  assign t_r27_c10_10 = t_r27_c10_7 + t_r27_c10_8;
  assign t_r27_c10_11 = t_r27_c10_9 + t_r27_c10_10;
  assign t_r27_c10_12 = t_r27_c10_11 + p_28_11;
  assign out_27_10 = t_r27_c10_12 >> 4;

  assign t_r27_c11_0 = p_26_11 << 1;
  assign t_r27_c11_1 = p_27_10 << 1;
  assign t_r27_c11_2 = p_27_11 << 2;
  assign t_r27_c11_3 = p_27_12 << 1;
  assign t_r27_c11_4 = p_28_11 << 1;
  assign t_r27_c11_5 = t_r27_c11_0 + p_26_10;
  assign t_r27_c11_6 = t_r27_c11_1 + p_26_12;
  assign t_r27_c11_7 = t_r27_c11_2 + t_r27_c11_3;
  assign t_r27_c11_8 = t_r27_c11_4 + p_28_10;
  assign t_r27_c11_9 = t_r27_c11_5 + t_r27_c11_6;
  assign t_r27_c11_10 = t_r27_c11_7 + t_r27_c11_8;
  assign t_r27_c11_11 = t_r27_c11_9 + t_r27_c11_10;
  assign t_r27_c11_12 = t_r27_c11_11 + p_28_12;
  assign out_27_11 = t_r27_c11_12 >> 4;

  assign t_r27_c12_0 = p_26_12 << 1;
  assign t_r27_c12_1 = p_27_11 << 1;
  assign t_r27_c12_2 = p_27_12 << 2;
  assign t_r27_c12_3 = p_27_13 << 1;
  assign t_r27_c12_4 = p_28_12 << 1;
  assign t_r27_c12_5 = t_r27_c12_0 + p_26_11;
  assign t_r27_c12_6 = t_r27_c12_1 + p_26_13;
  assign t_r27_c12_7 = t_r27_c12_2 + t_r27_c12_3;
  assign t_r27_c12_8 = t_r27_c12_4 + p_28_11;
  assign t_r27_c12_9 = t_r27_c12_5 + t_r27_c12_6;
  assign t_r27_c12_10 = t_r27_c12_7 + t_r27_c12_8;
  assign t_r27_c12_11 = t_r27_c12_9 + t_r27_c12_10;
  assign t_r27_c12_12 = t_r27_c12_11 + p_28_13;
  assign out_27_12 = t_r27_c12_12 >> 4;

  assign t_r27_c13_0 = p_26_13 << 1;
  assign t_r27_c13_1 = p_27_12 << 1;
  assign t_r27_c13_2 = p_27_13 << 2;
  assign t_r27_c13_3 = p_27_14 << 1;
  assign t_r27_c13_4 = p_28_13 << 1;
  assign t_r27_c13_5 = t_r27_c13_0 + p_26_12;
  assign t_r27_c13_6 = t_r27_c13_1 + p_26_14;
  assign t_r27_c13_7 = t_r27_c13_2 + t_r27_c13_3;
  assign t_r27_c13_8 = t_r27_c13_4 + p_28_12;
  assign t_r27_c13_9 = t_r27_c13_5 + t_r27_c13_6;
  assign t_r27_c13_10 = t_r27_c13_7 + t_r27_c13_8;
  assign t_r27_c13_11 = t_r27_c13_9 + t_r27_c13_10;
  assign t_r27_c13_12 = t_r27_c13_11 + p_28_14;
  assign out_27_13 = t_r27_c13_12 >> 4;

  assign t_r27_c14_0 = p_26_14 << 1;
  assign t_r27_c14_1 = p_27_13 << 1;
  assign t_r27_c14_2 = p_27_14 << 2;
  assign t_r27_c14_3 = p_27_15 << 1;
  assign t_r27_c14_4 = p_28_14 << 1;
  assign t_r27_c14_5 = t_r27_c14_0 + p_26_13;
  assign t_r27_c14_6 = t_r27_c14_1 + p_26_15;
  assign t_r27_c14_7 = t_r27_c14_2 + t_r27_c14_3;
  assign t_r27_c14_8 = t_r27_c14_4 + p_28_13;
  assign t_r27_c14_9 = t_r27_c14_5 + t_r27_c14_6;
  assign t_r27_c14_10 = t_r27_c14_7 + t_r27_c14_8;
  assign t_r27_c14_11 = t_r27_c14_9 + t_r27_c14_10;
  assign t_r27_c14_12 = t_r27_c14_11 + p_28_15;
  assign out_27_14 = t_r27_c14_12 >> 4;

  assign t_r27_c15_0 = p_26_15 << 1;
  assign t_r27_c15_1 = p_27_14 << 1;
  assign t_r27_c15_2 = p_27_15 << 2;
  assign t_r27_c15_3 = p_27_16 << 1;
  assign t_r27_c15_4 = p_28_15 << 1;
  assign t_r27_c15_5 = t_r27_c15_0 + p_26_14;
  assign t_r27_c15_6 = t_r27_c15_1 + p_26_16;
  assign t_r27_c15_7 = t_r27_c15_2 + t_r27_c15_3;
  assign t_r27_c15_8 = t_r27_c15_4 + p_28_14;
  assign t_r27_c15_9 = t_r27_c15_5 + t_r27_c15_6;
  assign t_r27_c15_10 = t_r27_c15_7 + t_r27_c15_8;
  assign t_r27_c15_11 = t_r27_c15_9 + t_r27_c15_10;
  assign t_r27_c15_12 = t_r27_c15_11 + p_28_16;
  assign out_27_15 = t_r27_c15_12 >> 4;

  assign t_r27_c16_0 = p_26_16 << 1;
  assign t_r27_c16_1 = p_27_15 << 1;
  assign t_r27_c16_2 = p_27_16 << 2;
  assign t_r27_c16_3 = p_27_17 << 1;
  assign t_r27_c16_4 = p_28_16 << 1;
  assign t_r27_c16_5 = t_r27_c16_0 + p_26_15;
  assign t_r27_c16_6 = t_r27_c16_1 + p_26_17;
  assign t_r27_c16_7 = t_r27_c16_2 + t_r27_c16_3;
  assign t_r27_c16_8 = t_r27_c16_4 + p_28_15;
  assign t_r27_c16_9 = t_r27_c16_5 + t_r27_c16_6;
  assign t_r27_c16_10 = t_r27_c16_7 + t_r27_c16_8;
  assign t_r27_c16_11 = t_r27_c16_9 + t_r27_c16_10;
  assign t_r27_c16_12 = t_r27_c16_11 + p_28_17;
  assign out_27_16 = t_r27_c16_12 >> 4;

  assign t_r27_c17_0 = p_26_17 << 1;
  assign t_r27_c17_1 = p_27_16 << 1;
  assign t_r27_c17_2 = p_27_17 << 2;
  assign t_r27_c17_3 = p_27_18 << 1;
  assign t_r27_c17_4 = p_28_17 << 1;
  assign t_r27_c17_5 = t_r27_c17_0 + p_26_16;
  assign t_r27_c17_6 = t_r27_c17_1 + p_26_18;
  assign t_r27_c17_7 = t_r27_c17_2 + t_r27_c17_3;
  assign t_r27_c17_8 = t_r27_c17_4 + p_28_16;
  assign t_r27_c17_9 = t_r27_c17_5 + t_r27_c17_6;
  assign t_r27_c17_10 = t_r27_c17_7 + t_r27_c17_8;
  assign t_r27_c17_11 = t_r27_c17_9 + t_r27_c17_10;
  assign t_r27_c17_12 = t_r27_c17_11 + p_28_18;
  assign out_27_17 = t_r27_c17_12 >> 4;

  assign t_r27_c18_0 = p_26_18 << 1;
  assign t_r27_c18_1 = p_27_17 << 1;
  assign t_r27_c18_2 = p_27_18 << 2;
  assign t_r27_c18_3 = p_27_19 << 1;
  assign t_r27_c18_4 = p_28_18 << 1;
  assign t_r27_c18_5 = t_r27_c18_0 + p_26_17;
  assign t_r27_c18_6 = t_r27_c18_1 + p_26_19;
  assign t_r27_c18_7 = t_r27_c18_2 + t_r27_c18_3;
  assign t_r27_c18_8 = t_r27_c18_4 + p_28_17;
  assign t_r27_c18_9 = t_r27_c18_5 + t_r27_c18_6;
  assign t_r27_c18_10 = t_r27_c18_7 + t_r27_c18_8;
  assign t_r27_c18_11 = t_r27_c18_9 + t_r27_c18_10;
  assign t_r27_c18_12 = t_r27_c18_11 + p_28_19;
  assign out_27_18 = t_r27_c18_12 >> 4;

  assign t_r27_c19_0 = p_26_19 << 1;
  assign t_r27_c19_1 = p_27_18 << 1;
  assign t_r27_c19_2 = p_27_19 << 2;
  assign t_r27_c19_3 = p_27_20 << 1;
  assign t_r27_c19_4 = p_28_19 << 1;
  assign t_r27_c19_5 = t_r27_c19_0 + p_26_18;
  assign t_r27_c19_6 = t_r27_c19_1 + p_26_20;
  assign t_r27_c19_7 = t_r27_c19_2 + t_r27_c19_3;
  assign t_r27_c19_8 = t_r27_c19_4 + p_28_18;
  assign t_r27_c19_9 = t_r27_c19_5 + t_r27_c19_6;
  assign t_r27_c19_10 = t_r27_c19_7 + t_r27_c19_8;
  assign t_r27_c19_11 = t_r27_c19_9 + t_r27_c19_10;
  assign t_r27_c19_12 = t_r27_c19_11 + p_28_20;
  assign out_27_19 = t_r27_c19_12 >> 4;

  assign t_r27_c20_0 = p_26_20 << 1;
  assign t_r27_c20_1 = p_27_19 << 1;
  assign t_r27_c20_2 = p_27_20 << 2;
  assign t_r27_c20_3 = p_27_21 << 1;
  assign t_r27_c20_4 = p_28_20 << 1;
  assign t_r27_c20_5 = t_r27_c20_0 + p_26_19;
  assign t_r27_c20_6 = t_r27_c20_1 + p_26_21;
  assign t_r27_c20_7 = t_r27_c20_2 + t_r27_c20_3;
  assign t_r27_c20_8 = t_r27_c20_4 + p_28_19;
  assign t_r27_c20_9 = t_r27_c20_5 + t_r27_c20_6;
  assign t_r27_c20_10 = t_r27_c20_7 + t_r27_c20_8;
  assign t_r27_c20_11 = t_r27_c20_9 + t_r27_c20_10;
  assign t_r27_c20_12 = t_r27_c20_11 + p_28_21;
  assign out_27_20 = t_r27_c20_12 >> 4;

  assign t_r27_c21_0 = p_26_21 << 1;
  assign t_r27_c21_1 = p_27_20 << 1;
  assign t_r27_c21_2 = p_27_21 << 2;
  assign t_r27_c21_3 = p_27_22 << 1;
  assign t_r27_c21_4 = p_28_21 << 1;
  assign t_r27_c21_5 = t_r27_c21_0 + p_26_20;
  assign t_r27_c21_6 = t_r27_c21_1 + p_26_22;
  assign t_r27_c21_7 = t_r27_c21_2 + t_r27_c21_3;
  assign t_r27_c21_8 = t_r27_c21_4 + p_28_20;
  assign t_r27_c21_9 = t_r27_c21_5 + t_r27_c21_6;
  assign t_r27_c21_10 = t_r27_c21_7 + t_r27_c21_8;
  assign t_r27_c21_11 = t_r27_c21_9 + t_r27_c21_10;
  assign t_r27_c21_12 = t_r27_c21_11 + p_28_22;
  assign out_27_21 = t_r27_c21_12 >> 4;

  assign t_r27_c22_0 = p_26_22 << 1;
  assign t_r27_c22_1 = p_27_21 << 1;
  assign t_r27_c22_2 = p_27_22 << 2;
  assign t_r27_c22_3 = p_27_23 << 1;
  assign t_r27_c22_4 = p_28_22 << 1;
  assign t_r27_c22_5 = t_r27_c22_0 + p_26_21;
  assign t_r27_c22_6 = t_r27_c22_1 + p_26_23;
  assign t_r27_c22_7 = t_r27_c22_2 + t_r27_c22_3;
  assign t_r27_c22_8 = t_r27_c22_4 + p_28_21;
  assign t_r27_c22_9 = t_r27_c22_5 + t_r27_c22_6;
  assign t_r27_c22_10 = t_r27_c22_7 + t_r27_c22_8;
  assign t_r27_c22_11 = t_r27_c22_9 + t_r27_c22_10;
  assign t_r27_c22_12 = t_r27_c22_11 + p_28_23;
  assign out_27_22 = t_r27_c22_12 >> 4;

  assign t_r27_c23_0 = p_26_23 << 1;
  assign t_r27_c23_1 = p_27_22 << 1;
  assign t_r27_c23_2 = p_27_23 << 2;
  assign t_r27_c23_3 = p_27_24 << 1;
  assign t_r27_c23_4 = p_28_23 << 1;
  assign t_r27_c23_5 = t_r27_c23_0 + p_26_22;
  assign t_r27_c23_6 = t_r27_c23_1 + p_26_24;
  assign t_r27_c23_7 = t_r27_c23_2 + t_r27_c23_3;
  assign t_r27_c23_8 = t_r27_c23_4 + p_28_22;
  assign t_r27_c23_9 = t_r27_c23_5 + t_r27_c23_6;
  assign t_r27_c23_10 = t_r27_c23_7 + t_r27_c23_8;
  assign t_r27_c23_11 = t_r27_c23_9 + t_r27_c23_10;
  assign t_r27_c23_12 = t_r27_c23_11 + p_28_24;
  assign out_27_23 = t_r27_c23_12 >> 4;

  assign t_r27_c24_0 = p_26_24 << 1;
  assign t_r27_c24_1 = p_27_23 << 1;
  assign t_r27_c24_2 = p_27_24 << 2;
  assign t_r27_c24_3 = p_27_25 << 1;
  assign t_r27_c24_4 = p_28_24 << 1;
  assign t_r27_c24_5 = t_r27_c24_0 + p_26_23;
  assign t_r27_c24_6 = t_r27_c24_1 + p_26_25;
  assign t_r27_c24_7 = t_r27_c24_2 + t_r27_c24_3;
  assign t_r27_c24_8 = t_r27_c24_4 + p_28_23;
  assign t_r27_c24_9 = t_r27_c24_5 + t_r27_c24_6;
  assign t_r27_c24_10 = t_r27_c24_7 + t_r27_c24_8;
  assign t_r27_c24_11 = t_r27_c24_9 + t_r27_c24_10;
  assign t_r27_c24_12 = t_r27_c24_11 + p_28_25;
  assign out_27_24 = t_r27_c24_12 >> 4;

  assign t_r27_c25_0 = p_26_25 << 1;
  assign t_r27_c25_1 = p_27_24 << 1;
  assign t_r27_c25_2 = p_27_25 << 2;
  assign t_r27_c25_3 = p_27_26 << 1;
  assign t_r27_c25_4 = p_28_25 << 1;
  assign t_r27_c25_5 = t_r27_c25_0 + p_26_24;
  assign t_r27_c25_6 = t_r27_c25_1 + p_26_26;
  assign t_r27_c25_7 = t_r27_c25_2 + t_r27_c25_3;
  assign t_r27_c25_8 = t_r27_c25_4 + p_28_24;
  assign t_r27_c25_9 = t_r27_c25_5 + t_r27_c25_6;
  assign t_r27_c25_10 = t_r27_c25_7 + t_r27_c25_8;
  assign t_r27_c25_11 = t_r27_c25_9 + t_r27_c25_10;
  assign t_r27_c25_12 = t_r27_c25_11 + p_28_26;
  assign out_27_25 = t_r27_c25_12 >> 4;

  assign t_r27_c26_0 = p_26_26 << 1;
  assign t_r27_c26_1 = p_27_25 << 1;
  assign t_r27_c26_2 = p_27_26 << 2;
  assign t_r27_c26_3 = p_27_27 << 1;
  assign t_r27_c26_4 = p_28_26 << 1;
  assign t_r27_c26_5 = t_r27_c26_0 + p_26_25;
  assign t_r27_c26_6 = t_r27_c26_1 + p_26_27;
  assign t_r27_c26_7 = t_r27_c26_2 + t_r27_c26_3;
  assign t_r27_c26_8 = t_r27_c26_4 + p_28_25;
  assign t_r27_c26_9 = t_r27_c26_5 + t_r27_c26_6;
  assign t_r27_c26_10 = t_r27_c26_7 + t_r27_c26_8;
  assign t_r27_c26_11 = t_r27_c26_9 + t_r27_c26_10;
  assign t_r27_c26_12 = t_r27_c26_11 + p_28_27;
  assign out_27_26 = t_r27_c26_12 >> 4;

  assign t_r27_c27_0 = p_26_27 << 1;
  assign t_r27_c27_1 = p_27_26 << 1;
  assign t_r27_c27_2 = p_27_27 << 2;
  assign t_r27_c27_3 = p_27_28 << 1;
  assign t_r27_c27_4 = p_28_27 << 1;
  assign t_r27_c27_5 = t_r27_c27_0 + p_26_26;
  assign t_r27_c27_6 = t_r27_c27_1 + p_26_28;
  assign t_r27_c27_7 = t_r27_c27_2 + t_r27_c27_3;
  assign t_r27_c27_8 = t_r27_c27_4 + p_28_26;
  assign t_r27_c27_9 = t_r27_c27_5 + t_r27_c27_6;
  assign t_r27_c27_10 = t_r27_c27_7 + t_r27_c27_8;
  assign t_r27_c27_11 = t_r27_c27_9 + t_r27_c27_10;
  assign t_r27_c27_12 = t_r27_c27_11 + p_28_28;
  assign out_27_27 = t_r27_c27_12 >> 4;

  assign t_r27_c28_0 = p_26_28 << 1;
  assign t_r27_c28_1 = p_27_27 << 1;
  assign t_r27_c28_2 = p_27_28 << 2;
  assign t_r27_c28_3 = p_27_29 << 1;
  assign t_r27_c28_4 = p_28_28 << 1;
  assign t_r27_c28_5 = t_r27_c28_0 + p_26_27;
  assign t_r27_c28_6 = t_r27_c28_1 + p_26_29;
  assign t_r27_c28_7 = t_r27_c28_2 + t_r27_c28_3;
  assign t_r27_c28_8 = t_r27_c28_4 + p_28_27;
  assign t_r27_c28_9 = t_r27_c28_5 + t_r27_c28_6;
  assign t_r27_c28_10 = t_r27_c28_7 + t_r27_c28_8;
  assign t_r27_c28_11 = t_r27_c28_9 + t_r27_c28_10;
  assign t_r27_c28_12 = t_r27_c28_11 + p_28_29;
  assign out_27_28 = t_r27_c28_12 >> 4;

  assign t_r27_c29_0 = p_26_29 << 1;
  assign t_r27_c29_1 = p_27_28 << 1;
  assign t_r27_c29_2 = p_27_29 << 2;
  assign t_r27_c29_3 = p_27_30 << 1;
  assign t_r27_c29_4 = p_28_29 << 1;
  assign t_r27_c29_5 = t_r27_c29_0 + p_26_28;
  assign t_r27_c29_6 = t_r27_c29_1 + p_26_30;
  assign t_r27_c29_7 = t_r27_c29_2 + t_r27_c29_3;
  assign t_r27_c29_8 = t_r27_c29_4 + p_28_28;
  assign t_r27_c29_9 = t_r27_c29_5 + t_r27_c29_6;
  assign t_r27_c29_10 = t_r27_c29_7 + t_r27_c29_8;
  assign t_r27_c29_11 = t_r27_c29_9 + t_r27_c29_10;
  assign t_r27_c29_12 = t_r27_c29_11 + p_28_30;
  assign out_27_29 = t_r27_c29_12 >> 4;

  assign t_r27_c30_0 = p_26_30 << 1;
  assign t_r27_c30_1 = p_27_29 << 1;
  assign t_r27_c30_2 = p_27_30 << 2;
  assign t_r27_c30_3 = p_27_31 << 1;
  assign t_r27_c30_4 = p_28_30 << 1;
  assign t_r27_c30_5 = t_r27_c30_0 + p_26_29;
  assign t_r27_c30_6 = t_r27_c30_1 + p_26_31;
  assign t_r27_c30_7 = t_r27_c30_2 + t_r27_c30_3;
  assign t_r27_c30_8 = t_r27_c30_4 + p_28_29;
  assign t_r27_c30_9 = t_r27_c30_5 + t_r27_c30_6;
  assign t_r27_c30_10 = t_r27_c30_7 + t_r27_c30_8;
  assign t_r27_c30_11 = t_r27_c30_9 + t_r27_c30_10;
  assign t_r27_c30_12 = t_r27_c30_11 + p_28_31;
  assign out_27_30 = t_r27_c30_12 >> 4;

  assign t_r27_c31_0 = p_26_31 << 1;
  assign t_r27_c31_1 = p_27_30 << 1;
  assign t_r27_c31_2 = p_27_31 << 2;
  assign t_r27_c31_3 = p_27_32 << 1;
  assign t_r27_c31_4 = p_28_31 << 1;
  assign t_r27_c31_5 = t_r27_c31_0 + p_26_30;
  assign t_r27_c31_6 = t_r27_c31_1 + p_26_32;
  assign t_r27_c31_7 = t_r27_c31_2 + t_r27_c31_3;
  assign t_r27_c31_8 = t_r27_c31_4 + p_28_30;
  assign t_r27_c31_9 = t_r27_c31_5 + t_r27_c31_6;
  assign t_r27_c31_10 = t_r27_c31_7 + t_r27_c31_8;
  assign t_r27_c31_11 = t_r27_c31_9 + t_r27_c31_10;
  assign t_r27_c31_12 = t_r27_c31_11 + p_28_32;
  assign out_27_31 = t_r27_c31_12 >> 4;

  assign t_r27_c32_0 = p_26_32 << 1;
  assign t_r27_c32_1 = p_27_31 << 1;
  assign t_r27_c32_2 = p_27_32 << 2;
  assign t_r27_c32_3 = p_27_33 << 1;
  assign t_r27_c32_4 = p_28_32 << 1;
  assign t_r27_c32_5 = t_r27_c32_0 + p_26_31;
  assign t_r27_c32_6 = t_r27_c32_1 + p_26_33;
  assign t_r27_c32_7 = t_r27_c32_2 + t_r27_c32_3;
  assign t_r27_c32_8 = t_r27_c32_4 + p_28_31;
  assign t_r27_c32_9 = t_r27_c32_5 + t_r27_c32_6;
  assign t_r27_c32_10 = t_r27_c32_7 + t_r27_c32_8;
  assign t_r27_c32_11 = t_r27_c32_9 + t_r27_c32_10;
  assign t_r27_c32_12 = t_r27_c32_11 + p_28_33;
  assign out_27_32 = t_r27_c32_12 >> 4;

  assign t_r27_c33_0 = p_26_33 << 1;
  assign t_r27_c33_1 = p_27_32 << 1;
  assign t_r27_c33_2 = p_27_33 << 2;
  assign t_r27_c33_3 = p_27_34 << 1;
  assign t_r27_c33_4 = p_28_33 << 1;
  assign t_r27_c33_5 = t_r27_c33_0 + p_26_32;
  assign t_r27_c33_6 = t_r27_c33_1 + p_26_34;
  assign t_r27_c33_7 = t_r27_c33_2 + t_r27_c33_3;
  assign t_r27_c33_8 = t_r27_c33_4 + p_28_32;
  assign t_r27_c33_9 = t_r27_c33_5 + t_r27_c33_6;
  assign t_r27_c33_10 = t_r27_c33_7 + t_r27_c33_8;
  assign t_r27_c33_11 = t_r27_c33_9 + t_r27_c33_10;
  assign t_r27_c33_12 = t_r27_c33_11 + p_28_34;
  assign out_27_33 = t_r27_c33_12 >> 4;

  assign t_r27_c34_0 = p_26_34 << 1;
  assign t_r27_c34_1 = p_27_33 << 1;
  assign t_r27_c34_2 = p_27_34 << 2;
  assign t_r27_c34_3 = p_27_35 << 1;
  assign t_r27_c34_4 = p_28_34 << 1;
  assign t_r27_c34_5 = t_r27_c34_0 + p_26_33;
  assign t_r27_c34_6 = t_r27_c34_1 + p_26_35;
  assign t_r27_c34_7 = t_r27_c34_2 + t_r27_c34_3;
  assign t_r27_c34_8 = t_r27_c34_4 + p_28_33;
  assign t_r27_c34_9 = t_r27_c34_5 + t_r27_c34_6;
  assign t_r27_c34_10 = t_r27_c34_7 + t_r27_c34_8;
  assign t_r27_c34_11 = t_r27_c34_9 + t_r27_c34_10;
  assign t_r27_c34_12 = t_r27_c34_11 + p_28_35;
  assign out_27_34 = t_r27_c34_12 >> 4;

  assign t_r27_c35_0 = p_26_35 << 1;
  assign t_r27_c35_1 = p_27_34 << 1;
  assign t_r27_c35_2 = p_27_35 << 2;
  assign t_r27_c35_3 = p_27_36 << 1;
  assign t_r27_c35_4 = p_28_35 << 1;
  assign t_r27_c35_5 = t_r27_c35_0 + p_26_34;
  assign t_r27_c35_6 = t_r27_c35_1 + p_26_36;
  assign t_r27_c35_7 = t_r27_c35_2 + t_r27_c35_3;
  assign t_r27_c35_8 = t_r27_c35_4 + p_28_34;
  assign t_r27_c35_9 = t_r27_c35_5 + t_r27_c35_6;
  assign t_r27_c35_10 = t_r27_c35_7 + t_r27_c35_8;
  assign t_r27_c35_11 = t_r27_c35_9 + t_r27_c35_10;
  assign t_r27_c35_12 = t_r27_c35_11 + p_28_36;
  assign out_27_35 = t_r27_c35_12 >> 4;

  assign t_r27_c36_0 = p_26_36 << 1;
  assign t_r27_c36_1 = p_27_35 << 1;
  assign t_r27_c36_2 = p_27_36 << 2;
  assign t_r27_c36_3 = p_27_37 << 1;
  assign t_r27_c36_4 = p_28_36 << 1;
  assign t_r27_c36_5 = t_r27_c36_0 + p_26_35;
  assign t_r27_c36_6 = t_r27_c36_1 + p_26_37;
  assign t_r27_c36_7 = t_r27_c36_2 + t_r27_c36_3;
  assign t_r27_c36_8 = t_r27_c36_4 + p_28_35;
  assign t_r27_c36_9 = t_r27_c36_5 + t_r27_c36_6;
  assign t_r27_c36_10 = t_r27_c36_7 + t_r27_c36_8;
  assign t_r27_c36_11 = t_r27_c36_9 + t_r27_c36_10;
  assign t_r27_c36_12 = t_r27_c36_11 + p_28_37;
  assign out_27_36 = t_r27_c36_12 >> 4;

  assign t_r27_c37_0 = p_26_37 << 1;
  assign t_r27_c37_1 = p_27_36 << 1;
  assign t_r27_c37_2 = p_27_37 << 2;
  assign t_r27_c37_3 = p_27_38 << 1;
  assign t_r27_c37_4 = p_28_37 << 1;
  assign t_r27_c37_5 = t_r27_c37_0 + p_26_36;
  assign t_r27_c37_6 = t_r27_c37_1 + p_26_38;
  assign t_r27_c37_7 = t_r27_c37_2 + t_r27_c37_3;
  assign t_r27_c37_8 = t_r27_c37_4 + p_28_36;
  assign t_r27_c37_9 = t_r27_c37_5 + t_r27_c37_6;
  assign t_r27_c37_10 = t_r27_c37_7 + t_r27_c37_8;
  assign t_r27_c37_11 = t_r27_c37_9 + t_r27_c37_10;
  assign t_r27_c37_12 = t_r27_c37_11 + p_28_38;
  assign out_27_37 = t_r27_c37_12 >> 4;

  assign t_r27_c38_0 = p_26_38 << 1;
  assign t_r27_c38_1 = p_27_37 << 1;
  assign t_r27_c38_2 = p_27_38 << 2;
  assign t_r27_c38_3 = p_27_39 << 1;
  assign t_r27_c38_4 = p_28_38 << 1;
  assign t_r27_c38_5 = t_r27_c38_0 + p_26_37;
  assign t_r27_c38_6 = t_r27_c38_1 + p_26_39;
  assign t_r27_c38_7 = t_r27_c38_2 + t_r27_c38_3;
  assign t_r27_c38_8 = t_r27_c38_4 + p_28_37;
  assign t_r27_c38_9 = t_r27_c38_5 + t_r27_c38_6;
  assign t_r27_c38_10 = t_r27_c38_7 + t_r27_c38_8;
  assign t_r27_c38_11 = t_r27_c38_9 + t_r27_c38_10;
  assign t_r27_c38_12 = t_r27_c38_11 + p_28_39;
  assign out_27_38 = t_r27_c38_12 >> 4;

  assign t_r27_c39_0 = p_26_39 << 1;
  assign t_r27_c39_1 = p_27_38 << 1;
  assign t_r27_c39_2 = p_27_39 << 2;
  assign t_r27_c39_3 = p_27_40 << 1;
  assign t_r27_c39_4 = p_28_39 << 1;
  assign t_r27_c39_5 = t_r27_c39_0 + p_26_38;
  assign t_r27_c39_6 = t_r27_c39_1 + p_26_40;
  assign t_r27_c39_7 = t_r27_c39_2 + t_r27_c39_3;
  assign t_r27_c39_8 = t_r27_c39_4 + p_28_38;
  assign t_r27_c39_9 = t_r27_c39_5 + t_r27_c39_6;
  assign t_r27_c39_10 = t_r27_c39_7 + t_r27_c39_8;
  assign t_r27_c39_11 = t_r27_c39_9 + t_r27_c39_10;
  assign t_r27_c39_12 = t_r27_c39_11 + p_28_40;
  assign out_27_39 = t_r27_c39_12 >> 4;

  assign t_r27_c40_0 = p_26_40 << 1;
  assign t_r27_c40_1 = p_27_39 << 1;
  assign t_r27_c40_2 = p_27_40 << 2;
  assign t_r27_c40_3 = p_27_41 << 1;
  assign t_r27_c40_4 = p_28_40 << 1;
  assign t_r27_c40_5 = t_r27_c40_0 + p_26_39;
  assign t_r27_c40_6 = t_r27_c40_1 + p_26_41;
  assign t_r27_c40_7 = t_r27_c40_2 + t_r27_c40_3;
  assign t_r27_c40_8 = t_r27_c40_4 + p_28_39;
  assign t_r27_c40_9 = t_r27_c40_5 + t_r27_c40_6;
  assign t_r27_c40_10 = t_r27_c40_7 + t_r27_c40_8;
  assign t_r27_c40_11 = t_r27_c40_9 + t_r27_c40_10;
  assign t_r27_c40_12 = t_r27_c40_11 + p_28_41;
  assign out_27_40 = t_r27_c40_12 >> 4;

  assign t_r27_c41_0 = p_26_41 << 1;
  assign t_r27_c41_1 = p_27_40 << 1;
  assign t_r27_c41_2 = p_27_41 << 2;
  assign t_r27_c41_3 = p_27_42 << 1;
  assign t_r27_c41_4 = p_28_41 << 1;
  assign t_r27_c41_5 = t_r27_c41_0 + p_26_40;
  assign t_r27_c41_6 = t_r27_c41_1 + p_26_42;
  assign t_r27_c41_7 = t_r27_c41_2 + t_r27_c41_3;
  assign t_r27_c41_8 = t_r27_c41_4 + p_28_40;
  assign t_r27_c41_9 = t_r27_c41_5 + t_r27_c41_6;
  assign t_r27_c41_10 = t_r27_c41_7 + t_r27_c41_8;
  assign t_r27_c41_11 = t_r27_c41_9 + t_r27_c41_10;
  assign t_r27_c41_12 = t_r27_c41_11 + p_28_42;
  assign out_27_41 = t_r27_c41_12 >> 4;

  assign t_r27_c42_0 = p_26_42 << 1;
  assign t_r27_c42_1 = p_27_41 << 1;
  assign t_r27_c42_2 = p_27_42 << 2;
  assign t_r27_c42_3 = p_27_43 << 1;
  assign t_r27_c42_4 = p_28_42 << 1;
  assign t_r27_c42_5 = t_r27_c42_0 + p_26_41;
  assign t_r27_c42_6 = t_r27_c42_1 + p_26_43;
  assign t_r27_c42_7 = t_r27_c42_2 + t_r27_c42_3;
  assign t_r27_c42_8 = t_r27_c42_4 + p_28_41;
  assign t_r27_c42_9 = t_r27_c42_5 + t_r27_c42_6;
  assign t_r27_c42_10 = t_r27_c42_7 + t_r27_c42_8;
  assign t_r27_c42_11 = t_r27_c42_9 + t_r27_c42_10;
  assign t_r27_c42_12 = t_r27_c42_11 + p_28_43;
  assign out_27_42 = t_r27_c42_12 >> 4;

  assign t_r27_c43_0 = p_26_43 << 1;
  assign t_r27_c43_1 = p_27_42 << 1;
  assign t_r27_c43_2 = p_27_43 << 2;
  assign t_r27_c43_3 = p_27_44 << 1;
  assign t_r27_c43_4 = p_28_43 << 1;
  assign t_r27_c43_5 = t_r27_c43_0 + p_26_42;
  assign t_r27_c43_6 = t_r27_c43_1 + p_26_44;
  assign t_r27_c43_7 = t_r27_c43_2 + t_r27_c43_3;
  assign t_r27_c43_8 = t_r27_c43_4 + p_28_42;
  assign t_r27_c43_9 = t_r27_c43_5 + t_r27_c43_6;
  assign t_r27_c43_10 = t_r27_c43_7 + t_r27_c43_8;
  assign t_r27_c43_11 = t_r27_c43_9 + t_r27_c43_10;
  assign t_r27_c43_12 = t_r27_c43_11 + p_28_44;
  assign out_27_43 = t_r27_c43_12 >> 4;

  assign t_r27_c44_0 = p_26_44 << 1;
  assign t_r27_c44_1 = p_27_43 << 1;
  assign t_r27_c44_2 = p_27_44 << 2;
  assign t_r27_c44_3 = p_27_45 << 1;
  assign t_r27_c44_4 = p_28_44 << 1;
  assign t_r27_c44_5 = t_r27_c44_0 + p_26_43;
  assign t_r27_c44_6 = t_r27_c44_1 + p_26_45;
  assign t_r27_c44_7 = t_r27_c44_2 + t_r27_c44_3;
  assign t_r27_c44_8 = t_r27_c44_4 + p_28_43;
  assign t_r27_c44_9 = t_r27_c44_5 + t_r27_c44_6;
  assign t_r27_c44_10 = t_r27_c44_7 + t_r27_c44_8;
  assign t_r27_c44_11 = t_r27_c44_9 + t_r27_c44_10;
  assign t_r27_c44_12 = t_r27_c44_11 + p_28_45;
  assign out_27_44 = t_r27_c44_12 >> 4;

  assign t_r27_c45_0 = p_26_45 << 1;
  assign t_r27_c45_1 = p_27_44 << 1;
  assign t_r27_c45_2 = p_27_45 << 2;
  assign t_r27_c45_3 = p_27_46 << 1;
  assign t_r27_c45_4 = p_28_45 << 1;
  assign t_r27_c45_5 = t_r27_c45_0 + p_26_44;
  assign t_r27_c45_6 = t_r27_c45_1 + p_26_46;
  assign t_r27_c45_7 = t_r27_c45_2 + t_r27_c45_3;
  assign t_r27_c45_8 = t_r27_c45_4 + p_28_44;
  assign t_r27_c45_9 = t_r27_c45_5 + t_r27_c45_6;
  assign t_r27_c45_10 = t_r27_c45_7 + t_r27_c45_8;
  assign t_r27_c45_11 = t_r27_c45_9 + t_r27_c45_10;
  assign t_r27_c45_12 = t_r27_c45_11 + p_28_46;
  assign out_27_45 = t_r27_c45_12 >> 4;

  assign t_r27_c46_0 = p_26_46 << 1;
  assign t_r27_c46_1 = p_27_45 << 1;
  assign t_r27_c46_2 = p_27_46 << 2;
  assign t_r27_c46_3 = p_27_47 << 1;
  assign t_r27_c46_4 = p_28_46 << 1;
  assign t_r27_c46_5 = t_r27_c46_0 + p_26_45;
  assign t_r27_c46_6 = t_r27_c46_1 + p_26_47;
  assign t_r27_c46_7 = t_r27_c46_2 + t_r27_c46_3;
  assign t_r27_c46_8 = t_r27_c46_4 + p_28_45;
  assign t_r27_c46_9 = t_r27_c46_5 + t_r27_c46_6;
  assign t_r27_c46_10 = t_r27_c46_7 + t_r27_c46_8;
  assign t_r27_c46_11 = t_r27_c46_9 + t_r27_c46_10;
  assign t_r27_c46_12 = t_r27_c46_11 + p_28_47;
  assign out_27_46 = t_r27_c46_12 >> 4;

  assign t_r27_c47_0 = p_26_47 << 1;
  assign t_r27_c47_1 = p_27_46 << 1;
  assign t_r27_c47_2 = p_27_47 << 2;
  assign t_r27_c47_3 = p_27_48 << 1;
  assign t_r27_c47_4 = p_28_47 << 1;
  assign t_r27_c47_5 = t_r27_c47_0 + p_26_46;
  assign t_r27_c47_6 = t_r27_c47_1 + p_26_48;
  assign t_r27_c47_7 = t_r27_c47_2 + t_r27_c47_3;
  assign t_r27_c47_8 = t_r27_c47_4 + p_28_46;
  assign t_r27_c47_9 = t_r27_c47_5 + t_r27_c47_6;
  assign t_r27_c47_10 = t_r27_c47_7 + t_r27_c47_8;
  assign t_r27_c47_11 = t_r27_c47_9 + t_r27_c47_10;
  assign t_r27_c47_12 = t_r27_c47_11 + p_28_48;
  assign out_27_47 = t_r27_c47_12 >> 4;

  assign t_r27_c48_0 = p_26_48 << 1;
  assign t_r27_c48_1 = p_27_47 << 1;
  assign t_r27_c48_2 = p_27_48 << 2;
  assign t_r27_c48_3 = p_27_49 << 1;
  assign t_r27_c48_4 = p_28_48 << 1;
  assign t_r27_c48_5 = t_r27_c48_0 + p_26_47;
  assign t_r27_c48_6 = t_r27_c48_1 + p_26_49;
  assign t_r27_c48_7 = t_r27_c48_2 + t_r27_c48_3;
  assign t_r27_c48_8 = t_r27_c48_4 + p_28_47;
  assign t_r27_c48_9 = t_r27_c48_5 + t_r27_c48_6;
  assign t_r27_c48_10 = t_r27_c48_7 + t_r27_c48_8;
  assign t_r27_c48_11 = t_r27_c48_9 + t_r27_c48_10;
  assign t_r27_c48_12 = t_r27_c48_11 + p_28_49;
  assign out_27_48 = t_r27_c48_12 >> 4;

  assign t_r27_c49_0 = p_26_49 << 1;
  assign t_r27_c49_1 = p_27_48 << 1;
  assign t_r27_c49_2 = p_27_49 << 2;
  assign t_r27_c49_3 = p_27_50 << 1;
  assign t_r27_c49_4 = p_28_49 << 1;
  assign t_r27_c49_5 = t_r27_c49_0 + p_26_48;
  assign t_r27_c49_6 = t_r27_c49_1 + p_26_50;
  assign t_r27_c49_7 = t_r27_c49_2 + t_r27_c49_3;
  assign t_r27_c49_8 = t_r27_c49_4 + p_28_48;
  assign t_r27_c49_9 = t_r27_c49_5 + t_r27_c49_6;
  assign t_r27_c49_10 = t_r27_c49_7 + t_r27_c49_8;
  assign t_r27_c49_11 = t_r27_c49_9 + t_r27_c49_10;
  assign t_r27_c49_12 = t_r27_c49_11 + p_28_50;
  assign out_27_49 = t_r27_c49_12 >> 4;

  assign t_r27_c50_0 = p_26_50 << 1;
  assign t_r27_c50_1 = p_27_49 << 1;
  assign t_r27_c50_2 = p_27_50 << 2;
  assign t_r27_c50_3 = p_27_51 << 1;
  assign t_r27_c50_4 = p_28_50 << 1;
  assign t_r27_c50_5 = t_r27_c50_0 + p_26_49;
  assign t_r27_c50_6 = t_r27_c50_1 + p_26_51;
  assign t_r27_c50_7 = t_r27_c50_2 + t_r27_c50_3;
  assign t_r27_c50_8 = t_r27_c50_4 + p_28_49;
  assign t_r27_c50_9 = t_r27_c50_5 + t_r27_c50_6;
  assign t_r27_c50_10 = t_r27_c50_7 + t_r27_c50_8;
  assign t_r27_c50_11 = t_r27_c50_9 + t_r27_c50_10;
  assign t_r27_c50_12 = t_r27_c50_11 + p_28_51;
  assign out_27_50 = t_r27_c50_12 >> 4;

  assign t_r27_c51_0 = p_26_51 << 1;
  assign t_r27_c51_1 = p_27_50 << 1;
  assign t_r27_c51_2 = p_27_51 << 2;
  assign t_r27_c51_3 = p_27_52 << 1;
  assign t_r27_c51_4 = p_28_51 << 1;
  assign t_r27_c51_5 = t_r27_c51_0 + p_26_50;
  assign t_r27_c51_6 = t_r27_c51_1 + p_26_52;
  assign t_r27_c51_7 = t_r27_c51_2 + t_r27_c51_3;
  assign t_r27_c51_8 = t_r27_c51_4 + p_28_50;
  assign t_r27_c51_9 = t_r27_c51_5 + t_r27_c51_6;
  assign t_r27_c51_10 = t_r27_c51_7 + t_r27_c51_8;
  assign t_r27_c51_11 = t_r27_c51_9 + t_r27_c51_10;
  assign t_r27_c51_12 = t_r27_c51_11 + p_28_52;
  assign out_27_51 = t_r27_c51_12 >> 4;

  assign t_r27_c52_0 = p_26_52 << 1;
  assign t_r27_c52_1 = p_27_51 << 1;
  assign t_r27_c52_2 = p_27_52 << 2;
  assign t_r27_c52_3 = p_27_53 << 1;
  assign t_r27_c52_4 = p_28_52 << 1;
  assign t_r27_c52_5 = t_r27_c52_0 + p_26_51;
  assign t_r27_c52_6 = t_r27_c52_1 + p_26_53;
  assign t_r27_c52_7 = t_r27_c52_2 + t_r27_c52_3;
  assign t_r27_c52_8 = t_r27_c52_4 + p_28_51;
  assign t_r27_c52_9 = t_r27_c52_5 + t_r27_c52_6;
  assign t_r27_c52_10 = t_r27_c52_7 + t_r27_c52_8;
  assign t_r27_c52_11 = t_r27_c52_9 + t_r27_c52_10;
  assign t_r27_c52_12 = t_r27_c52_11 + p_28_53;
  assign out_27_52 = t_r27_c52_12 >> 4;

  assign t_r27_c53_0 = p_26_53 << 1;
  assign t_r27_c53_1 = p_27_52 << 1;
  assign t_r27_c53_2 = p_27_53 << 2;
  assign t_r27_c53_3 = p_27_54 << 1;
  assign t_r27_c53_4 = p_28_53 << 1;
  assign t_r27_c53_5 = t_r27_c53_0 + p_26_52;
  assign t_r27_c53_6 = t_r27_c53_1 + p_26_54;
  assign t_r27_c53_7 = t_r27_c53_2 + t_r27_c53_3;
  assign t_r27_c53_8 = t_r27_c53_4 + p_28_52;
  assign t_r27_c53_9 = t_r27_c53_5 + t_r27_c53_6;
  assign t_r27_c53_10 = t_r27_c53_7 + t_r27_c53_8;
  assign t_r27_c53_11 = t_r27_c53_9 + t_r27_c53_10;
  assign t_r27_c53_12 = t_r27_c53_11 + p_28_54;
  assign out_27_53 = t_r27_c53_12 >> 4;

  assign t_r27_c54_0 = p_26_54 << 1;
  assign t_r27_c54_1 = p_27_53 << 1;
  assign t_r27_c54_2 = p_27_54 << 2;
  assign t_r27_c54_3 = p_27_55 << 1;
  assign t_r27_c54_4 = p_28_54 << 1;
  assign t_r27_c54_5 = t_r27_c54_0 + p_26_53;
  assign t_r27_c54_6 = t_r27_c54_1 + p_26_55;
  assign t_r27_c54_7 = t_r27_c54_2 + t_r27_c54_3;
  assign t_r27_c54_8 = t_r27_c54_4 + p_28_53;
  assign t_r27_c54_9 = t_r27_c54_5 + t_r27_c54_6;
  assign t_r27_c54_10 = t_r27_c54_7 + t_r27_c54_8;
  assign t_r27_c54_11 = t_r27_c54_9 + t_r27_c54_10;
  assign t_r27_c54_12 = t_r27_c54_11 + p_28_55;
  assign out_27_54 = t_r27_c54_12 >> 4;

  assign t_r27_c55_0 = p_26_55 << 1;
  assign t_r27_c55_1 = p_27_54 << 1;
  assign t_r27_c55_2 = p_27_55 << 2;
  assign t_r27_c55_3 = p_27_56 << 1;
  assign t_r27_c55_4 = p_28_55 << 1;
  assign t_r27_c55_5 = t_r27_c55_0 + p_26_54;
  assign t_r27_c55_6 = t_r27_c55_1 + p_26_56;
  assign t_r27_c55_7 = t_r27_c55_2 + t_r27_c55_3;
  assign t_r27_c55_8 = t_r27_c55_4 + p_28_54;
  assign t_r27_c55_9 = t_r27_c55_5 + t_r27_c55_6;
  assign t_r27_c55_10 = t_r27_c55_7 + t_r27_c55_8;
  assign t_r27_c55_11 = t_r27_c55_9 + t_r27_c55_10;
  assign t_r27_c55_12 = t_r27_c55_11 + p_28_56;
  assign out_27_55 = t_r27_c55_12 >> 4;

  assign t_r27_c56_0 = p_26_56 << 1;
  assign t_r27_c56_1 = p_27_55 << 1;
  assign t_r27_c56_2 = p_27_56 << 2;
  assign t_r27_c56_3 = p_27_57 << 1;
  assign t_r27_c56_4 = p_28_56 << 1;
  assign t_r27_c56_5 = t_r27_c56_0 + p_26_55;
  assign t_r27_c56_6 = t_r27_c56_1 + p_26_57;
  assign t_r27_c56_7 = t_r27_c56_2 + t_r27_c56_3;
  assign t_r27_c56_8 = t_r27_c56_4 + p_28_55;
  assign t_r27_c56_9 = t_r27_c56_5 + t_r27_c56_6;
  assign t_r27_c56_10 = t_r27_c56_7 + t_r27_c56_8;
  assign t_r27_c56_11 = t_r27_c56_9 + t_r27_c56_10;
  assign t_r27_c56_12 = t_r27_c56_11 + p_28_57;
  assign out_27_56 = t_r27_c56_12 >> 4;

  assign t_r27_c57_0 = p_26_57 << 1;
  assign t_r27_c57_1 = p_27_56 << 1;
  assign t_r27_c57_2 = p_27_57 << 2;
  assign t_r27_c57_3 = p_27_58 << 1;
  assign t_r27_c57_4 = p_28_57 << 1;
  assign t_r27_c57_5 = t_r27_c57_0 + p_26_56;
  assign t_r27_c57_6 = t_r27_c57_1 + p_26_58;
  assign t_r27_c57_7 = t_r27_c57_2 + t_r27_c57_3;
  assign t_r27_c57_8 = t_r27_c57_4 + p_28_56;
  assign t_r27_c57_9 = t_r27_c57_5 + t_r27_c57_6;
  assign t_r27_c57_10 = t_r27_c57_7 + t_r27_c57_8;
  assign t_r27_c57_11 = t_r27_c57_9 + t_r27_c57_10;
  assign t_r27_c57_12 = t_r27_c57_11 + p_28_58;
  assign out_27_57 = t_r27_c57_12 >> 4;

  assign t_r27_c58_0 = p_26_58 << 1;
  assign t_r27_c58_1 = p_27_57 << 1;
  assign t_r27_c58_2 = p_27_58 << 2;
  assign t_r27_c58_3 = p_27_59 << 1;
  assign t_r27_c58_4 = p_28_58 << 1;
  assign t_r27_c58_5 = t_r27_c58_0 + p_26_57;
  assign t_r27_c58_6 = t_r27_c58_1 + p_26_59;
  assign t_r27_c58_7 = t_r27_c58_2 + t_r27_c58_3;
  assign t_r27_c58_8 = t_r27_c58_4 + p_28_57;
  assign t_r27_c58_9 = t_r27_c58_5 + t_r27_c58_6;
  assign t_r27_c58_10 = t_r27_c58_7 + t_r27_c58_8;
  assign t_r27_c58_11 = t_r27_c58_9 + t_r27_c58_10;
  assign t_r27_c58_12 = t_r27_c58_11 + p_28_59;
  assign out_27_58 = t_r27_c58_12 >> 4;

  assign t_r27_c59_0 = p_26_59 << 1;
  assign t_r27_c59_1 = p_27_58 << 1;
  assign t_r27_c59_2 = p_27_59 << 2;
  assign t_r27_c59_3 = p_27_60 << 1;
  assign t_r27_c59_4 = p_28_59 << 1;
  assign t_r27_c59_5 = t_r27_c59_0 + p_26_58;
  assign t_r27_c59_6 = t_r27_c59_1 + p_26_60;
  assign t_r27_c59_7 = t_r27_c59_2 + t_r27_c59_3;
  assign t_r27_c59_8 = t_r27_c59_4 + p_28_58;
  assign t_r27_c59_9 = t_r27_c59_5 + t_r27_c59_6;
  assign t_r27_c59_10 = t_r27_c59_7 + t_r27_c59_8;
  assign t_r27_c59_11 = t_r27_c59_9 + t_r27_c59_10;
  assign t_r27_c59_12 = t_r27_c59_11 + p_28_60;
  assign out_27_59 = t_r27_c59_12 >> 4;

  assign t_r27_c60_0 = p_26_60 << 1;
  assign t_r27_c60_1 = p_27_59 << 1;
  assign t_r27_c60_2 = p_27_60 << 2;
  assign t_r27_c60_3 = p_27_61 << 1;
  assign t_r27_c60_4 = p_28_60 << 1;
  assign t_r27_c60_5 = t_r27_c60_0 + p_26_59;
  assign t_r27_c60_6 = t_r27_c60_1 + p_26_61;
  assign t_r27_c60_7 = t_r27_c60_2 + t_r27_c60_3;
  assign t_r27_c60_8 = t_r27_c60_4 + p_28_59;
  assign t_r27_c60_9 = t_r27_c60_5 + t_r27_c60_6;
  assign t_r27_c60_10 = t_r27_c60_7 + t_r27_c60_8;
  assign t_r27_c60_11 = t_r27_c60_9 + t_r27_c60_10;
  assign t_r27_c60_12 = t_r27_c60_11 + p_28_61;
  assign out_27_60 = t_r27_c60_12 >> 4;

  assign t_r27_c61_0 = p_26_61 << 1;
  assign t_r27_c61_1 = p_27_60 << 1;
  assign t_r27_c61_2 = p_27_61 << 2;
  assign t_r27_c61_3 = p_27_62 << 1;
  assign t_r27_c61_4 = p_28_61 << 1;
  assign t_r27_c61_5 = t_r27_c61_0 + p_26_60;
  assign t_r27_c61_6 = t_r27_c61_1 + p_26_62;
  assign t_r27_c61_7 = t_r27_c61_2 + t_r27_c61_3;
  assign t_r27_c61_8 = t_r27_c61_4 + p_28_60;
  assign t_r27_c61_9 = t_r27_c61_5 + t_r27_c61_6;
  assign t_r27_c61_10 = t_r27_c61_7 + t_r27_c61_8;
  assign t_r27_c61_11 = t_r27_c61_9 + t_r27_c61_10;
  assign t_r27_c61_12 = t_r27_c61_11 + p_28_62;
  assign out_27_61 = t_r27_c61_12 >> 4;

  assign t_r27_c62_0 = p_26_62 << 1;
  assign t_r27_c62_1 = p_27_61 << 1;
  assign t_r27_c62_2 = p_27_62 << 2;
  assign t_r27_c62_3 = p_27_63 << 1;
  assign t_r27_c62_4 = p_28_62 << 1;
  assign t_r27_c62_5 = t_r27_c62_0 + p_26_61;
  assign t_r27_c62_6 = t_r27_c62_1 + p_26_63;
  assign t_r27_c62_7 = t_r27_c62_2 + t_r27_c62_3;
  assign t_r27_c62_8 = t_r27_c62_4 + p_28_61;
  assign t_r27_c62_9 = t_r27_c62_5 + t_r27_c62_6;
  assign t_r27_c62_10 = t_r27_c62_7 + t_r27_c62_8;
  assign t_r27_c62_11 = t_r27_c62_9 + t_r27_c62_10;
  assign t_r27_c62_12 = t_r27_c62_11 + p_28_63;
  assign out_27_62 = t_r27_c62_12 >> 4;

  assign t_r27_c63_0 = p_26_63 << 1;
  assign t_r27_c63_1 = p_27_62 << 1;
  assign t_r27_c63_2 = p_27_63 << 2;
  assign t_r27_c63_3 = p_27_64 << 1;
  assign t_r27_c63_4 = p_28_63 << 1;
  assign t_r27_c63_5 = t_r27_c63_0 + p_26_62;
  assign t_r27_c63_6 = t_r27_c63_1 + p_26_64;
  assign t_r27_c63_7 = t_r27_c63_2 + t_r27_c63_3;
  assign t_r27_c63_8 = t_r27_c63_4 + p_28_62;
  assign t_r27_c63_9 = t_r27_c63_5 + t_r27_c63_6;
  assign t_r27_c63_10 = t_r27_c63_7 + t_r27_c63_8;
  assign t_r27_c63_11 = t_r27_c63_9 + t_r27_c63_10;
  assign t_r27_c63_12 = t_r27_c63_11 + p_28_64;
  assign out_27_63 = t_r27_c63_12 >> 4;

  assign t_r27_c64_0 = p_26_64 << 1;
  assign t_r27_c64_1 = p_27_63 << 1;
  assign t_r27_c64_2 = p_27_64 << 2;
  assign t_r27_c64_3 = p_27_65 << 1;
  assign t_r27_c64_4 = p_28_64 << 1;
  assign t_r27_c64_5 = t_r27_c64_0 + p_26_63;
  assign t_r27_c64_6 = t_r27_c64_1 + p_26_65;
  assign t_r27_c64_7 = t_r27_c64_2 + t_r27_c64_3;
  assign t_r27_c64_8 = t_r27_c64_4 + p_28_63;
  assign t_r27_c64_9 = t_r27_c64_5 + t_r27_c64_6;
  assign t_r27_c64_10 = t_r27_c64_7 + t_r27_c64_8;
  assign t_r27_c64_11 = t_r27_c64_9 + t_r27_c64_10;
  assign t_r27_c64_12 = t_r27_c64_11 + p_28_65;
  assign out_27_64 = t_r27_c64_12 >> 4;

  assign t_r28_c1_0 = p_27_1 << 1;
  assign t_r28_c1_1 = p_28_0 << 1;
  assign t_r28_c1_2 = p_28_1 << 2;
  assign t_r28_c1_3 = p_28_2 << 1;
  assign t_r28_c1_4 = p_29_1 << 1;
  assign t_r28_c1_5 = t_r28_c1_0 + p_27_0;
  assign t_r28_c1_6 = t_r28_c1_1 + p_27_2;
  assign t_r28_c1_7 = t_r28_c1_2 + t_r28_c1_3;
  assign t_r28_c1_8 = t_r28_c1_4 + p_29_0;
  assign t_r28_c1_9 = t_r28_c1_5 + t_r28_c1_6;
  assign t_r28_c1_10 = t_r28_c1_7 + t_r28_c1_8;
  assign t_r28_c1_11 = t_r28_c1_9 + t_r28_c1_10;
  assign t_r28_c1_12 = t_r28_c1_11 + p_29_2;
  assign out_28_1 = t_r28_c1_12 >> 4;

  assign t_r28_c2_0 = p_27_2 << 1;
  assign t_r28_c2_1 = p_28_1 << 1;
  assign t_r28_c2_2 = p_28_2 << 2;
  assign t_r28_c2_3 = p_28_3 << 1;
  assign t_r28_c2_4 = p_29_2 << 1;
  assign t_r28_c2_5 = t_r28_c2_0 + p_27_1;
  assign t_r28_c2_6 = t_r28_c2_1 + p_27_3;
  assign t_r28_c2_7 = t_r28_c2_2 + t_r28_c2_3;
  assign t_r28_c2_8 = t_r28_c2_4 + p_29_1;
  assign t_r28_c2_9 = t_r28_c2_5 + t_r28_c2_6;
  assign t_r28_c2_10 = t_r28_c2_7 + t_r28_c2_8;
  assign t_r28_c2_11 = t_r28_c2_9 + t_r28_c2_10;
  assign t_r28_c2_12 = t_r28_c2_11 + p_29_3;
  assign out_28_2 = t_r28_c2_12 >> 4;

  assign t_r28_c3_0 = p_27_3 << 1;
  assign t_r28_c3_1 = p_28_2 << 1;
  assign t_r28_c3_2 = p_28_3 << 2;
  assign t_r28_c3_3 = p_28_4 << 1;
  assign t_r28_c3_4 = p_29_3 << 1;
  assign t_r28_c3_5 = t_r28_c3_0 + p_27_2;
  assign t_r28_c3_6 = t_r28_c3_1 + p_27_4;
  assign t_r28_c3_7 = t_r28_c3_2 + t_r28_c3_3;
  assign t_r28_c3_8 = t_r28_c3_4 + p_29_2;
  assign t_r28_c3_9 = t_r28_c3_5 + t_r28_c3_6;
  assign t_r28_c3_10 = t_r28_c3_7 + t_r28_c3_8;
  assign t_r28_c3_11 = t_r28_c3_9 + t_r28_c3_10;
  assign t_r28_c3_12 = t_r28_c3_11 + p_29_4;
  assign out_28_3 = t_r28_c3_12 >> 4;

  assign t_r28_c4_0 = p_27_4 << 1;
  assign t_r28_c4_1 = p_28_3 << 1;
  assign t_r28_c4_2 = p_28_4 << 2;
  assign t_r28_c4_3 = p_28_5 << 1;
  assign t_r28_c4_4 = p_29_4 << 1;
  assign t_r28_c4_5 = t_r28_c4_0 + p_27_3;
  assign t_r28_c4_6 = t_r28_c4_1 + p_27_5;
  assign t_r28_c4_7 = t_r28_c4_2 + t_r28_c4_3;
  assign t_r28_c4_8 = t_r28_c4_4 + p_29_3;
  assign t_r28_c4_9 = t_r28_c4_5 + t_r28_c4_6;
  assign t_r28_c4_10 = t_r28_c4_7 + t_r28_c4_8;
  assign t_r28_c4_11 = t_r28_c4_9 + t_r28_c4_10;
  assign t_r28_c4_12 = t_r28_c4_11 + p_29_5;
  assign out_28_4 = t_r28_c4_12 >> 4;

  assign t_r28_c5_0 = p_27_5 << 1;
  assign t_r28_c5_1 = p_28_4 << 1;
  assign t_r28_c5_2 = p_28_5 << 2;
  assign t_r28_c5_3 = p_28_6 << 1;
  assign t_r28_c5_4 = p_29_5 << 1;
  assign t_r28_c5_5 = t_r28_c5_0 + p_27_4;
  assign t_r28_c5_6 = t_r28_c5_1 + p_27_6;
  assign t_r28_c5_7 = t_r28_c5_2 + t_r28_c5_3;
  assign t_r28_c5_8 = t_r28_c5_4 + p_29_4;
  assign t_r28_c5_9 = t_r28_c5_5 + t_r28_c5_6;
  assign t_r28_c5_10 = t_r28_c5_7 + t_r28_c5_8;
  assign t_r28_c5_11 = t_r28_c5_9 + t_r28_c5_10;
  assign t_r28_c5_12 = t_r28_c5_11 + p_29_6;
  assign out_28_5 = t_r28_c5_12 >> 4;

  assign t_r28_c6_0 = p_27_6 << 1;
  assign t_r28_c6_1 = p_28_5 << 1;
  assign t_r28_c6_2 = p_28_6 << 2;
  assign t_r28_c6_3 = p_28_7 << 1;
  assign t_r28_c6_4 = p_29_6 << 1;
  assign t_r28_c6_5 = t_r28_c6_0 + p_27_5;
  assign t_r28_c6_6 = t_r28_c6_1 + p_27_7;
  assign t_r28_c6_7 = t_r28_c6_2 + t_r28_c6_3;
  assign t_r28_c6_8 = t_r28_c6_4 + p_29_5;
  assign t_r28_c6_9 = t_r28_c6_5 + t_r28_c6_6;
  assign t_r28_c6_10 = t_r28_c6_7 + t_r28_c6_8;
  assign t_r28_c6_11 = t_r28_c6_9 + t_r28_c6_10;
  assign t_r28_c6_12 = t_r28_c6_11 + p_29_7;
  assign out_28_6 = t_r28_c6_12 >> 4;

  assign t_r28_c7_0 = p_27_7 << 1;
  assign t_r28_c7_1 = p_28_6 << 1;
  assign t_r28_c7_2 = p_28_7 << 2;
  assign t_r28_c7_3 = p_28_8 << 1;
  assign t_r28_c7_4 = p_29_7 << 1;
  assign t_r28_c7_5 = t_r28_c7_0 + p_27_6;
  assign t_r28_c7_6 = t_r28_c7_1 + p_27_8;
  assign t_r28_c7_7 = t_r28_c7_2 + t_r28_c7_3;
  assign t_r28_c7_8 = t_r28_c7_4 + p_29_6;
  assign t_r28_c7_9 = t_r28_c7_5 + t_r28_c7_6;
  assign t_r28_c7_10 = t_r28_c7_7 + t_r28_c7_8;
  assign t_r28_c7_11 = t_r28_c7_9 + t_r28_c7_10;
  assign t_r28_c7_12 = t_r28_c7_11 + p_29_8;
  assign out_28_7 = t_r28_c7_12 >> 4;

  assign t_r28_c8_0 = p_27_8 << 1;
  assign t_r28_c8_1 = p_28_7 << 1;
  assign t_r28_c8_2 = p_28_8 << 2;
  assign t_r28_c8_3 = p_28_9 << 1;
  assign t_r28_c8_4 = p_29_8 << 1;
  assign t_r28_c8_5 = t_r28_c8_0 + p_27_7;
  assign t_r28_c8_6 = t_r28_c8_1 + p_27_9;
  assign t_r28_c8_7 = t_r28_c8_2 + t_r28_c8_3;
  assign t_r28_c8_8 = t_r28_c8_4 + p_29_7;
  assign t_r28_c8_9 = t_r28_c8_5 + t_r28_c8_6;
  assign t_r28_c8_10 = t_r28_c8_7 + t_r28_c8_8;
  assign t_r28_c8_11 = t_r28_c8_9 + t_r28_c8_10;
  assign t_r28_c8_12 = t_r28_c8_11 + p_29_9;
  assign out_28_8 = t_r28_c8_12 >> 4;

  assign t_r28_c9_0 = p_27_9 << 1;
  assign t_r28_c9_1 = p_28_8 << 1;
  assign t_r28_c9_2 = p_28_9 << 2;
  assign t_r28_c9_3 = p_28_10 << 1;
  assign t_r28_c9_4 = p_29_9 << 1;
  assign t_r28_c9_5 = t_r28_c9_0 + p_27_8;
  assign t_r28_c9_6 = t_r28_c9_1 + p_27_10;
  assign t_r28_c9_7 = t_r28_c9_2 + t_r28_c9_3;
  assign t_r28_c9_8 = t_r28_c9_4 + p_29_8;
  assign t_r28_c9_9 = t_r28_c9_5 + t_r28_c9_6;
  assign t_r28_c9_10 = t_r28_c9_7 + t_r28_c9_8;
  assign t_r28_c9_11 = t_r28_c9_9 + t_r28_c9_10;
  assign t_r28_c9_12 = t_r28_c9_11 + p_29_10;
  assign out_28_9 = t_r28_c9_12 >> 4;

  assign t_r28_c10_0 = p_27_10 << 1;
  assign t_r28_c10_1 = p_28_9 << 1;
  assign t_r28_c10_2 = p_28_10 << 2;
  assign t_r28_c10_3 = p_28_11 << 1;
  assign t_r28_c10_4 = p_29_10 << 1;
  assign t_r28_c10_5 = t_r28_c10_0 + p_27_9;
  assign t_r28_c10_6 = t_r28_c10_1 + p_27_11;
  assign t_r28_c10_7 = t_r28_c10_2 + t_r28_c10_3;
  assign t_r28_c10_8 = t_r28_c10_4 + p_29_9;
  assign t_r28_c10_9 = t_r28_c10_5 + t_r28_c10_6;
  assign t_r28_c10_10 = t_r28_c10_7 + t_r28_c10_8;
  assign t_r28_c10_11 = t_r28_c10_9 + t_r28_c10_10;
  assign t_r28_c10_12 = t_r28_c10_11 + p_29_11;
  assign out_28_10 = t_r28_c10_12 >> 4;

  assign t_r28_c11_0 = p_27_11 << 1;
  assign t_r28_c11_1 = p_28_10 << 1;
  assign t_r28_c11_2 = p_28_11 << 2;
  assign t_r28_c11_3 = p_28_12 << 1;
  assign t_r28_c11_4 = p_29_11 << 1;
  assign t_r28_c11_5 = t_r28_c11_0 + p_27_10;
  assign t_r28_c11_6 = t_r28_c11_1 + p_27_12;
  assign t_r28_c11_7 = t_r28_c11_2 + t_r28_c11_3;
  assign t_r28_c11_8 = t_r28_c11_4 + p_29_10;
  assign t_r28_c11_9 = t_r28_c11_5 + t_r28_c11_6;
  assign t_r28_c11_10 = t_r28_c11_7 + t_r28_c11_8;
  assign t_r28_c11_11 = t_r28_c11_9 + t_r28_c11_10;
  assign t_r28_c11_12 = t_r28_c11_11 + p_29_12;
  assign out_28_11 = t_r28_c11_12 >> 4;

  assign t_r28_c12_0 = p_27_12 << 1;
  assign t_r28_c12_1 = p_28_11 << 1;
  assign t_r28_c12_2 = p_28_12 << 2;
  assign t_r28_c12_3 = p_28_13 << 1;
  assign t_r28_c12_4 = p_29_12 << 1;
  assign t_r28_c12_5 = t_r28_c12_0 + p_27_11;
  assign t_r28_c12_6 = t_r28_c12_1 + p_27_13;
  assign t_r28_c12_7 = t_r28_c12_2 + t_r28_c12_3;
  assign t_r28_c12_8 = t_r28_c12_4 + p_29_11;
  assign t_r28_c12_9 = t_r28_c12_5 + t_r28_c12_6;
  assign t_r28_c12_10 = t_r28_c12_7 + t_r28_c12_8;
  assign t_r28_c12_11 = t_r28_c12_9 + t_r28_c12_10;
  assign t_r28_c12_12 = t_r28_c12_11 + p_29_13;
  assign out_28_12 = t_r28_c12_12 >> 4;

  assign t_r28_c13_0 = p_27_13 << 1;
  assign t_r28_c13_1 = p_28_12 << 1;
  assign t_r28_c13_2 = p_28_13 << 2;
  assign t_r28_c13_3 = p_28_14 << 1;
  assign t_r28_c13_4 = p_29_13 << 1;
  assign t_r28_c13_5 = t_r28_c13_0 + p_27_12;
  assign t_r28_c13_6 = t_r28_c13_1 + p_27_14;
  assign t_r28_c13_7 = t_r28_c13_2 + t_r28_c13_3;
  assign t_r28_c13_8 = t_r28_c13_4 + p_29_12;
  assign t_r28_c13_9 = t_r28_c13_5 + t_r28_c13_6;
  assign t_r28_c13_10 = t_r28_c13_7 + t_r28_c13_8;
  assign t_r28_c13_11 = t_r28_c13_9 + t_r28_c13_10;
  assign t_r28_c13_12 = t_r28_c13_11 + p_29_14;
  assign out_28_13 = t_r28_c13_12 >> 4;

  assign t_r28_c14_0 = p_27_14 << 1;
  assign t_r28_c14_1 = p_28_13 << 1;
  assign t_r28_c14_2 = p_28_14 << 2;
  assign t_r28_c14_3 = p_28_15 << 1;
  assign t_r28_c14_4 = p_29_14 << 1;
  assign t_r28_c14_5 = t_r28_c14_0 + p_27_13;
  assign t_r28_c14_6 = t_r28_c14_1 + p_27_15;
  assign t_r28_c14_7 = t_r28_c14_2 + t_r28_c14_3;
  assign t_r28_c14_8 = t_r28_c14_4 + p_29_13;
  assign t_r28_c14_9 = t_r28_c14_5 + t_r28_c14_6;
  assign t_r28_c14_10 = t_r28_c14_7 + t_r28_c14_8;
  assign t_r28_c14_11 = t_r28_c14_9 + t_r28_c14_10;
  assign t_r28_c14_12 = t_r28_c14_11 + p_29_15;
  assign out_28_14 = t_r28_c14_12 >> 4;

  assign t_r28_c15_0 = p_27_15 << 1;
  assign t_r28_c15_1 = p_28_14 << 1;
  assign t_r28_c15_2 = p_28_15 << 2;
  assign t_r28_c15_3 = p_28_16 << 1;
  assign t_r28_c15_4 = p_29_15 << 1;
  assign t_r28_c15_5 = t_r28_c15_0 + p_27_14;
  assign t_r28_c15_6 = t_r28_c15_1 + p_27_16;
  assign t_r28_c15_7 = t_r28_c15_2 + t_r28_c15_3;
  assign t_r28_c15_8 = t_r28_c15_4 + p_29_14;
  assign t_r28_c15_9 = t_r28_c15_5 + t_r28_c15_6;
  assign t_r28_c15_10 = t_r28_c15_7 + t_r28_c15_8;
  assign t_r28_c15_11 = t_r28_c15_9 + t_r28_c15_10;
  assign t_r28_c15_12 = t_r28_c15_11 + p_29_16;
  assign out_28_15 = t_r28_c15_12 >> 4;

  assign t_r28_c16_0 = p_27_16 << 1;
  assign t_r28_c16_1 = p_28_15 << 1;
  assign t_r28_c16_2 = p_28_16 << 2;
  assign t_r28_c16_3 = p_28_17 << 1;
  assign t_r28_c16_4 = p_29_16 << 1;
  assign t_r28_c16_5 = t_r28_c16_0 + p_27_15;
  assign t_r28_c16_6 = t_r28_c16_1 + p_27_17;
  assign t_r28_c16_7 = t_r28_c16_2 + t_r28_c16_3;
  assign t_r28_c16_8 = t_r28_c16_4 + p_29_15;
  assign t_r28_c16_9 = t_r28_c16_5 + t_r28_c16_6;
  assign t_r28_c16_10 = t_r28_c16_7 + t_r28_c16_8;
  assign t_r28_c16_11 = t_r28_c16_9 + t_r28_c16_10;
  assign t_r28_c16_12 = t_r28_c16_11 + p_29_17;
  assign out_28_16 = t_r28_c16_12 >> 4;

  assign t_r28_c17_0 = p_27_17 << 1;
  assign t_r28_c17_1 = p_28_16 << 1;
  assign t_r28_c17_2 = p_28_17 << 2;
  assign t_r28_c17_3 = p_28_18 << 1;
  assign t_r28_c17_4 = p_29_17 << 1;
  assign t_r28_c17_5 = t_r28_c17_0 + p_27_16;
  assign t_r28_c17_6 = t_r28_c17_1 + p_27_18;
  assign t_r28_c17_7 = t_r28_c17_2 + t_r28_c17_3;
  assign t_r28_c17_8 = t_r28_c17_4 + p_29_16;
  assign t_r28_c17_9 = t_r28_c17_5 + t_r28_c17_6;
  assign t_r28_c17_10 = t_r28_c17_7 + t_r28_c17_8;
  assign t_r28_c17_11 = t_r28_c17_9 + t_r28_c17_10;
  assign t_r28_c17_12 = t_r28_c17_11 + p_29_18;
  assign out_28_17 = t_r28_c17_12 >> 4;

  assign t_r28_c18_0 = p_27_18 << 1;
  assign t_r28_c18_1 = p_28_17 << 1;
  assign t_r28_c18_2 = p_28_18 << 2;
  assign t_r28_c18_3 = p_28_19 << 1;
  assign t_r28_c18_4 = p_29_18 << 1;
  assign t_r28_c18_5 = t_r28_c18_0 + p_27_17;
  assign t_r28_c18_6 = t_r28_c18_1 + p_27_19;
  assign t_r28_c18_7 = t_r28_c18_2 + t_r28_c18_3;
  assign t_r28_c18_8 = t_r28_c18_4 + p_29_17;
  assign t_r28_c18_9 = t_r28_c18_5 + t_r28_c18_6;
  assign t_r28_c18_10 = t_r28_c18_7 + t_r28_c18_8;
  assign t_r28_c18_11 = t_r28_c18_9 + t_r28_c18_10;
  assign t_r28_c18_12 = t_r28_c18_11 + p_29_19;
  assign out_28_18 = t_r28_c18_12 >> 4;

  assign t_r28_c19_0 = p_27_19 << 1;
  assign t_r28_c19_1 = p_28_18 << 1;
  assign t_r28_c19_2 = p_28_19 << 2;
  assign t_r28_c19_3 = p_28_20 << 1;
  assign t_r28_c19_4 = p_29_19 << 1;
  assign t_r28_c19_5 = t_r28_c19_0 + p_27_18;
  assign t_r28_c19_6 = t_r28_c19_1 + p_27_20;
  assign t_r28_c19_7 = t_r28_c19_2 + t_r28_c19_3;
  assign t_r28_c19_8 = t_r28_c19_4 + p_29_18;
  assign t_r28_c19_9 = t_r28_c19_5 + t_r28_c19_6;
  assign t_r28_c19_10 = t_r28_c19_7 + t_r28_c19_8;
  assign t_r28_c19_11 = t_r28_c19_9 + t_r28_c19_10;
  assign t_r28_c19_12 = t_r28_c19_11 + p_29_20;
  assign out_28_19 = t_r28_c19_12 >> 4;

  assign t_r28_c20_0 = p_27_20 << 1;
  assign t_r28_c20_1 = p_28_19 << 1;
  assign t_r28_c20_2 = p_28_20 << 2;
  assign t_r28_c20_3 = p_28_21 << 1;
  assign t_r28_c20_4 = p_29_20 << 1;
  assign t_r28_c20_5 = t_r28_c20_0 + p_27_19;
  assign t_r28_c20_6 = t_r28_c20_1 + p_27_21;
  assign t_r28_c20_7 = t_r28_c20_2 + t_r28_c20_3;
  assign t_r28_c20_8 = t_r28_c20_4 + p_29_19;
  assign t_r28_c20_9 = t_r28_c20_5 + t_r28_c20_6;
  assign t_r28_c20_10 = t_r28_c20_7 + t_r28_c20_8;
  assign t_r28_c20_11 = t_r28_c20_9 + t_r28_c20_10;
  assign t_r28_c20_12 = t_r28_c20_11 + p_29_21;
  assign out_28_20 = t_r28_c20_12 >> 4;

  assign t_r28_c21_0 = p_27_21 << 1;
  assign t_r28_c21_1 = p_28_20 << 1;
  assign t_r28_c21_2 = p_28_21 << 2;
  assign t_r28_c21_3 = p_28_22 << 1;
  assign t_r28_c21_4 = p_29_21 << 1;
  assign t_r28_c21_5 = t_r28_c21_0 + p_27_20;
  assign t_r28_c21_6 = t_r28_c21_1 + p_27_22;
  assign t_r28_c21_7 = t_r28_c21_2 + t_r28_c21_3;
  assign t_r28_c21_8 = t_r28_c21_4 + p_29_20;
  assign t_r28_c21_9 = t_r28_c21_5 + t_r28_c21_6;
  assign t_r28_c21_10 = t_r28_c21_7 + t_r28_c21_8;
  assign t_r28_c21_11 = t_r28_c21_9 + t_r28_c21_10;
  assign t_r28_c21_12 = t_r28_c21_11 + p_29_22;
  assign out_28_21 = t_r28_c21_12 >> 4;

  assign t_r28_c22_0 = p_27_22 << 1;
  assign t_r28_c22_1 = p_28_21 << 1;
  assign t_r28_c22_2 = p_28_22 << 2;
  assign t_r28_c22_3 = p_28_23 << 1;
  assign t_r28_c22_4 = p_29_22 << 1;
  assign t_r28_c22_5 = t_r28_c22_0 + p_27_21;
  assign t_r28_c22_6 = t_r28_c22_1 + p_27_23;
  assign t_r28_c22_7 = t_r28_c22_2 + t_r28_c22_3;
  assign t_r28_c22_8 = t_r28_c22_4 + p_29_21;
  assign t_r28_c22_9 = t_r28_c22_5 + t_r28_c22_6;
  assign t_r28_c22_10 = t_r28_c22_7 + t_r28_c22_8;
  assign t_r28_c22_11 = t_r28_c22_9 + t_r28_c22_10;
  assign t_r28_c22_12 = t_r28_c22_11 + p_29_23;
  assign out_28_22 = t_r28_c22_12 >> 4;

  assign t_r28_c23_0 = p_27_23 << 1;
  assign t_r28_c23_1 = p_28_22 << 1;
  assign t_r28_c23_2 = p_28_23 << 2;
  assign t_r28_c23_3 = p_28_24 << 1;
  assign t_r28_c23_4 = p_29_23 << 1;
  assign t_r28_c23_5 = t_r28_c23_0 + p_27_22;
  assign t_r28_c23_6 = t_r28_c23_1 + p_27_24;
  assign t_r28_c23_7 = t_r28_c23_2 + t_r28_c23_3;
  assign t_r28_c23_8 = t_r28_c23_4 + p_29_22;
  assign t_r28_c23_9 = t_r28_c23_5 + t_r28_c23_6;
  assign t_r28_c23_10 = t_r28_c23_7 + t_r28_c23_8;
  assign t_r28_c23_11 = t_r28_c23_9 + t_r28_c23_10;
  assign t_r28_c23_12 = t_r28_c23_11 + p_29_24;
  assign out_28_23 = t_r28_c23_12 >> 4;

  assign t_r28_c24_0 = p_27_24 << 1;
  assign t_r28_c24_1 = p_28_23 << 1;
  assign t_r28_c24_2 = p_28_24 << 2;
  assign t_r28_c24_3 = p_28_25 << 1;
  assign t_r28_c24_4 = p_29_24 << 1;
  assign t_r28_c24_5 = t_r28_c24_0 + p_27_23;
  assign t_r28_c24_6 = t_r28_c24_1 + p_27_25;
  assign t_r28_c24_7 = t_r28_c24_2 + t_r28_c24_3;
  assign t_r28_c24_8 = t_r28_c24_4 + p_29_23;
  assign t_r28_c24_9 = t_r28_c24_5 + t_r28_c24_6;
  assign t_r28_c24_10 = t_r28_c24_7 + t_r28_c24_8;
  assign t_r28_c24_11 = t_r28_c24_9 + t_r28_c24_10;
  assign t_r28_c24_12 = t_r28_c24_11 + p_29_25;
  assign out_28_24 = t_r28_c24_12 >> 4;

  assign t_r28_c25_0 = p_27_25 << 1;
  assign t_r28_c25_1 = p_28_24 << 1;
  assign t_r28_c25_2 = p_28_25 << 2;
  assign t_r28_c25_3 = p_28_26 << 1;
  assign t_r28_c25_4 = p_29_25 << 1;
  assign t_r28_c25_5 = t_r28_c25_0 + p_27_24;
  assign t_r28_c25_6 = t_r28_c25_1 + p_27_26;
  assign t_r28_c25_7 = t_r28_c25_2 + t_r28_c25_3;
  assign t_r28_c25_8 = t_r28_c25_4 + p_29_24;
  assign t_r28_c25_9 = t_r28_c25_5 + t_r28_c25_6;
  assign t_r28_c25_10 = t_r28_c25_7 + t_r28_c25_8;
  assign t_r28_c25_11 = t_r28_c25_9 + t_r28_c25_10;
  assign t_r28_c25_12 = t_r28_c25_11 + p_29_26;
  assign out_28_25 = t_r28_c25_12 >> 4;

  assign t_r28_c26_0 = p_27_26 << 1;
  assign t_r28_c26_1 = p_28_25 << 1;
  assign t_r28_c26_2 = p_28_26 << 2;
  assign t_r28_c26_3 = p_28_27 << 1;
  assign t_r28_c26_4 = p_29_26 << 1;
  assign t_r28_c26_5 = t_r28_c26_0 + p_27_25;
  assign t_r28_c26_6 = t_r28_c26_1 + p_27_27;
  assign t_r28_c26_7 = t_r28_c26_2 + t_r28_c26_3;
  assign t_r28_c26_8 = t_r28_c26_4 + p_29_25;
  assign t_r28_c26_9 = t_r28_c26_5 + t_r28_c26_6;
  assign t_r28_c26_10 = t_r28_c26_7 + t_r28_c26_8;
  assign t_r28_c26_11 = t_r28_c26_9 + t_r28_c26_10;
  assign t_r28_c26_12 = t_r28_c26_11 + p_29_27;
  assign out_28_26 = t_r28_c26_12 >> 4;

  assign t_r28_c27_0 = p_27_27 << 1;
  assign t_r28_c27_1 = p_28_26 << 1;
  assign t_r28_c27_2 = p_28_27 << 2;
  assign t_r28_c27_3 = p_28_28 << 1;
  assign t_r28_c27_4 = p_29_27 << 1;
  assign t_r28_c27_5 = t_r28_c27_0 + p_27_26;
  assign t_r28_c27_6 = t_r28_c27_1 + p_27_28;
  assign t_r28_c27_7 = t_r28_c27_2 + t_r28_c27_3;
  assign t_r28_c27_8 = t_r28_c27_4 + p_29_26;
  assign t_r28_c27_9 = t_r28_c27_5 + t_r28_c27_6;
  assign t_r28_c27_10 = t_r28_c27_7 + t_r28_c27_8;
  assign t_r28_c27_11 = t_r28_c27_9 + t_r28_c27_10;
  assign t_r28_c27_12 = t_r28_c27_11 + p_29_28;
  assign out_28_27 = t_r28_c27_12 >> 4;

  assign t_r28_c28_0 = p_27_28 << 1;
  assign t_r28_c28_1 = p_28_27 << 1;
  assign t_r28_c28_2 = p_28_28 << 2;
  assign t_r28_c28_3 = p_28_29 << 1;
  assign t_r28_c28_4 = p_29_28 << 1;
  assign t_r28_c28_5 = t_r28_c28_0 + p_27_27;
  assign t_r28_c28_6 = t_r28_c28_1 + p_27_29;
  assign t_r28_c28_7 = t_r28_c28_2 + t_r28_c28_3;
  assign t_r28_c28_8 = t_r28_c28_4 + p_29_27;
  assign t_r28_c28_9 = t_r28_c28_5 + t_r28_c28_6;
  assign t_r28_c28_10 = t_r28_c28_7 + t_r28_c28_8;
  assign t_r28_c28_11 = t_r28_c28_9 + t_r28_c28_10;
  assign t_r28_c28_12 = t_r28_c28_11 + p_29_29;
  assign out_28_28 = t_r28_c28_12 >> 4;

  assign t_r28_c29_0 = p_27_29 << 1;
  assign t_r28_c29_1 = p_28_28 << 1;
  assign t_r28_c29_2 = p_28_29 << 2;
  assign t_r28_c29_3 = p_28_30 << 1;
  assign t_r28_c29_4 = p_29_29 << 1;
  assign t_r28_c29_5 = t_r28_c29_0 + p_27_28;
  assign t_r28_c29_6 = t_r28_c29_1 + p_27_30;
  assign t_r28_c29_7 = t_r28_c29_2 + t_r28_c29_3;
  assign t_r28_c29_8 = t_r28_c29_4 + p_29_28;
  assign t_r28_c29_9 = t_r28_c29_5 + t_r28_c29_6;
  assign t_r28_c29_10 = t_r28_c29_7 + t_r28_c29_8;
  assign t_r28_c29_11 = t_r28_c29_9 + t_r28_c29_10;
  assign t_r28_c29_12 = t_r28_c29_11 + p_29_30;
  assign out_28_29 = t_r28_c29_12 >> 4;

  assign t_r28_c30_0 = p_27_30 << 1;
  assign t_r28_c30_1 = p_28_29 << 1;
  assign t_r28_c30_2 = p_28_30 << 2;
  assign t_r28_c30_3 = p_28_31 << 1;
  assign t_r28_c30_4 = p_29_30 << 1;
  assign t_r28_c30_5 = t_r28_c30_0 + p_27_29;
  assign t_r28_c30_6 = t_r28_c30_1 + p_27_31;
  assign t_r28_c30_7 = t_r28_c30_2 + t_r28_c30_3;
  assign t_r28_c30_8 = t_r28_c30_4 + p_29_29;
  assign t_r28_c30_9 = t_r28_c30_5 + t_r28_c30_6;
  assign t_r28_c30_10 = t_r28_c30_7 + t_r28_c30_8;
  assign t_r28_c30_11 = t_r28_c30_9 + t_r28_c30_10;
  assign t_r28_c30_12 = t_r28_c30_11 + p_29_31;
  assign out_28_30 = t_r28_c30_12 >> 4;

  assign t_r28_c31_0 = p_27_31 << 1;
  assign t_r28_c31_1 = p_28_30 << 1;
  assign t_r28_c31_2 = p_28_31 << 2;
  assign t_r28_c31_3 = p_28_32 << 1;
  assign t_r28_c31_4 = p_29_31 << 1;
  assign t_r28_c31_5 = t_r28_c31_0 + p_27_30;
  assign t_r28_c31_6 = t_r28_c31_1 + p_27_32;
  assign t_r28_c31_7 = t_r28_c31_2 + t_r28_c31_3;
  assign t_r28_c31_8 = t_r28_c31_4 + p_29_30;
  assign t_r28_c31_9 = t_r28_c31_5 + t_r28_c31_6;
  assign t_r28_c31_10 = t_r28_c31_7 + t_r28_c31_8;
  assign t_r28_c31_11 = t_r28_c31_9 + t_r28_c31_10;
  assign t_r28_c31_12 = t_r28_c31_11 + p_29_32;
  assign out_28_31 = t_r28_c31_12 >> 4;

  assign t_r28_c32_0 = p_27_32 << 1;
  assign t_r28_c32_1 = p_28_31 << 1;
  assign t_r28_c32_2 = p_28_32 << 2;
  assign t_r28_c32_3 = p_28_33 << 1;
  assign t_r28_c32_4 = p_29_32 << 1;
  assign t_r28_c32_5 = t_r28_c32_0 + p_27_31;
  assign t_r28_c32_6 = t_r28_c32_1 + p_27_33;
  assign t_r28_c32_7 = t_r28_c32_2 + t_r28_c32_3;
  assign t_r28_c32_8 = t_r28_c32_4 + p_29_31;
  assign t_r28_c32_9 = t_r28_c32_5 + t_r28_c32_6;
  assign t_r28_c32_10 = t_r28_c32_7 + t_r28_c32_8;
  assign t_r28_c32_11 = t_r28_c32_9 + t_r28_c32_10;
  assign t_r28_c32_12 = t_r28_c32_11 + p_29_33;
  assign out_28_32 = t_r28_c32_12 >> 4;

  assign t_r28_c33_0 = p_27_33 << 1;
  assign t_r28_c33_1 = p_28_32 << 1;
  assign t_r28_c33_2 = p_28_33 << 2;
  assign t_r28_c33_3 = p_28_34 << 1;
  assign t_r28_c33_4 = p_29_33 << 1;
  assign t_r28_c33_5 = t_r28_c33_0 + p_27_32;
  assign t_r28_c33_6 = t_r28_c33_1 + p_27_34;
  assign t_r28_c33_7 = t_r28_c33_2 + t_r28_c33_3;
  assign t_r28_c33_8 = t_r28_c33_4 + p_29_32;
  assign t_r28_c33_9 = t_r28_c33_5 + t_r28_c33_6;
  assign t_r28_c33_10 = t_r28_c33_7 + t_r28_c33_8;
  assign t_r28_c33_11 = t_r28_c33_9 + t_r28_c33_10;
  assign t_r28_c33_12 = t_r28_c33_11 + p_29_34;
  assign out_28_33 = t_r28_c33_12 >> 4;

  assign t_r28_c34_0 = p_27_34 << 1;
  assign t_r28_c34_1 = p_28_33 << 1;
  assign t_r28_c34_2 = p_28_34 << 2;
  assign t_r28_c34_3 = p_28_35 << 1;
  assign t_r28_c34_4 = p_29_34 << 1;
  assign t_r28_c34_5 = t_r28_c34_0 + p_27_33;
  assign t_r28_c34_6 = t_r28_c34_1 + p_27_35;
  assign t_r28_c34_7 = t_r28_c34_2 + t_r28_c34_3;
  assign t_r28_c34_8 = t_r28_c34_4 + p_29_33;
  assign t_r28_c34_9 = t_r28_c34_5 + t_r28_c34_6;
  assign t_r28_c34_10 = t_r28_c34_7 + t_r28_c34_8;
  assign t_r28_c34_11 = t_r28_c34_9 + t_r28_c34_10;
  assign t_r28_c34_12 = t_r28_c34_11 + p_29_35;
  assign out_28_34 = t_r28_c34_12 >> 4;

  assign t_r28_c35_0 = p_27_35 << 1;
  assign t_r28_c35_1 = p_28_34 << 1;
  assign t_r28_c35_2 = p_28_35 << 2;
  assign t_r28_c35_3 = p_28_36 << 1;
  assign t_r28_c35_4 = p_29_35 << 1;
  assign t_r28_c35_5 = t_r28_c35_0 + p_27_34;
  assign t_r28_c35_6 = t_r28_c35_1 + p_27_36;
  assign t_r28_c35_7 = t_r28_c35_2 + t_r28_c35_3;
  assign t_r28_c35_8 = t_r28_c35_4 + p_29_34;
  assign t_r28_c35_9 = t_r28_c35_5 + t_r28_c35_6;
  assign t_r28_c35_10 = t_r28_c35_7 + t_r28_c35_8;
  assign t_r28_c35_11 = t_r28_c35_9 + t_r28_c35_10;
  assign t_r28_c35_12 = t_r28_c35_11 + p_29_36;
  assign out_28_35 = t_r28_c35_12 >> 4;

  assign t_r28_c36_0 = p_27_36 << 1;
  assign t_r28_c36_1 = p_28_35 << 1;
  assign t_r28_c36_2 = p_28_36 << 2;
  assign t_r28_c36_3 = p_28_37 << 1;
  assign t_r28_c36_4 = p_29_36 << 1;
  assign t_r28_c36_5 = t_r28_c36_0 + p_27_35;
  assign t_r28_c36_6 = t_r28_c36_1 + p_27_37;
  assign t_r28_c36_7 = t_r28_c36_2 + t_r28_c36_3;
  assign t_r28_c36_8 = t_r28_c36_4 + p_29_35;
  assign t_r28_c36_9 = t_r28_c36_5 + t_r28_c36_6;
  assign t_r28_c36_10 = t_r28_c36_7 + t_r28_c36_8;
  assign t_r28_c36_11 = t_r28_c36_9 + t_r28_c36_10;
  assign t_r28_c36_12 = t_r28_c36_11 + p_29_37;
  assign out_28_36 = t_r28_c36_12 >> 4;

  assign t_r28_c37_0 = p_27_37 << 1;
  assign t_r28_c37_1 = p_28_36 << 1;
  assign t_r28_c37_2 = p_28_37 << 2;
  assign t_r28_c37_3 = p_28_38 << 1;
  assign t_r28_c37_4 = p_29_37 << 1;
  assign t_r28_c37_5 = t_r28_c37_0 + p_27_36;
  assign t_r28_c37_6 = t_r28_c37_1 + p_27_38;
  assign t_r28_c37_7 = t_r28_c37_2 + t_r28_c37_3;
  assign t_r28_c37_8 = t_r28_c37_4 + p_29_36;
  assign t_r28_c37_9 = t_r28_c37_5 + t_r28_c37_6;
  assign t_r28_c37_10 = t_r28_c37_7 + t_r28_c37_8;
  assign t_r28_c37_11 = t_r28_c37_9 + t_r28_c37_10;
  assign t_r28_c37_12 = t_r28_c37_11 + p_29_38;
  assign out_28_37 = t_r28_c37_12 >> 4;

  assign t_r28_c38_0 = p_27_38 << 1;
  assign t_r28_c38_1 = p_28_37 << 1;
  assign t_r28_c38_2 = p_28_38 << 2;
  assign t_r28_c38_3 = p_28_39 << 1;
  assign t_r28_c38_4 = p_29_38 << 1;
  assign t_r28_c38_5 = t_r28_c38_0 + p_27_37;
  assign t_r28_c38_6 = t_r28_c38_1 + p_27_39;
  assign t_r28_c38_7 = t_r28_c38_2 + t_r28_c38_3;
  assign t_r28_c38_8 = t_r28_c38_4 + p_29_37;
  assign t_r28_c38_9 = t_r28_c38_5 + t_r28_c38_6;
  assign t_r28_c38_10 = t_r28_c38_7 + t_r28_c38_8;
  assign t_r28_c38_11 = t_r28_c38_9 + t_r28_c38_10;
  assign t_r28_c38_12 = t_r28_c38_11 + p_29_39;
  assign out_28_38 = t_r28_c38_12 >> 4;

  assign t_r28_c39_0 = p_27_39 << 1;
  assign t_r28_c39_1 = p_28_38 << 1;
  assign t_r28_c39_2 = p_28_39 << 2;
  assign t_r28_c39_3 = p_28_40 << 1;
  assign t_r28_c39_4 = p_29_39 << 1;
  assign t_r28_c39_5 = t_r28_c39_0 + p_27_38;
  assign t_r28_c39_6 = t_r28_c39_1 + p_27_40;
  assign t_r28_c39_7 = t_r28_c39_2 + t_r28_c39_3;
  assign t_r28_c39_8 = t_r28_c39_4 + p_29_38;
  assign t_r28_c39_9 = t_r28_c39_5 + t_r28_c39_6;
  assign t_r28_c39_10 = t_r28_c39_7 + t_r28_c39_8;
  assign t_r28_c39_11 = t_r28_c39_9 + t_r28_c39_10;
  assign t_r28_c39_12 = t_r28_c39_11 + p_29_40;
  assign out_28_39 = t_r28_c39_12 >> 4;

  assign t_r28_c40_0 = p_27_40 << 1;
  assign t_r28_c40_1 = p_28_39 << 1;
  assign t_r28_c40_2 = p_28_40 << 2;
  assign t_r28_c40_3 = p_28_41 << 1;
  assign t_r28_c40_4 = p_29_40 << 1;
  assign t_r28_c40_5 = t_r28_c40_0 + p_27_39;
  assign t_r28_c40_6 = t_r28_c40_1 + p_27_41;
  assign t_r28_c40_7 = t_r28_c40_2 + t_r28_c40_3;
  assign t_r28_c40_8 = t_r28_c40_4 + p_29_39;
  assign t_r28_c40_9 = t_r28_c40_5 + t_r28_c40_6;
  assign t_r28_c40_10 = t_r28_c40_7 + t_r28_c40_8;
  assign t_r28_c40_11 = t_r28_c40_9 + t_r28_c40_10;
  assign t_r28_c40_12 = t_r28_c40_11 + p_29_41;
  assign out_28_40 = t_r28_c40_12 >> 4;

  assign t_r28_c41_0 = p_27_41 << 1;
  assign t_r28_c41_1 = p_28_40 << 1;
  assign t_r28_c41_2 = p_28_41 << 2;
  assign t_r28_c41_3 = p_28_42 << 1;
  assign t_r28_c41_4 = p_29_41 << 1;
  assign t_r28_c41_5 = t_r28_c41_0 + p_27_40;
  assign t_r28_c41_6 = t_r28_c41_1 + p_27_42;
  assign t_r28_c41_7 = t_r28_c41_2 + t_r28_c41_3;
  assign t_r28_c41_8 = t_r28_c41_4 + p_29_40;
  assign t_r28_c41_9 = t_r28_c41_5 + t_r28_c41_6;
  assign t_r28_c41_10 = t_r28_c41_7 + t_r28_c41_8;
  assign t_r28_c41_11 = t_r28_c41_9 + t_r28_c41_10;
  assign t_r28_c41_12 = t_r28_c41_11 + p_29_42;
  assign out_28_41 = t_r28_c41_12 >> 4;

  assign t_r28_c42_0 = p_27_42 << 1;
  assign t_r28_c42_1 = p_28_41 << 1;
  assign t_r28_c42_2 = p_28_42 << 2;
  assign t_r28_c42_3 = p_28_43 << 1;
  assign t_r28_c42_4 = p_29_42 << 1;
  assign t_r28_c42_5 = t_r28_c42_0 + p_27_41;
  assign t_r28_c42_6 = t_r28_c42_1 + p_27_43;
  assign t_r28_c42_7 = t_r28_c42_2 + t_r28_c42_3;
  assign t_r28_c42_8 = t_r28_c42_4 + p_29_41;
  assign t_r28_c42_9 = t_r28_c42_5 + t_r28_c42_6;
  assign t_r28_c42_10 = t_r28_c42_7 + t_r28_c42_8;
  assign t_r28_c42_11 = t_r28_c42_9 + t_r28_c42_10;
  assign t_r28_c42_12 = t_r28_c42_11 + p_29_43;
  assign out_28_42 = t_r28_c42_12 >> 4;

  assign t_r28_c43_0 = p_27_43 << 1;
  assign t_r28_c43_1 = p_28_42 << 1;
  assign t_r28_c43_2 = p_28_43 << 2;
  assign t_r28_c43_3 = p_28_44 << 1;
  assign t_r28_c43_4 = p_29_43 << 1;
  assign t_r28_c43_5 = t_r28_c43_0 + p_27_42;
  assign t_r28_c43_6 = t_r28_c43_1 + p_27_44;
  assign t_r28_c43_7 = t_r28_c43_2 + t_r28_c43_3;
  assign t_r28_c43_8 = t_r28_c43_4 + p_29_42;
  assign t_r28_c43_9 = t_r28_c43_5 + t_r28_c43_6;
  assign t_r28_c43_10 = t_r28_c43_7 + t_r28_c43_8;
  assign t_r28_c43_11 = t_r28_c43_9 + t_r28_c43_10;
  assign t_r28_c43_12 = t_r28_c43_11 + p_29_44;
  assign out_28_43 = t_r28_c43_12 >> 4;

  assign t_r28_c44_0 = p_27_44 << 1;
  assign t_r28_c44_1 = p_28_43 << 1;
  assign t_r28_c44_2 = p_28_44 << 2;
  assign t_r28_c44_3 = p_28_45 << 1;
  assign t_r28_c44_4 = p_29_44 << 1;
  assign t_r28_c44_5 = t_r28_c44_0 + p_27_43;
  assign t_r28_c44_6 = t_r28_c44_1 + p_27_45;
  assign t_r28_c44_7 = t_r28_c44_2 + t_r28_c44_3;
  assign t_r28_c44_8 = t_r28_c44_4 + p_29_43;
  assign t_r28_c44_9 = t_r28_c44_5 + t_r28_c44_6;
  assign t_r28_c44_10 = t_r28_c44_7 + t_r28_c44_8;
  assign t_r28_c44_11 = t_r28_c44_9 + t_r28_c44_10;
  assign t_r28_c44_12 = t_r28_c44_11 + p_29_45;
  assign out_28_44 = t_r28_c44_12 >> 4;

  assign t_r28_c45_0 = p_27_45 << 1;
  assign t_r28_c45_1 = p_28_44 << 1;
  assign t_r28_c45_2 = p_28_45 << 2;
  assign t_r28_c45_3 = p_28_46 << 1;
  assign t_r28_c45_4 = p_29_45 << 1;
  assign t_r28_c45_5 = t_r28_c45_0 + p_27_44;
  assign t_r28_c45_6 = t_r28_c45_1 + p_27_46;
  assign t_r28_c45_7 = t_r28_c45_2 + t_r28_c45_3;
  assign t_r28_c45_8 = t_r28_c45_4 + p_29_44;
  assign t_r28_c45_9 = t_r28_c45_5 + t_r28_c45_6;
  assign t_r28_c45_10 = t_r28_c45_7 + t_r28_c45_8;
  assign t_r28_c45_11 = t_r28_c45_9 + t_r28_c45_10;
  assign t_r28_c45_12 = t_r28_c45_11 + p_29_46;
  assign out_28_45 = t_r28_c45_12 >> 4;

  assign t_r28_c46_0 = p_27_46 << 1;
  assign t_r28_c46_1 = p_28_45 << 1;
  assign t_r28_c46_2 = p_28_46 << 2;
  assign t_r28_c46_3 = p_28_47 << 1;
  assign t_r28_c46_4 = p_29_46 << 1;
  assign t_r28_c46_5 = t_r28_c46_0 + p_27_45;
  assign t_r28_c46_6 = t_r28_c46_1 + p_27_47;
  assign t_r28_c46_7 = t_r28_c46_2 + t_r28_c46_3;
  assign t_r28_c46_8 = t_r28_c46_4 + p_29_45;
  assign t_r28_c46_9 = t_r28_c46_5 + t_r28_c46_6;
  assign t_r28_c46_10 = t_r28_c46_7 + t_r28_c46_8;
  assign t_r28_c46_11 = t_r28_c46_9 + t_r28_c46_10;
  assign t_r28_c46_12 = t_r28_c46_11 + p_29_47;
  assign out_28_46 = t_r28_c46_12 >> 4;

  assign t_r28_c47_0 = p_27_47 << 1;
  assign t_r28_c47_1 = p_28_46 << 1;
  assign t_r28_c47_2 = p_28_47 << 2;
  assign t_r28_c47_3 = p_28_48 << 1;
  assign t_r28_c47_4 = p_29_47 << 1;
  assign t_r28_c47_5 = t_r28_c47_0 + p_27_46;
  assign t_r28_c47_6 = t_r28_c47_1 + p_27_48;
  assign t_r28_c47_7 = t_r28_c47_2 + t_r28_c47_3;
  assign t_r28_c47_8 = t_r28_c47_4 + p_29_46;
  assign t_r28_c47_9 = t_r28_c47_5 + t_r28_c47_6;
  assign t_r28_c47_10 = t_r28_c47_7 + t_r28_c47_8;
  assign t_r28_c47_11 = t_r28_c47_9 + t_r28_c47_10;
  assign t_r28_c47_12 = t_r28_c47_11 + p_29_48;
  assign out_28_47 = t_r28_c47_12 >> 4;

  assign t_r28_c48_0 = p_27_48 << 1;
  assign t_r28_c48_1 = p_28_47 << 1;
  assign t_r28_c48_2 = p_28_48 << 2;
  assign t_r28_c48_3 = p_28_49 << 1;
  assign t_r28_c48_4 = p_29_48 << 1;
  assign t_r28_c48_5 = t_r28_c48_0 + p_27_47;
  assign t_r28_c48_6 = t_r28_c48_1 + p_27_49;
  assign t_r28_c48_7 = t_r28_c48_2 + t_r28_c48_3;
  assign t_r28_c48_8 = t_r28_c48_4 + p_29_47;
  assign t_r28_c48_9 = t_r28_c48_5 + t_r28_c48_6;
  assign t_r28_c48_10 = t_r28_c48_7 + t_r28_c48_8;
  assign t_r28_c48_11 = t_r28_c48_9 + t_r28_c48_10;
  assign t_r28_c48_12 = t_r28_c48_11 + p_29_49;
  assign out_28_48 = t_r28_c48_12 >> 4;

  assign t_r28_c49_0 = p_27_49 << 1;
  assign t_r28_c49_1 = p_28_48 << 1;
  assign t_r28_c49_2 = p_28_49 << 2;
  assign t_r28_c49_3 = p_28_50 << 1;
  assign t_r28_c49_4 = p_29_49 << 1;
  assign t_r28_c49_5 = t_r28_c49_0 + p_27_48;
  assign t_r28_c49_6 = t_r28_c49_1 + p_27_50;
  assign t_r28_c49_7 = t_r28_c49_2 + t_r28_c49_3;
  assign t_r28_c49_8 = t_r28_c49_4 + p_29_48;
  assign t_r28_c49_9 = t_r28_c49_5 + t_r28_c49_6;
  assign t_r28_c49_10 = t_r28_c49_7 + t_r28_c49_8;
  assign t_r28_c49_11 = t_r28_c49_9 + t_r28_c49_10;
  assign t_r28_c49_12 = t_r28_c49_11 + p_29_50;
  assign out_28_49 = t_r28_c49_12 >> 4;

  assign t_r28_c50_0 = p_27_50 << 1;
  assign t_r28_c50_1 = p_28_49 << 1;
  assign t_r28_c50_2 = p_28_50 << 2;
  assign t_r28_c50_3 = p_28_51 << 1;
  assign t_r28_c50_4 = p_29_50 << 1;
  assign t_r28_c50_5 = t_r28_c50_0 + p_27_49;
  assign t_r28_c50_6 = t_r28_c50_1 + p_27_51;
  assign t_r28_c50_7 = t_r28_c50_2 + t_r28_c50_3;
  assign t_r28_c50_8 = t_r28_c50_4 + p_29_49;
  assign t_r28_c50_9 = t_r28_c50_5 + t_r28_c50_6;
  assign t_r28_c50_10 = t_r28_c50_7 + t_r28_c50_8;
  assign t_r28_c50_11 = t_r28_c50_9 + t_r28_c50_10;
  assign t_r28_c50_12 = t_r28_c50_11 + p_29_51;
  assign out_28_50 = t_r28_c50_12 >> 4;

  assign t_r28_c51_0 = p_27_51 << 1;
  assign t_r28_c51_1 = p_28_50 << 1;
  assign t_r28_c51_2 = p_28_51 << 2;
  assign t_r28_c51_3 = p_28_52 << 1;
  assign t_r28_c51_4 = p_29_51 << 1;
  assign t_r28_c51_5 = t_r28_c51_0 + p_27_50;
  assign t_r28_c51_6 = t_r28_c51_1 + p_27_52;
  assign t_r28_c51_7 = t_r28_c51_2 + t_r28_c51_3;
  assign t_r28_c51_8 = t_r28_c51_4 + p_29_50;
  assign t_r28_c51_9 = t_r28_c51_5 + t_r28_c51_6;
  assign t_r28_c51_10 = t_r28_c51_7 + t_r28_c51_8;
  assign t_r28_c51_11 = t_r28_c51_9 + t_r28_c51_10;
  assign t_r28_c51_12 = t_r28_c51_11 + p_29_52;
  assign out_28_51 = t_r28_c51_12 >> 4;

  assign t_r28_c52_0 = p_27_52 << 1;
  assign t_r28_c52_1 = p_28_51 << 1;
  assign t_r28_c52_2 = p_28_52 << 2;
  assign t_r28_c52_3 = p_28_53 << 1;
  assign t_r28_c52_4 = p_29_52 << 1;
  assign t_r28_c52_5 = t_r28_c52_0 + p_27_51;
  assign t_r28_c52_6 = t_r28_c52_1 + p_27_53;
  assign t_r28_c52_7 = t_r28_c52_2 + t_r28_c52_3;
  assign t_r28_c52_8 = t_r28_c52_4 + p_29_51;
  assign t_r28_c52_9 = t_r28_c52_5 + t_r28_c52_6;
  assign t_r28_c52_10 = t_r28_c52_7 + t_r28_c52_8;
  assign t_r28_c52_11 = t_r28_c52_9 + t_r28_c52_10;
  assign t_r28_c52_12 = t_r28_c52_11 + p_29_53;
  assign out_28_52 = t_r28_c52_12 >> 4;

  assign t_r28_c53_0 = p_27_53 << 1;
  assign t_r28_c53_1 = p_28_52 << 1;
  assign t_r28_c53_2 = p_28_53 << 2;
  assign t_r28_c53_3 = p_28_54 << 1;
  assign t_r28_c53_4 = p_29_53 << 1;
  assign t_r28_c53_5 = t_r28_c53_0 + p_27_52;
  assign t_r28_c53_6 = t_r28_c53_1 + p_27_54;
  assign t_r28_c53_7 = t_r28_c53_2 + t_r28_c53_3;
  assign t_r28_c53_8 = t_r28_c53_4 + p_29_52;
  assign t_r28_c53_9 = t_r28_c53_5 + t_r28_c53_6;
  assign t_r28_c53_10 = t_r28_c53_7 + t_r28_c53_8;
  assign t_r28_c53_11 = t_r28_c53_9 + t_r28_c53_10;
  assign t_r28_c53_12 = t_r28_c53_11 + p_29_54;
  assign out_28_53 = t_r28_c53_12 >> 4;

  assign t_r28_c54_0 = p_27_54 << 1;
  assign t_r28_c54_1 = p_28_53 << 1;
  assign t_r28_c54_2 = p_28_54 << 2;
  assign t_r28_c54_3 = p_28_55 << 1;
  assign t_r28_c54_4 = p_29_54 << 1;
  assign t_r28_c54_5 = t_r28_c54_0 + p_27_53;
  assign t_r28_c54_6 = t_r28_c54_1 + p_27_55;
  assign t_r28_c54_7 = t_r28_c54_2 + t_r28_c54_3;
  assign t_r28_c54_8 = t_r28_c54_4 + p_29_53;
  assign t_r28_c54_9 = t_r28_c54_5 + t_r28_c54_6;
  assign t_r28_c54_10 = t_r28_c54_7 + t_r28_c54_8;
  assign t_r28_c54_11 = t_r28_c54_9 + t_r28_c54_10;
  assign t_r28_c54_12 = t_r28_c54_11 + p_29_55;
  assign out_28_54 = t_r28_c54_12 >> 4;

  assign t_r28_c55_0 = p_27_55 << 1;
  assign t_r28_c55_1 = p_28_54 << 1;
  assign t_r28_c55_2 = p_28_55 << 2;
  assign t_r28_c55_3 = p_28_56 << 1;
  assign t_r28_c55_4 = p_29_55 << 1;
  assign t_r28_c55_5 = t_r28_c55_0 + p_27_54;
  assign t_r28_c55_6 = t_r28_c55_1 + p_27_56;
  assign t_r28_c55_7 = t_r28_c55_2 + t_r28_c55_3;
  assign t_r28_c55_8 = t_r28_c55_4 + p_29_54;
  assign t_r28_c55_9 = t_r28_c55_5 + t_r28_c55_6;
  assign t_r28_c55_10 = t_r28_c55_7 + t_r28_c55_8;
  assign t_r28_c55_11 = t_r28_c55_9 + t_r28_c55_10;
  assign t_r28_c55_12 = t_r28_c55_11 + p_29_56;
  assign out_28_55 = t_r28_c55_12 >> 4;

  assign t_r28_c56_0 = p_27_56 << 1;
  assign t_r28_c56_1 = p_28_55 << 1;
  assign t_r28_c56_2 = p_28_56 << 2;
  assign t_r28_c56_3 = p_28_57 << 1;
  assign t_r28_c56_4 = p_29_56 << 1;
  assign t_r28_c56_5 = t_r28_c56_0 + p_27_55;
  assign t_r28_c56_6 = t_r28_c56_1 + p_27_57;
  assign t_r28_c56_7 = t_r28_c56_2 + t_r28_c56_3;
  assign t_r28_c56_8 = t_r28_c56_4 + p_29_55;
  assign t_r28_c56_9 = t_r28_c56_5 + t_r28_c56_6;
  assign t_r28_c56_10 = t_r28_c56_7 + t_r28_c56_8;
  assign t_r28_c56_11 = t_r28_c56_9 + t_r28_c56_10;
  assign t_r28_c56_12 = t_r28_c56_11 + p_29_57;
  assign out_28_56 = t_r28_c56_12 >> 4;

  assign t_r28_c57_0 = p_27_57 << 1;
  assign t_r28_c57_1 = p_28_56 << 1;
  assign t_r28_c57_2 = p_28_57 << 2;
  assign t_r28_c57_3 = p_28_58 << 1;
  assign t_r28_c57_4 = p_29_57 << 1;
  assign t_r28_c57_5 = t_r28_c57_0 + p_27_56;
  assign t_r28_c57_6 = t_r28_c57_1 + p_27_58;
  assign t_r28_c57_7 = t_r28_c57_2 + t_r28_c57_3;
  assign t_r28_c57_8 = t_r28_c57_4 + p_29_56;
  assign t_r28_c57_9 = t_r28_c57_5 + t_r28_c57_6;
  assign t_r28_c57_10 = t_r28_c57_7 + t_r28_c57_8;
  assign t_r28_c57_11 = t_r28_c57_9 + t_r28_c57_10;
  assign t_r28_c57_12 = t_r28_c57_11 + p_29_58;
  assign out_28_57 = t_r28_c57_12 >> 4;

  assign t_r28_c58_0 = p_27_58 << 1;
  assign t_r28_c58_1 = p_28_57 << 1;
  assign t_r28_c58_2 = p_28_58 << 2;
  assign t_r28_c58_3 = p_28_59 << 1;
  assign t_r28_c58_4 = p_29_58 << 1;
  assign t_r28_c58_5 = t_r28_c58_0 + p_27_57;
  assign t_r28_c58_6 = t_r28_c58_1 + p_27_59;
  assign t_r28_c58_7 = t_r28_c58_2 + t_r28_c58_3;
  assign t_r28_c58_8 = t_r28_c58_4 + p_29_57;
  assign t_r28_c58_9 = t_r28_c58_5 + t_r28_c58_6;
  assign t_r28_c58_10 = t_r28_c58_7 + t_r28_c58_8;
  assign t_r28_c58_11 = t_r28_c58_9 + t_r28_c58_10;
  assign t_r28_c58_12 = t_r28_c58_11 + p_29_59;
  assign out_28_58 = t_r28_c58_12 >> 4;

  assign t_r28_c59_0 = p_27_59 << 1;
  assign t_r28_c59_1 = p_28_58 << 1;
  assign t_r28_c59_2 = p_28_59 << 2;
  assign t_r28_c59_3 = p_28_60 << 1;
  assign t_r28_c59_4 = p_29_59 << 1;
  assign t_r28_c59_5 = t_r28_c59_0 + p_27_58;
  assign t_r28_c59_6 = t_r28_c59_1 + p_27_60;
  assign t_r28_c59_7 = t_r28_c59_2 + t_r28_c59_3;
  assign t_r28_c59_8 = t_r28_c59_4 + p_29_58;
  assign t_r28_c59_9 = t_r28_c59_5 + t_r28_c59_6;
  assign t_r28_c59_10 = t_r28_c59_7 + t_r28_c59_8;
  assign t_r28_c59_11 = t_r28_c59_9 + t_r28_c59_10;
  assign t_r28_c59_12 = t_r28_c59_11 + p_29_60;
  assign out_28_59 = t_r28_c59_12 >> 4;

  assign t_r28_c60_0 = p_27_60 << 1;
  assign t_r28_c60_1 = p_28_59 << 1;
  assign t_r28_c60_2 = p_28_60 << 2;
  assign t_r28_c60_3 = p_28_61 << 1;
  assign t_r28_c60_4 = p_29_60 << 1;
  assign t_r28_c60_5 = t_r28_c60_0 + p_27_59;
  assign t_r28_c60_6 = t_r28_c60_1 + p_27_61;
  assign t_r28_c60_7 = t_r28_c60_2 + t_r28_c60_3;
  assign t_r28_c60_8 = t_r28_c60_4 + p_29_59;
  assign t_r28_c60_9 = t_r28_c60_5 + t_r28_c60_6;
  assign t_r28_c60_10 = t_r28_c60_7 + t_r28_c60_8;
  assign t_r28_c60_11 = t_r28_c60_9 + t_r28_c60_10;
  assign t_r28_c60_12 = t_r28_c60_11 + p_29_61;
  assign out_28_60 = t_r28_c60_12 >> 4;

  assign t_r28_c61_0 = p_27_61 << 1;
  assign t_r28_c61_1 = p_28_60 << 1;
  assign t_r28_c61_2 = p_28_61 << 2;
  assign t_r28_c61_3 = p_28_62 << 1;
  assign t_r28_c61_4 = p_29_61 << 1;
  assign t_r28_c61_5 = t_r28_c61_0 + p_27_60;
  assign t_r28_c61_6 = t_r28_c61_1 + p_27_62;
  assign t_r28_c61_7 = t_r28_c61_2 + t_r28_c61_3;
  assign t_r28_c61_8 = t_r28_c61_4 + p_29_60;
  assign t_r28_c61_9 = t_r28_c61_5 + t_r28_c61_6;
  assign t_r28_c61_10 = t_r28_c61_7 + t_r28_c61_8;
  assign t_r28_c61_11 = t_r28_c61_9 + t_r28_c61_10;
  assign t_r28_c61_12 = t_r28_c61_11 + p_29_62;
  assign out_28_61 = t_r28_c61_12 >> 4;

  assign t_r28_c62_0 = p_27_62 << 1;
  assign t_r28_c62_1 = p_28_61 << 1;
  assign t_r28_c62_2 = p_28_62 << 2;
  assign t_r28_c62_3 = p_28_63 << 1;
  assign t_r28_c62_4 = p_29_62 << 1;
  assign t_r28_c62_5 = t_r28_c62_0 + p_27_61;
  assign t_r28_c62_6 = t_r28_c62_1 + p_27_63;
  assign t_r28_c62_7 = t_r28_c62_2 + t_r28_c62_3;
  assign t_r28_c62_8 = t_r28_c62_4 + p_29_61;
  assign t_r28_c62_9 = t_r28_c62_5 + t_r28_c62_6;
  assign t_r28_c62_10 = t_r28_c62_7 + t_r28_c62_8;
  assign t_r28_c62_11 = t_r28_c62_9 + t_r28_c62_10;
  assign t_r28_c62_12 = t_r28_c62_11 + p_29_63;
  assign out_28_62 = t_r28_c62_12 >> 4;

  assign t_r28_c63_0 = p_27_63 << 1;
  assign t_r28_c63_1 = p_28_62 << 1;
  assign t_r28_c63_2 = p_28_63 << 2;
  assign t_r28_c63_3 = p_28_64 << 1;
  assign t_r28_c63_4 = p_29_63 << 1;
  assign t_r28_c63_5 = t_r28_c63_0 + p_27_62;
  assign t_r28_c63_6 = t_r28_c63_1 + p_27_64;
  assign t_r28_c63_7 = t_r28_c63_2 + t_r28_c63_3;
  assign t_r28_c63_8 = t_r28_c63_4 + p_29_62;
  assign t_r28_c63_9 = t_r28_c63_5 + t_r28_c63_6;
  assign t_r28_c63_10 = t_r28_c63_7 + t_r28_c63_8;
  assign t_r28_c63_11 = t_r28_c63_9 + t_r28_c63_10;
  assign t_r28_c63_12 = t_r28_c63_11 + p_29_64;
  assign out_28_63 = t_r28_c63_12 >> 4;

  assign t_r28_c64_0 = p_27_64 << 1;
  assign t_r28_c64_1 = p_28_63 << 1;
  assign t_r28_c64_2 = p_28_64 << 2;
  assign t_r28_c64_3 = p_28_65 << 1;
  assign t_r28_c64_4 = p_29_64 << 1;
  assign t_r28_c64_5 = t_r28_c64_0 + p_27_63;
  assign t_r28_c64_6 = t_r28_c64_1 + p_27_65;
  assign t_r28_c64_7 = t_r28_c64_2 + t_r28_c64_3;
  assign t_r28_c64_8 = t_r28_c64_4 + p_29_63;
  assign t_r28_c64_9 = t_r28_c64_5 + t_r28_c64_6;
  assign t_r28_c64_10 = t_r28_c64_7 + t_r28_c64_8;
  assign t_r28_c64_11 = t_r28_c64_9 + t_r28_c64_10;
  assign t_r28_c64_12 = t_r28_c64_11 + p_29_65;
  assign out_28_64 = t_r28_c64_12 >> 4;

  assign t_r29_c1_0 = p_28_1 << 1;
  assign t_r29_c1_1 = p_29_0 << 1;
  assign t_r29_c1_2 = p_29_1 << 2;
  assign t_r29_c1_3 = p_29_2 << 1;
  assign t_r29_c1_4 = p_30_1 << 1;
  assign t_r29_c1_5 = t_r29_c1_0 + p_28_0;
  assign t_r29_c1_6 = t_r29_c1_1 + p_28_2;
  assign t_r29_c1_7 = t_r29_c1_2 + t_r29_c1_3;
  assign t_r29_c1_8 = t_r29_c1_4 + p_30_0;
  assign t_r29_c1_9 = t_r29_c1_5 + t_r29_c1_6;
  assign t_r29_c1_10 = t_r29_c1_7 + t_r29_c1_8;
  assign t_r29_c1_11 = t_r29_c1_9 + t_r29_c1_10;
  assign t_r29_c1_12 = t_r29_c1_11 + p_30_2;
  assign out_29_1 = t_r29_c1_12 >> 4;

  assign t_r29_c2_0 = p_28_2 << 1;
  assign t_r29_c2_1 = p_29_1 << 1;
  assign t_r29_c2_2 = p_29_2 << 2;
  assign t_r29_c2_3 = p_29_3 << 1;
  assign t_r29_c2_4 = p_30_2 << 1;
  assign t_r29_c2_5 = t_r29_c2_0 + p_28_1;
  assign t_r29_c2_6 = t_r29_c2_1 + p_28_3;
  assign t_r29_c2_7 = t_r29_c2_2 + t_r29_c2_3;
  assign t_r29_c2_8 = t_r29_c2_4 + p_30_1;
  assign t_r29_c2_9 = t_r29_c2_5 + t_r29_c2_6;
  assign t_r29_c2_10 = t_r29_c2_7 + t_r29_c2_8;
  assign t_r29_c2_11 = t_r29_c2_9 + t_r29_c2_10;
  assign t_r29_c2_12 = t_r29_c2_11 + p_30_3;
  assign out_29_2 = t_r29_c2_12 >> 4;

  assign t_r29_c3_0 = p_28_3 << 1;
  assign t_r29_c3_1 = p_29_2 << 1;
  assign t_r29_c3_2 = p_29_3 << 2;
  assign t_r29_c3_3 = p_29_4 << 1;
  assign t_r29_c3_4 = p_30_3 << 1;
  assign t_r29_c3_5 = t_r29_c3_0 + p_28_2;
  assign t_r29_c3_6 = t_r29_c3_1 + p_28_4;
  assign t_r29_c3_7 = t_r29_c3_2 + t_r29_c3_3;
  assign t_r29_c3_8 = t_r29_c3_4 + p_30_2;
  assign t_r29_c3_9 = t_r29_c3_5 + t_r29_c3_6;
  assign t_r29_c3_10 = t_r29_c3_7 + t_r29_c3_8;
  assign t_r29_c3_11 = t_r29_c3_9 + t_r29_c3_10;
  assign t_r29_c3_12 = t_r29_c3_11 + p_30_4;
  assign out_29_3 = t_r29_c3_12 >> 4;

  assign t_r29_c4_0 = p_28_4 << 1;
  assign t_r29_c4_1 = p_29_3 << 1;
  assign t_r29_c4_2 = p_29_4 << 2;
  assign t_r29_c4_3 = p_29_5 << 1;
  assign t_r29_c4_4 = p_30_4 << 1;
  assign t_r29_c4_5 = t_r29_c4_0 + p_28_3;
  assign t_r29_c4_6 = t_r29_c4_1 + p_28_5;
  assign t_r29_c4_7 = t_r29_c4_2 + t_r29_c4_3;
  assign t_r29_c4_8 = t_r29_c4_4 + p_30_3;
  assign t_r29_c4_9 = t_r29_c4_5 + t_r29_c4_6;
  assign t_r29_c4_10 = t_r29_c4_7 + t_r29_c4_8;
  assign t_r29_c4_11 = t_r29_c4_9 + t_r29_c4_10;
  assign t_r29_c4_12 = t_r29_c4_11 + p_30_5;
  assign out_29_4 = t_r29_c4_12 >> 4;

  assign t_r29_c5_0 = p_28_5 << 1;
  assign t_r29_c5_1 = p_29_4 << 1;
  assign t_r29_c5_2 = p_29_5 << 2;
  assign t_r29_c5_3 = p_29_6 << 1;
  assign t_r29_c5_4 = p_30_5 << 1;
  assign t_r29_c5_5 = t_r29_c5_0 + p_28_4;
  assign t_r29_c5_6 = t_r29_c5_1 + p_28_6;
  assign t_r29_c5_7 = t_r29_c5_2 + t_r29_c5_3;
  assign t_r29_c5_8 = t_r29_c5_4 + p_30_4;
  assign t_r29_c5_9 = t_r29_c5_5 + t_r29_c5_6;
  assign t_r29_c5_10 = t_r29_c5_7 + t_r29_c5_8;
  assign t_r29_c5_11 = t_r29_c5_9 + t_r29_c5_10;
  assign t_r29_c5_12 = t_r29_c5_11 + p_30_6;
  assign out_29_5 = t_r29_c5_12 >> 4;

  assign t_r29_c6_0 = p_28_6 << 1;
  assign t_r29_c6_1 = p_29_5 << 1;
  assign t_r29_c6_2 = p_29_6 << 2;
  assign t_r29_c6_3 = p_29_7 << 1;
  assign t_r29_c6_4 = p_30_6 << 1;
  assign t_r29_c6_5 = t_r29_c6_0 + p_28_5;
  assign t_r29_c6_6 = t_r29_c6_1 + p_28_7;
  assign t_r29_c6_7 = t_r29_c6_2 + t_r29_c6_3;
  assign t_r29_c6_8 = t_r29_c6_4 + p_30_5;
  assign t_r29_c6_9 = t_r29_c6_5 + t_r29_c6_6;
  assign t_r29_c6_10 = t_r29_c6_7 + t_r29_c6_8;
  assign t_r29_c6_11 = t_r29_c6_9 + t_r29_c6_10;
  assign t_r29_c6_12 = t_r29_c6_11 + p_30_7;
  assign out_29_6 = t_r29_c6_12 >> 4;

  assign t_r29_c7_0 = p_28_7 << 1;
  assign t_r29_c7_1 = p_29_6 << 1;
  assign t_r29_c7_2 = p_29_7 << 2;
  assign t_r29_c7_3 = p_29_8 << 1;
  assign t_r29_c7_4 = p_30_7 << 1;
  assign t_r29_c7_5 = t_r29_c7_0 + p_28_6;
  assign t_r29_c7_6 = t_r29_c7_1 + p_28_8;
  assign t_r29_c7_7 = t_r29_c7_2 + t_r29_c7_3;
  assign t_r29_c7_8 = t_r29_c7_4 + p_30_6;
  assign t_r29_c7_9 = t_r29_c7_5 + t_r29_c7_6;
  assign t_r29_c7_10 = t_r29_c7_7 + t_r29_c7_8;
  assign t_r29_c7_11 = t_r29_c7_9 + t_r29_c7_10;
  assign t_r29_c7_12 = t_r29_c7_11 + p_30_8;
  assign out_29_7 = t_r29_c7_12 >> 4;

  assign t_r29_c8_0 = p_28_8 << 1;
  assign t_r29_c8_1 = p_29_7 << 1;
  assign t_r29_c8_2 = p_29_8 << 2;
  assign t_r29_c8_3 = p_29_9 << 1;
  assign t_r29_c8_4 = p_30_8 << 1;
  assign t_r29_c8_5 = t_r29_c8_0 + p_28_7;
  assign t_r29_c8_6 = t_r29_c8_1 + p_28_9;
  assign t_r29_c8_7 = t_r29_c8_2 + t_r29_c8_3;
  assign t_r29_c8_8 = t_r29_c8_4 + p_30_7;
  assign t_r29_c8_9 = t_r29_c8_5 + t_r29_c8_6;
  assign t_r29_c8_10 = t_r29_c8_7 + t_r29_c8_8;
  assign t_r29_c8_11 = t_r29_c8_9 + t_r29_c8_10;
  assign t_r29_c8_12 = t_r29_c8_11 + p_30_9;
  assign out_29_8 = t_r29_c8_12 >> 4;

  assign t_r29_c9_0 = p_28_9 << 1;
  assign t_r29_c9_1 = p_29_8 << 1;
  assign t_r29_c9_2 = p_29_9 << 2;
  assign t_r29_c9_3 = p_29_10 << 1;
  assign t_r29_c9_4 = p_30_9 << 1;
  assign t_r29_c9_5 = t_r29_c9_0 + p_28_8;
  assign t_r29_c9_6 = t_r29_c9_1 + p_28_10;
  assign t_r29_c9_7 = t_r29_c9_2 + t_r29_c9_3;
  assign t_r29_c9_8 = t_r29_c9_4 + p_30_8;
  assign t_r29_c9_9 = t_r29_c9_5 + t_r29_c9_6;
  assign t_r29_c9_10 = t_r29_c9_7 + t_r29_c9_8;
  assign t_r29_c9_11 = t_r29_c9_9 + t_r29_c9_10;
  assign t_r29_c9_12 = t_r29_c9_11 + p_30_10;
  assign out_29_9 = t_r29_c9_12 >> 4;

  assign t_r29_c10_0 = p_28_10 << 1;
  assign t_r29_c10_1 = p_29_9 << 1;
  assign t_r29_c10_2 = p_29_10 << 2;
  assign t_r29_c10_3 = p_29_11 << 1;
  assign t_r29_c10_4 = p_30_10 << 1;
  assign t_r29_c10_5 = t_r29_c10_0 + p_28_9;
  assign t_r29_c10_6 = t_r29_c10_1 + p_28_11;
  assign t_r29_c10_7 = t_r29_c10_2 + t_r29_c10_3;
  assign t_r29_c10_8 = t_r29_c10_4 + p_30_9;
  assign t_r29_c10_9 = t_r29_c10_5 + t_r29_c10_6;
  assign t_r29_c10_10 = t_r29_c10_7 + t_r29_c10_8;
  assign t_r29_c10_11 = t_r29_c10_9 + t_r29_c10_10;
  assign t_r29_c10_12 = t_r29_c10_11 + p_30_11;
  assign out_29_10 = t_r29_c10_12 >> 4;

  assign t_r29_c11_0 = p_28_11 << 1;
  assign t_r29_c11_1 = p_29_10 << 1;
  assign t_r29_c11_2 = p_29_11 << 2;
  assign t_r29_c11_3 = p_29_12 << 1;
  assign t_r29_c11_4 = p_30_11 << 1;
  assign t_r29_c11_5 = t_r29_c11_0 + p_28_10;
  assign t_r29_c11_6 = t_r29_c11_1 + p_28_12;
  assign t_r29_c11_7 = t_r29_c11_2 + t_r29_c11_3;
  assign t_r29_c11_8 = t_r29_c11_4 + p_30_10;
  assign t_r29_c11_9 = t_r29_c11_5 + t_r29_c11_6;
  assign t_r29_c11_10 = t_r29_c11_7 + t_r29_c11_8;
  assign t_r29_c11_11 = t_r29_c11_9 + t_r29_c11_10;
  assign t_r29_c11_12 = t_r29_c11_11 + p_30_12;
  assign out_29_11 = t_r29_c11_12 >> 4;

  assign t_r29_c12_0 = p_28_12 << 1;
  assign t_r29_c12_1 = p_29_11 << 1;
  assign t_r29_c12_2 = p_29_12 << 2;
  assign t_r29_c12_3 = p_29_13 << 1;
  assign t_r29_c12_4 = p_30_12 << 1;
  assign t_r29_c12_5 = t_r29_c12_0 + p_28_11;
  assign t_r29_c12_6 = t_r29_c12_1 + p_28_13;
  assign t_r29_c12_7 = t_r29_c12_2 + t_r29_c12_3;
  assign t_r29_c12_8 = t_r29_c12_4 + p_30_11;
  assign t_r29_c12_9 = t_r29_c12_5 + t_r29_c12_6;
  assign t_r29_c12_10 = t_r29_c12_7 + t_r29_c12_8;
  assign t_r29_c12_11 = t_r29_c12_9 + t_r29_c12_10;
  assign t_r29_c12_12 = t_r29_c12_11 + p_30_13;
  assign out_29_12 = t_r29_c12_12 >> 4;

  assign t_r29_c13_0 = p_28_13 << 1;
  assign t_r29_c13_1 = p_29_12 << 1;
  assign t_r29_c13_2 = p_29_13 << 2;
  assign t_r29_c13_3 = p_29_14 << 1;
  assign t_r29_c13_4 = p_30_13 << 1;
  assign t_r29_c13_5 = t_r29_c13_0 + p_28_12;
  assign t_r29_c13_6 = t_r29_c13_1 + p_28_14;
  assign t_r29_c13_7 = t_r29_c13_2 + t_r29_c13_3;
  assign t_r29_c13_8 = t_r29_c13_4 + p_30_12;
  assign t_r29_c13_9 = t_r29_c13_5 + t_r29_c13_6;
  assign t_r29_c13_10 = t_r29_c13_7 + t_r29_c13_8;
  assign t_r29_c13_11 = t_r29_c13_9 + t_r29_c13_10;
  assign t_r29_c13_12 = t_r29_c13_11 + p_30_14;
  assign out_29_13 = t_r29_c13_12 >> 4;

  assign t_r29_c14_0 = p_28_14 << 1;
  assign t_r29_c14_1 = p_29_13 << 1;
  assign t_r29_c14_2 = p_29_14 << 2;
  assign t_r29_c14_3 = p_29_15 << 1;
  assign t_r29_c14_4 = p_30_14 << 1;
  assign t_r29_c14_5 = t_r29_c14_0 + p_28_13;
  assign t_r29_c14_6 = t_r29_c14_1 + p_28_15;
  assign t_r29_c14_7 = t_r29_c14_2 + t_r29_c14_3;
  assign t_r29_c14_8 = t_r29_c14_4 + p_30_13;
  assign t_r29_c14_9 = t_r29_c14_5 + t_r29_c14_6;
  assign t_r29_c14_10 = t_r29_c14_7 + t_r29_c14_8;
  assign t_r29_c14_11 = t_r29_c14_9 + t_r29_c14_10;
  assign t_r29_c14_12 = t_r29_c14_11 + p_30_15;
  assign out_29_14 = t_r29_c14_12 >> 4;

  assign t_r29_c15_0 = p_28_15 << 1;
  assign t_r29_c15_1 = p_29_14 << 1;
  assign t_r29_c15_2 = p_29_15 << 2;
  assign t_r29_c15_3 = p_29_16 << 1;
  assign t_r29_c15_4 = p_30_15 << 1;
  assign t_r29_c15_5 = t_r29_c15_0 + p_28_14;
  assign t_r29_c15_6 = t_r29_c15_1 + p_28_16;
  assign t_r29_c15_7 = t_r29_c15_2 + t_r29_c15_3;
  assign t_r29_c15_8 = t_r29_c15_4 + p_30_14;
  assign t_r29_c15_9 = t_r29_c15_5 + t_r29_c15_6;
  assign t_r29_c15_10 = t_r29_c15_7 + t_r29_c15_8;
  assign t_r29_c15_11 = t_r29_c15_9 + t_r29_c15_10;
  assign t_r29_c15_12 = t_r29_c15_11 + p_30_16;
  assign out_29_15 = t_r29_c15_12 >> 4;

  assign t_r29_c16_0 = p_28_16 << 1;
  assign t_r29_c16_1 = p_29_15 << 1;
  assign t_r29_c16_2 = p_29_16 << 2;
  assign t_r29_c16_3 = p_29_17 << 1;
  assign t_r29_c16_4 = p_30_16 << 1;
  assign t_r29_c16_5 = t_r29_c16_0 + p_28_15;
  assign t_r29_c16_6 = t_r29_c16_1 + p_28_17;
  assign t_r29_c16_7 = t_r29_c16_2 + t_r29_c16_3;
  assign t_r29_c16_8 = t_r29_c16_4 + p_30_15;
  assign t_r29_c16_9 = t_r29_c16_5 + t_r29_c16_6;
  assign t_r29_c16_10 = t_r29_c16_7 + t_r29_c16_8;
  assign t_r29_c16_11 = t_r29_c16_9 + t_r29_c16_10;
  assign t_r29_c16_12 = t_r29_c16_11 + p_30_17;
  assign out_29_16 = t_r29_c16_12 >> 4;

  assign t_r29_c17_0 = p_28_17 << 1;
  assign t_r29_c17_1 = p_29_16 << 1;
  assign t_r29_c17_2 = p_29_17 << 2;
  assign t_r29_c17_3 = p_29_18 << 1;
  assign t_r29_c17_4 = p_30_17 << 1;
  assign t_r29_c17_5 = t_r29_c17_0 + p_28_16;
  assign t_r29_c17_6 = t_r29_c17_1 + p_28_18;
  assign t_r29_c17_7 = t_r29_c17_2 + t_r29_c17_3;
  assign t_r29_c17_8 = t_r29_c17_4 + p_30_16;
  assign t_r29_c17_9 = t_r29_c17_5 + t_r29_c17_6;
  assign t_r29_c17_10 = t_r29_c17_7 + t_r29_c17_8;
  assign t_r29_c17_11 = t_r29_c17_9 + t_r29_c17_10;
  assign t_r29_c17_12 = t_r29_c17_11 + p_30_18;
  assign out_29_17 = t_r29_c17_12 >> 4;

  assign t_r29_c18_0 = p_28_18 << 1;
  assign t_r29_c18_1 = p_29_17 << 1;
  assign t_r29_c18_2 = p_29_18 << 2;
  assign t_r29_c18_3 = p_29_19 << 1;
  assign t_r29_c18_4 = p_30_18 << 1;
  assign t_r29_c18_5 = t_r29_c18_0 + p_28_17;
  assign t_r29_c18_6 = t_r29_c18_1 + p_28_19;
  assign t_r29_c18_7 = t_r29_c18_2 + t_r29_c18_3;
  assign t_r29_c18_8 = t_r29_c18_4 + p_30_17;
  assign t_r29_c18_9 = t_r29_c18_5 + t_r29_c18_6;
  assign t_r29_c18_10 = t_r29_c18_7 + t_r29_c18_8;
  assign t_r29_c18_11 = t_r29_c18_9 + t_r29_c18_10;
  assign t_r29_c18_12 = t_r29_c18_11 + p_30_19;
  assign out_29_18 = t_r29_c18_12 >> 4;

  assign t_r29_c19_0 = p_28_19 << 1;
  assign t_r29_c19_1 = p_29_18 << 1;
  assign t_r29_c19_2 = p_29_19 << 2;
  assign t_r29_c19_3 = p_29_20 << 1;
  assign t_r29_c19_4 = p_30_19 << 1;
  assign t_r29_c19_5 = t_r29_c19_0 + p_28_18;
  assign t_r29_c19_6 = t_r29_c19_1 + p_28_20;
  assign t_r29_c19_7 = t_r29_c19_2 + t_r29_c19_3;
  assign t_r29_c19_8 = t_r29_c19_4 + p_30_18;
  assign t_r29_c19_9 = t_r29_c19_5 + t_r29_c19_6;
  assign t_r29_c19_10 = t_r29_c19_7 + t_r29_c19_8;
  assign t_r29_c19_11 = t_r29_c19_9 + t_r29_c19_10;
  assign t_r29_c19_12 = t_r29_c19_11 + p_30_20;
  assign out_29_19 = t_r29_c19_12 >> 4;

  assign t_r29_c20_0 = p_28_20 << 1;
  assign t_r29_c20_1 = p_29_19 << 1;
  assign t_r29_c20_2 = p_29_20 << 2;
  assign t_r29_c20_3 = p_29_21 << 1;
  assign t_r29_c20_4 = p_30_20 << 1;
  assign t_r29_c20_5 = t_r29_c20_0 + p_28_19;
  assign t_r29_c20_6 = t_r29_c20_1 + p_28_21;
  assign t_r29_c20_7 = t_r29_c20_2 + t_r29_c20_3;
  assign t_r29_c20_8 = t_r29_c20_4 + p_30_19;
  assign t_r29_c20_9 = t_r29_c20_5 + t_r29_c20_6;
  assign t_r29_c20_10 = t_r29_c20_7 + t_r29_c20_8;
  assign t_r29_c20_11 = t_r29_c20_9 + t_r29_c20_10;
  assign t_r29_c20_12 = t_r29_c20_11 + p_30_21;
  assign out_29_20 = t_r29_c20_12 >> 4;

  assign t_r29_c21_0 = p_28_21 << 1;
  assign t_r29_c21_1 = p_29_20 << 1;
  assign t_r29_c21_2 = p_29_21 << 2;
  assign t_r29_c21_3 = p_29_22 << 1;
  assign t_r29_c21_4 = p_30_21 << 1;
  assign t_r29_c21_5 = t_r29_c21_0 + p_28_20;
  assign t_r29_c21_6 = t_r29_c21_1 + p_28_22;
  assign t_r29_c21_7 = t_r29_c21_2 + t_r29_c21_3;
  assign t_r29_c21_8 = t_r29_c21_4 + p_30_20;
  assign t_r29_c21_9 = t_r29_c21_5 + t_r29_c21_6;
  assign t_r29_c21_10 = t_r29_c21_7 + t_r29_c21_8;
  assign t_r29_c21_11 = t_r29_c21_9 + t_r29_c21_10;
  assign t_r29_c21_12 = t_r29_c21_11 + p_30_22;
  assign out_29_21 = t_r29_c21_12 >> 4;

  assign t_r29_c22_0 = p_28_22 << 1;
  assign t_r29_c22_1 = p_29_21 << 1;
  assign t_r29_c22_2 = p_29_22 << 2;
  assign t_r29_c22_3 = p_29_23 << 1;
  assign t_r29_c22_4 = p_30_22 << 1;
  assign t_r29_c22_5 = t_r29_c22_0 + p_28_21;
  assign t_r29_c22_6 = t_r29_c22_1 + p_28_23;
  assign t_r29_c22_7 = t_r29_c22_2 + t_r29_c22_3;
  assign t_r29_c22_8 = t_r29_c22_4 + p_30_21;
  assign t_r29_c22_9 = t_r29_c22_5 + t_r29_c22_6;
  assign t_r29_c22_10 = t_r29_c22_7 + t_r29_c22_8;
  assign t_r29_c22_11 = t_r29_c22_9 + t_r29_c22_10;
  assign t_r29_c22_12 = t_r29_c22_11 + p_30_23;
  assign out_29_22 = t_r29_c22_12 >> 4;

  assign t_r29_c23_0 = p_28_23 << 1;
  assign t_r29_c23_1 = p_29_22 << 1;
  assign t_r29_c23_2 = p_29_23 << 2;
  assign t_r29_c23_3 = p_29_24 << 1;
  assign t_r29_c23_4 = p_30_23 << 1;
  assign t_r29_c23_5 = t_r29_c23_0 + p_28_22;
  assign t_r29_c23_6 = t_r29_c23_1 + p_28_24;
  assign t_r29_c23_7 = t_r29_c23_2 + t_r29_c23_3;
  assign t_r29_c23_8 = t_r29_c23_4 + p_30_22;
  assign t_r29_c23_9 = t_r29_c23_5 + t_r29_c23_6;
  assign t_r29_c23_10 = t_r29_c23_7 + t_r29_c23_8;
  assign t_r29_c23_11 = t_r29_c23_9 + t_r29_c23_10;
  assign t_r29_c23_12 = t_r29_c23_11 + p_30_24;
  assign out_29_23 = t_r29_c23_12 >> 4;

  assign t_r29_c24_0 = p_28_24 << 1;
  assign t_r29_c24_1 = p_29_23 << 1;
  assign t_r29_c24_2 = p_29_24 << 2;
  assign t_r29_c24_3 = p_29_25 << 1;
  assign t_r29_c24_4 = p_30_24 << 1;
  assign t_r29_c24_5 = t_r29_c24_0 + p_28_23;
  assign t_r29_c24_6 = t_r29_c24_1 + p_28_25;
  assign t_r29_c24_7 = t_r29_c24_2 + t_r29_c24_3;
  assign t_r29_c24_8 = t_r29_c24_4 + p_30_23;
  assign t_r29_c24_9 = t_r29_c24_5 + t_r29_c24_6;
  assign t_r29_c24_10 = t_r29_c24_7 + t_r29_c24_8;
  assign t_r29_c24_11 = t_r29_c24_9 + t_r29_c24_10;
  assign t_r29_c24_12 = t_r29_c24_11 + p_30_25;
  assign out_29_24 = t_r29_c24_12 >> 4;

  assign t_r29_c25_0 = p_28_25 << 1;
  assign t_r29_c25_1 = p_29_24 << 1;
  assign t_r29_c25_2 = p_29_25 << 2;
  assign t_r29_c25_3 = p_29_26 << 1;
  assign t_r29_c25_4 = p_30_25 << 1;
  assign t_r29_c25_5 = t_r29_c25_0 + p_28_24;
  assign t_r29_c25_6 = t_r29_c25_1 + p_28_26;
  assign t_r29_c25_7 = t_r29_c25_2 + t_r29_c25_3;
  assign t_r29_c25_8 = t_r29_c25_4 + p_30_24;
  assign t_r29_c25_9 = t_r29_c25_5 + t_r29_c25_6;
  assign t_r29_c25_10 = t_r29_c25_7 + t_r29_c25_8;
  assign t_r29_c25_11 = t_r29_c25_9 + t_r29_c25_10;
  assign t_r29_c25_12 = t_r29_c25_11 + p_30_26;
  assign out_29_25 = t_r29_c25_12 >> 4;

  assign t_r29_c26_0 = p_28_26 << 1;
  assign t_r29_c26_1 = p_29_25 << 1;
  assign t_r29_c26_2 = p_29_26 << 2;
  assign t_r29_c26_3 = p_29_27 << 1;
  assign t_r29_c26_4 = p_30_26 << 1;
  assign t_r29_c26_5 = t_r29_c26_0 + p_28_25;
  assign t_r29_c26_6 = t_r29_c26_1 + p_28_27;
  assign t_r29_c26_7 = t_r29_c26_2 + t_r29_c26_3;
  assign t_r29_c26_8 = t_r29_c26_4 + p_30_25;
  assign t_r29_c26_9 = t_r29_c26_5 + t_r29_c26_6;
  assign t_r29_c26_10 = t_r29_c26_7 + t_r29_c26_8;
  assign t_r29_c26_11 = t_r29_c26_9 + t_r29_c26_10;
  assign t_r29_c26_12 = t_r29_c26_11 + p_30_27;
  assign out_29_26 = t_r29_c26_12 >> 4;

  assign t_r29_c27_0 = p_28_27 << 1;
  assign t_r29_c27_1 = p_29_26 << 1;
  assign t_r29_c27_2 = p_29_27 << 2;
  assign t_r29_c27_3 = p_29_28 << 1;
  assign t_r29_c27_4 = p_30_27 << 1;
  assign t_r29_c27_5 = t_r29_c27_0 + p_28_26;
  assign t_r29_c27_6 = t_r29_c27_1 + p_28_28;
  assign t_r29_c27_7 = t_r29_c27_2 + t_r29_c27_3;
  assign t_r29_c27_8 = t_r29_c27_4 + p_30_26;
  assign t_r29_c27_9 = t_r29_c27_5 + t_r29_c27_6;
  assign t_r29_c27_10 = t_r29_c27_7 + t_r29_c27_8;
  assign t_r29_c27_11 = t_r29_c27_9 + t_r29_c27_10;
  assign t_r29_c27_12 = t_r29_c27_11 + p_30_28;
  assign out_29_27 = t_r29_c27_12 >> 4;

  assign t_r29_c28_0 = p_28_28 << 1;
  assign t_r29_c28_1 = p_29_27 << 1;
  assign t_r29_c28_2 = p_29_28 << 2;
  assign t_r29_c28_3 = p_29_29 << 1;
  assign t_r29_c28_4 = p_30_28 << 1;
  assign t_r29_c28_5 = t_r29_c28_0 + p_28_27;
  assign t_r29_c28_6 = t_r29_c28_1 + p_28_29;
  assign t_r29_c28_7 = t_r29_c28_2 + t_r29_c28_3;
  assign t_r29_c28_8 = t_r29_c28_4 + p_30_27;
  assign t_r29_c28_9 = t_r29_c28_5 + t_r29_c28_6;
  assign t_r29_c28_10 = t_r29_c28_7 + t_r29_c28_8;
  assign t_r29_c28_11 = t_r29_c28_9 + t_r29_c28_10;
  assign t_r29_c28_12 = t_r29_c28_11 + p_30_29;
  assign out_29_28 = t_r29_c28_12 >> 4;

  assign t_r29_c29_0 = p_28_29 << 1;
  assign t_r29_c29_1 = p_29_28 << 1;
  assign t_r29_c29_2 = p_29_29 << 2;
  assign t_r29_c29_3 = p_29_30 << 1;
  assign t_r29_c29_4 = p_30_29 << 1;
  assign t_r29_c29_5 = t_r29_c29_0 + p_28_28;
  assign t_r29_c29_6 = t_r29_c29_1 + p_28_30;
  assign t_r29_c29_7 = t_r29_c29_2 + t_r29_c29_3;
  assign t_r29_c29_8 = t_r29_c29_4 + p_30_28;
  assign t_r29_c29_9 = t_r29_c29_5 + t_r29_c29_6;
  assign t_r29_c29_10 = t_r29_c29_7 + t_r29_c29_8;
  assign t_r29_c29_11 = t_r29_c29_9 + t_r29_c29_10;
  assign t_r29_c29_12 = t_r29_c29_11 + p_30_30;
  assign out_29_29 = t_r29_c29_12 >> 4;

  assign t_r29_c30_0 = p_28_30 << 1;
  assign t_r29_c30_1 = p_29_29 << 1;
  assign t_r29_c30_2 = p_29_30 << 2;
  assign t_r29_c30_3 = p_29_31 << 1;
  assign t_r29_c30_4 = p_30_30 << 1;
  assign t_r29_c30_5 = t_r29_c30_0 + p_28_29;
  assign t_r29_c30_6 = t_r29_c30_1 + p_28_31;
  assign t_r29_c30_7 = t_r29_c30_2 + t_r29_c30_3;
  assign t_r29_c30_8 = t_r29_c30_4 + p_30_29;
  assign t_r29_c30_9 = t_r29_c30_5 + t_r29_c30_6;
  assign t_r29_c30_10 = t_r29_c30_7 + t_r29_c30_8;
  assign t_r29_c30_11 = t_r29_c30_9 + t_r29_c30_10;
  assign t_r29_c30_12 = t_r29_c30_11 + p_30_31;
  assign out_29_30 = t_r29_c30_12 >> 4;

  assign t_r29_c31_0 = p_28_31 << 1;
  assign t_r29_c31_1 = p_29_30 << 1;
  assign t_r29_c31_2 = p_29_31 << 2;
  assign t_r29_c31_3 = p_29_32 << 1;
  assign t_r29_c31_4 = p_30_31 << 1;
  assign t_r29_c31_5 = t_r29_c31_0 + p_28_30;
  assign t_r29_c31_6 = t_r29_c31_1 + p_28_32;
  assign t_r29_c31_7 = t_r29_c31_2 + t_r29_c31_3;
  assign t_r29_c31_8 = t_r29_c31_4 + p_30_30;
  assign t_r29_c31_9 = t_r29_c31_5 + t_r29_c31_6;
  assign t_r29_c31_10 = t_r29_c31_7 + t_r29_c31_8;
  assign t_r29_c31_11 = t_r29_c31_9 + t_r29_c31_10;
  assign t_r29_c31_12 = t_r29_c31_11 + p_30_32;
  assign out_29_31 = t_r29_c31_12 >> 4;

  assign t_r29_c32_0 = p_28_32 << 1;
  assign t_r29_c32_1 = p_29_31 << 1;
  assign t_r29_c32_2 = p_29_32 << 2;
  assign t_r29_c32_3 = p_29_33 << 1;
  assign t_r29_c32_4 = p_30_32 << 1;
  assign t_r29_c32_5 = t_r29_c32_0 + p_28_31;
  assign t_r29_c32_6 = t_r29_c32_1 + p_28_33;
  assign t_r29_c32_7 = t_r29_c32_2 + t_r29_c32_3;
  assign t_r29_c32_8 = t_r29_c32_4 + p_30_31;
  assign t_r29_c32_9 = t_r29_c32_5 + t_r29_c32_6;
  assign t_r29_c32_10 = t_r29_c32_7 + t_r29_c32_8;
  assign t_r29_c32_11 = t_r29_c32_9 + t_r29_c32_10;
  assign t_r29_c32_12 = t_r29_c32_11 + p_30_33;
  assign out_29_32 = t_r29_c32_12 >> 4;

  assign t_r29_c33_0 = p_28_33 << 1;
  assign t_r29_c33_1 = p_29_32 << 1;
  assign t_r29_c33_2 = p_29_33 << 2;
  assign t_r29_c33_3 = p_29_34 << 1;
  assign t_r29_c33_4 = p_30_33 << 1;
  assign t_r29_c33_5 = t_r29_c33_0 + p_28_32;
  assign t_r29_c33_6 = t_r29_c33_1 + p_28_34;
  assign t_r29_c33_7 = t_r29_c33_2 + t_r29_c33_3;
  assign t_r29_c33_8 = t_r29_c33_4 + p_30_32;
  assign t_r29_c33_9 = t_r29_c33_5 + t_r29_c33_6;
  assign t_r29_c33_10 = t_r29_c33_7 + t_r29_c33_8;
  assign t_r29_c33_11 = t_r29_c33_9 + t_r29_c33_10;
  assign t_r29_c33_12 = t_r29_c33_11 + p_30_34;
  assign out_29_33 = t_r29_c33_12 >> 4;

  assign t_r29_c34_0 = p_28_34 << 1;
  assign t_r29_c34_1 = p_29_33 << 1;
  assign t_r29_c34_2 = p_29_34 << 2;
  assign t_r29_c34_3 = p_29_35 << 1;
  assign t_r29_c34_4 = p_30_34 << 1;
  assign t_r29_c34_5 = t_r29_c34_0 + p_28_33;
  assign t_r29_c34_6 = t_r29_c34_1 + p_28_35;
  assign t_r29_c34_7 = t_r29_c34_2 + t_r29_c34_3;
  assign t_r29_c34_8 = t_r29_c34_4 + p_30_33;
  assign t_r29_c34_9 = t_r29_c34_5 + t_r29_c34_6;
  assign t_r29_c34_10 = t_r29_c34_7 + t_r29_c34_8;
  assign t_r29_c34_11 = t_r29_c34_9 + t_r29_c34_10;
  assign t_r29_c34_12 = t_r29_c34_11 + p_30_35;
  assign out_29_34 = t_r29_c34_12 >> 4;

  assign t_r29_c35_0 = p_28_35 << 1;
  assign t_r29_c35_1 = p_29_34 << 1;
  assign t_r29_c35_2 = p_29_35 << 2;
  assign t_r29_c35_3 = p_29_36 << 1;
  assign t_r29_c35_4 = p_30_35 << 1;
  assign t_r29_c35_5 = t_r29_c35_0 + p_28_34;
  assign t_r29_c35_6 = t_r29_c35_1 + p_28_36;
  assign t_r29_c35_7 = t_r29_c35_2 + t_r29_c35_3;
  assign t_r29_c35_8 = t_r29_c35_4 + p_30_34;
  assign t_r29_c35_9 = t_r29_c35_5 + t_r29_c35_6;
  assign t_r29_c35_10 = t_r29_c35_7 + t_r29_c35_8;
  assign t_r29_c35_11 = t_r29_c35_9 + t_r29_c35_10;
  assign t_r29_c35_12 = t_r29_c35_11 + p_30_36;
  assign out_29_35 = t_r29_c35_12 >> 4;

  assign t_r29_c36_0 = p_28_36 << 1;
  assign t_r29_c36_1 = p_29_35 << 1;
  assign t_r29_c36_2 = p_29_36 << 2;
  assign t_r29_c36_3 = p_29_37 << 1;
  assign t_r29_c36_4 = p_30_36 << 1;
  assign t_r29_c36_5 = t_r29_c36_0 + p_28_35;
  assign t_r29_c36_6 = t_r29_c36_1 + p_28_37;
  assign t_r29_c36_7 = t_r29_c36_2 + t_r29_c36_3;
  assign t_r29_c36_8 = t_r29_c36_4 + p_30_35;
  assign t_r29_c36_9 = t_r29_c36_5 + t_r29_c36_6;
  assign t_r29_c36_10 = t_r29_c36_7 + t_r29_c36_8;
  assign t_r29_c36_11 = t_r29_c36_9 + t_r29_c36_10;
  assign t_r29_c36_12 = t_r29_c36_11 + p_30_37;
  assign out_29_36 = t_r29_c36_12 >> 4;

  assign t_r29_c37_0 = p_28_37 << 1;
  assign t_r29_c37_1 = p_29_36 << 1;
  assign t_r29_c37_2 = p_29_37 << 2;
  assign t_r29_c37_3 = p_29_38 << 1;
  assign t_r29_c37_4 = p_30_37 << 1;
  assign t_r29_c37_5 = t_r29_c37_0 + p_28_36;
  assign t_r29_c37_6 = t_r29_c37_1 + p_28_38;
  assign t_r29_c37_7 = t_r29_c37_2 + t_r29_c37_3;
  assign t_r29_c37_8 = t_r29_c37_4 + p_30_36;
  assign t_r29_c37_9 = t_r29_c37_5 + t_r29_c37_6;
  assign t_r29_c37_10 = t_r29_c37_7 + t_r29_c37_8;
  assign t_r29_c37_11 = t_r29_c37_9 + t_r29_c37_10;
  assign t_r29_c37_12 = t_r29_c37_11 + p_30_38;
  assign out_29_37 = t_r29_c37_12 >> 4;

  assign t_r29_c38_0 = p_28_38 << 1;
  assign t_r29_c38_1 = p_29_37 << 1;
  assign t_r29_c38_2 = p_29_38 << 2;
  assign t_r29_c38_3 = p_29_39 << 1;
  assign t_r29_c38_4 = p_30_38 << 1;
  assign t_r29_c38_5 = t_r29_c38_0 + p_28_37;
  assign t_r29_c38_6 = t_r29_c38_1 + p_28_39;
  assign t_r29_c38_7 = t_r29_c38_2 + t_r29_c38_3;
  assign t_r29_c38_8 = t_r29_c38_4 + p_30_37;
  assign t_r29_c38_9 = t_r29_c38_5 + t_r29_c38_6;
  assign t_r29_c38_10 = t_r29_c38_7 + t_r29_c38_8;
  assign t_r29_c38_11 = t_r29_c38_9 + t_r29_c38_10;
  assign t_r29_c38_12 = t_r29_c38_11 + p_30_39;
  assign out_29_38 = t_r29_c38_12 >> 4;

  assign t_r29_c39_0 = p_28_39 << 1;
  assign t_r29_c39_1 = p_29_38 << 1;
  assign t_r29_c39_2 = p_29_39 << 2;
  assign t_r29_c39_3 = p_29_40 << 1;
  assign t_r29_c39_4 = p_30_39 << 1;
  assign t_r29_c39_5 = t_r29_c39_0 + p_28_38;
  assign t_r29_c39_6 = t_r29_c39_1 + p_28_40;
  assign t_r29_c39_7 = t_r29_c39_2 + t_r29_c39_3;
  assign t_r29_c39_8 = t_r29_c39_4 + p_30_38;
  assign t_r29_c39_9 = t_r29_c39_5 + t_r29_c39_6;
  assign t_r29_c39_10 = t_r29_c39_7 + t_r29_c39_8;
  assign t_r29_c39_11 = t_r29_c39_9 + t_r29_c39_10;
  assign t_r29_c39_12 = t_r29_c39_11 + p_30_40;
  assign out_29_39 = t_r29_c39_12 >> 4;

  assign t_r29_c40_0 = p_28_40 << 1;
  assign t_r29_c40_1 = p_29_39 << 1;
  assign t_r29_c40_2 = p_29_40 << 2;
  assign t_r29_c40_3 = p_29_41 << 1;
  assign t_r29_c40_4 = p_30_40 << 1;
  assign t_r29_c40_5 = t_r29_c40_0 + p_28_39;
  assign t_r29_c40_6 = t_r29_c40_1 + p_28_41;
  assign t_r29_c40_7 = t_r29_c40_2 + t_r29_c40_3;
  assign t_r29_c40_8 = t_r29_c40_4 + p_30_39;
  assign t_r29_c40_9 = t_r29_c40_5 + t_r29_c40_6;
  assign t_r29_c40_10 = t_r29_c40_7 + t_r29_c40_8;
  assign t_r29_c40_11 = t_r29_c40_9 + t_r29_c40_10;
  assign t_r29_c40_12 = t_r29_c40_11 + p_30_41;
  assign out_29_40 = t_r29_c40_12 >> 4;

  assign t_r29_c41_0 = p_28_41 << 1;
  assign t_r29_c41_1 = p_29_40 << 1;
  assign t_r29_c41_2 = p_29_41 << 2;
  assign t_r29_c41_3 = p_29_42 << 1;
  assign t_r29_c41_4 = p_30_41 << 1;
  assign t_r29_c41_5 = t_r29_c41_0 + p_28_40;
  assign t_r29_c41_6 = t_r29_c41_1 + p_28_42;
  assign t_r29_c41_7 = t_r29_c41_2 + t_r29_c41_3;
  assign t_r29_c41_8 = t_r29_c41_4 + p_30_40;
  assign t_r29_c41_9 = t_r29_c41_5 + t_r29_c41_6;
  assign t_r29_c41_10 = t_r29_c41_7 + t_r29_c41_8;
  assign t_r29_c41_11 = t_r29_c41_9 + t_r29_c41_10;
  assign t_r29_c41_12 = t_r29_c41_11 + p_30_42;
  assign out_29_41 = t_r29_c41_12 >> 4;

  assign t_r29_c42_0 = p_28_42 << 1;
  assign t_r29_c42_1 = p_29_41 << 1;
  assign t_r29_c42_2 = p_29_42 << 2;
  assign t_r29_c42_3 = p_29_43 << 1;
  assign t_r29_c42_4 = p_30_42 << 1;
  assign t_r29_c42_5 = t_r29_c42_0 + p_28_41;
  assign t_r29_c42_6 = t_r29_c42_1 + p_28_43;
  assign t_r29_c42_7 = t_r29_c42_2 + t_r29_c42_3;
  assign t_r29_c42_8 = t_r29_c42_4 + p_30_41;
  assign t_r29_c42_9 = t_r29_c42_5 + t_r29_c42_6;
  assign t_r29_c42_10 = t_r29_c42_7 + t_r29_c42_8;
  assign t_r29_c42_11 = t_r29_c42_9 + t_r29_c42_10;
  assign t_r29_c42_12 = t_r29_c42_11 + p_30_43;
  assign out_29_42 = t_r29_c42_12 >> 4;

  assign t_r29_c43_0 = p_28_43 << 1;
  assign t_r29_c43_1 = p_29_42 << 1;
  assign t_r29_c43_2 = p_29_43 << 2;
  assign t_r29_c43_3 = p_29_44 << 1;
  assign t_r29_c43_4 = p_30_43 << 1;
  assign t_r29_c43_5 = t_r29_c43_0 + p_28_42;
  assign t_r29_c43_6 = t_r29_c43_1 + p_28_44;
  assign t_r29_c43_7 = t_r29_c43_2 + t_r29_c43_3;
  assign t_r29_c43_8 = t_r29_c43_4 + p_30_42;
  assign t_r29_c43_9 = t_r29_c43_5 + t_r29_c43_6;
  assign t_r29_c43_10 = t_r29_c43_7 + t_r29_c43_8;
  assign t_r29_c43_11 = t_r29_c43_9 + t_r29_c43_10;
  assign t_r29_c43_12 = t_r29_c43_11 + p_30_44;
  assign out_29_43 = t_r29_c43_12 >> 4;

  assign t_r29_c44_0 = p_28_44 << 1;
  assign t_r29_c44_1 = p_29_43 << 1;
  assign t_r29_c44_2 = p_29_44 << 2;
  assign t_r29_c44_3 = p_29_45 << 1;
  assign t_r29_c44_4 = p_30_44 << 1;
  assign t_r29_c44_5 = t_r29_c44_0 + p_28_43;
  assign t_r29_c44_6 = t_r29_c44_1 + p_28_45;
  assign t_r29_c44_7 = t_r29_c44_2 + t_r29_c44_3;
  assign t_r29_c44_8 = t_r29_c44_4 + p_30_43;
  assign t_r29_c44_9 = t_r29_c44_5 + t_r29_c44_6;
  assign t_r29_c44_10 = t_r29_c44_7 + t_r29_c44_8;
  assign t_r29_c44_11 = t_r29_c44_9 + t_r29_c44_10;
  assign t_r29_c44_12 = t_r29_c44_11 + p_30_45;
  assign out_29_44 = t_r29_c44_12 >> 4;

  assign t_r29_c45_0 = p_28_45 << 1;
  assign t_r29_c45_1 = p_29_44 << 1;
  assign t_r29_c45_2 = p_29_45 << 2;
  assign t_r29_c45_3 = p_29_46 << 1;
  assign t_r29_c45_4 = p_30_45 << 1;
  assign t_r29_c45_5 = t_r29_c45_0 + p_28_44;
  assign t_r29_c45_6 = t_r29_c45_1 + p_28_46;
  assign t_r29_c45_7 = t_r29_c45_2 + t_r29_c45_3;
  assign t_r29_c45_8 = t_r29_c45_4 + p_30_44;
  assign t_r29_c45_9 = t_r29_c45_5 + t_r29_c45_6;
  assign t_r29_c45_10 = t_r29_c45_7 + t_r29_c45_8;
  assign t_r29_c45_11 = t_r29_c45_9 + t_r29_c45_10;
  assign t_r29_c45_12 = t_r29_c45_11 + p_30_46;
  assign out_29_45 = t_r29_c45_12 >> 4;

  assign t_r29_c46_0 = p_28_46 << 1;
  assign t_r29_c46_1 = p_29_45 << 1;
  assign t_r29_c46_2 = p_29_46 << 2;
  assign t_r29_c46_3 = p_29_47 << 1;
  assign t_r29_c46_4 = p_30_46 << 1;
  assign t_r29_c46_5 = t_r29_c46_0 + p_28_45;
  assign t_r29_c46_6 = t_r29_c46_1 + p_28_47;
  assign t_r29_c46_7 = t_r29_c46_2 + t_r29_c46_3;
  assign t_r29_c46_8 = t_r29_c46_4 + p_30_45;
  assign t_r29_c46_9 = t_r29_c46_5 + t_r29_c46_6;
  assign t_r29_c46_10 = t_r29_c46_7 + t_r29_c46_8;
  assign t_r29_c46_11 = t_r29_c46_9 + t_r29_c46_10;
  assign t_r29_c46_12 = t_r29_c46_11 + p_30_47;
  assign out_29_46 = t_r29_c46_12 >> 4;

  assign t_r29_c47_0 = p_28_47 << 1;
  assign t_r29_c47_1 = p_29_46 << 1;
  assign t_r29_c47_2 = p_29_47 << 2;
  assign t_r29_c47_3 = p_29_48 << 1;
  assign t_r29_c47_4 = p_30_47 << 1;
  assign t_r29_c47_5 = t_r29_c47_0 + p_28_46;
  assign t_r29_c47_6 = t_r29_c47_1 + p_28_48;
  assign t_r29_c47_7 = t_r29_c47_2 + t_r29_c47_3;
  assign t_r29_c47_8 = t_r29_c47_4 + p_30_46;
  assign t_r29_c47_9 = t_r29_c47_5 + t_r29_c47_6;
  assign t_r29_c47_10 = t_r29_c47_7 + t_r29_c47_8;
  assign t_r29_c47_11 = t_r29_c47_9 + t_r29_c47_10;
  assign t_r29_c47_12 = t_r29_c47_11 + p_30_48;
  assign out_29_47 = t_r29_c47_12 >> 4;

  assign t_r29_c48_0 = p_28_48 << 1;
  assign t_r29_c48_1 = p_29_47 << 1;
  assign t_r29_c48_2 = p_29_48 << 2;
  assign t_r29_c48_3 = p_29_49 << 1;
  assign t_r29_c48_4 = p_30_48 << 1;
  assign t_r29_c48_5 = t_r29_c48_0 + p_28_47;
  assign t_r29_c48_6 = t_r29_c48_1 + p_28_49;
  assign t_r29_c48_7 = t_r29_c48_2 + t_r29_c48_3;
  assign t_r29_c48_8 = t_r29_c48_4 + p_30_47;
  assign t_r29_c48_9 = t_r29_c48_5 + t_r29_c48_6;
  assign t_r29_c48_10 = t_r29_c48_7 + t_r29_c48_8;
  assign t_r29_c48_11 = t_r29_c48_9 + t_r29_c48_10;
  assign t_r29_c48_12 = t_r29_c48_11 + p_30_49;
  assign out_29_48 = t_r29_c48_12 >> 4;

  assign t_r29_c49_0 = p_28_49 << 1;
  assign t_r29_c49_1 = p_29_48 << 1;
  assign t_r29_c49_2 = p_29_49 << 2;
  assign t_r29_c49_3 = p_29_50 << 1;
  assign t_r29_c49_4 = p_30_49 << 1;
  assign t_r29_c49_5 = t_r29_c49_0 + p_28_48;
  assign t_r29_c49_6 = t_r29_c49_1 + p_28_50;
  assign t_r29_c49_7 = t_r29_c49_2 + t_r29_c49_3;
  assign t_r29_c49_8 = t_r29_c49_4 + p_30_48;
  assign t_r29_c49_9 = t_r29_c49_5 + t_r29_c49_6;
  assign t_r29_c49_10 = t_r29_c49_7 + t_r29_c49_8;
  assign t_r29_c49_11 = t_r29_c49_9 + t_r29_c49_10;
  assign t_r29_c49_12 = t_r29_c49_11 + p_30_50;
  assign out_29_49 = t_r29_c49_12 >> 4;

  assign t_r29_c50_0 = p_28_50 << 1;
  assign t_r29_c50_1 = p_29_49 << 1;
  assign t_r29_c50_2 = p_29_50 << 2;
  assign t_r29_c50_3 = p_29_51 << 1;
  assign t_r29_c50_4 = p_30_50 << 1;
  assign t_r29_c50_5 = t_r29_c50_0 + p_28_49;
  assign t_r29_c50_6 = t_r29_c50_1 + p_28_51;
  assign t_r29_c50_7 = t_r29_c50_2 + t_r29_c50_3;
  assign t_r29_c50_8 = t_r29_c50_4 + p_30_49;
  assign t_r29_c50_9 = t_r29_c50_5 + t_r29_c50_6;
  assign t_r29_c50_10 = t_r29_c50_7 + t_r29_c50_8;
  assign t_r29_c50_11 = t_r29_c50_9 + t_r29_c50_10;
  assign t_r29_c50_12 = t_r29_c50_11 + p_30_51;
  assign out_29_50 = t_r29_c50_12 >> 4;

  assign t_r29_c51_0 = p_28_51 << 1;
  assign t_r29_c51_1 = p_29_50 << 1;
  assign t_r29_c51_2 = p_29_51 << 2;
  assign t_r29_c51_3 = p_29_52 << 1;
  assign t_r29_c51_4 = p_30_51 << 1;
  assign t_r29_c51_5 = t_r29_c51_0 + p_28_50;
  assign t_r29_c51_6 = t_r29_c51_1 + p_28_52;
  assign t_r29_c51_7 = t_r29_c51_2 + t_r29_c51_3;
  assign t_r29_c51_8 = t_r29_c51_4 + p_30_50;
  assign t_r29_c51_9 = t_r29_c51_5 + t_r29_c51_6;
  assign t_r29_c51_10 = t_r29_c51_7 + t_r29_c51_8;
  assign t_r29_c51_11 = t_r29_c51_9 + t_r29_c51_10;
  assign t_r29_c51_12 = t_r29_c51_11 + p_30_52;
  assign out_29_51 = t_r29_c51_12 >> 4;

  assign t_r29_c52_0 = p_28_52 << 1;
  assign t_r29_c52_1 = p_29_51 << 1;
  assign t_r29_c52_2 = p_29_52 << 2;
  assign t_r29_c52_3 = p_29_53 << 1;
  assign t_r29_c52_4 = p_30_52 << 1;
  assign t_r29_c52_5 = t_r29_c52_0 + p_28_51;
  assign t_r29_c52_6 = t_r29_c52_1 + p_28_53;
  assign t_r29_c52_7 = t_r29_c52_2 + t_r29_c52_3;
  assign t_r29_c52_8 = t_r29_c52_4 + p_30_51;
  assign t_r29_c52_9 = t_r29_c52_5 + t_r29_c52_6;
  assign t_r29_c52_10 = t_r29_c52_7 + t_r29_c52_8;
  assign t_r29_c52_11 = t_r29_c52_9 + t_r29_c52_10;
  assign t_r29_c52_12 = t_r29_c52_11 + p_30_53;
  assign out_29_52 = t_r29_c52_12 >> 4;

  assign t_r29_c53_0 = p_28_53 << 1;
  assign t_r29_c53_1 = p_29_52 << 1;
  assign t_r29_c53_2 = p_29_53 << 2;
  assign t_r29_c53_3 = p_29_54 << 1;
  assign t_r29_c53_4 = p_30_53 << 1;
  assign t_r29_c53_5 = t_r29_c53_0 + p_28_52;
  assign t_r29_c53_6 = t_r29_c53_1 + p_28_54;
  assign t_r29_c53_7 = t_r29_c53_2 + t_r29_c53_3;
  assign t_r29_c53_8 = t_r29_c53_4 + p_30_52;
  assign t_r29_c53_9 = t_r29_c53_5 + t_r29_c53_6;
  assign t_r29_c53_10 = t_r29_c53_7 + t_r29_c53_8;
  assign t_r29_c53_11 = t_r29_c53_9 + t_r29_c53_10;
  assign t_r29_c53_12 = t_r29_c53_11 + p_30_54;
  assign out_29_53 = t_r29_c53_12 >> 4;

  assign t_r29_c54_0 = p_28_54 << 1;
  assign t_r29_c54_1 = p_29_53 << 1;
  assign t_r29_c54_2 = p_29_54 << 2;
  assign t_r29_c54_3 = p_29_55 << 1;
  assign t_r29_c54_4 = p_30_54 << 1;
  assign t_r29_c54_5 = t_r29_c54_0 + p_28_53;
  assign t_r29_c54_6 = t_r29_c54_1 + p_28_55;
  assign t_r29_c54_7 = t_r29_c54_2 + t_r29_c54_3;
  assign t_r29_c54_8 = t_r29_c54_4 + p_30_53;
  assign t_r29_c54_9 = t_r29_c54_5 + t_r29_c54_6;
  assign t_r29_c54_10 = t_r29_c54_7 + t_r29_c54_8;
  assign t_r29_c54_11 = t_r29_c54_9 + t_r29_c54_10;
  assign t_r29_c54_12 = t_r29_c54_11 + p_30_55;
  assign out_29_54 = t_r29_c54_12 >> 4;

  assign t_r29_c55_0 = p_28_55 << 1;
  assign t_r29_c55_1 = p_29_54 << 1;
  assign t_r29_c55_2 = p_29_55 << 2;
  assign t_r29_c55_3 = p_29_56 << 1;
  assign t_r29_c55_4 = p_30_55 << 1;
  assign t_r29_c55_5 = t_r29_c55_0 + p_28_54;
  assign t_r29_c55_6 = t_r29_c55_1 + p_28_56;
  assign t_r29_c55_7 = t_r29_c55_2 + t_r29_c55_3;
  assign t_r29_c55_8 = t_r29_c55_4 + p_30_54;
  assign t_r29_c55_9 = t_r29_c55_5 + t_r29_c55_6;
  assign t_r29_c55_10 = t_r29_c55_7 + t_r29_c55_8;
  assign t_r29_c55_11 = t_r29_c55_9 + t_r29_c55_10;
  assign t_r29_c55_12 = t_r29_c55_11 + p_30_56;
  assign out_29_55 = t_r29_c55_12 >> 4;

  assign t_r29_c56_0 = p_28_56 << 1;
  assign t_r29_c56_1 = p_29_55 << 1;
  assign t_r29_c56_2 = p_29_56 << 2;
  assign t_r29_c56_3 = p_29_57 << 1;
  assign t_r29_c56_4 = p_30_56 << 1;
  assign t_r29_c56_5 = t_r29_c56_0 + p_28_55;
  assign t_r29_c56_6 = t_r29_c56_1 + p_28_57;
  assign t_r29_c56_7 = t_r29_c56_2 + t_r29_c56_3;
  assign t_r29_c56_8 = t_r29_c56_4 + p_30_55;
  assign t_r29_c56_9 = t_r29_c56_5 + t_r29_c56_6;
  assign t_r29_c56_10 = t_r29_c56_7 + t_r29_c56_8;
  assign t_r29_c56_11 = t_r29_c56_9 + t_r29_c56_10;
  assign t_r29_c56_12 = t_r29_c56_11 + p_30_57;
  assign out_29_56 = t_r29_c56_12 >> 4;

  assign t_r29_c57_0 = p_28_57 << 1;
  assign t_r29_c57_1 = p_29_56 << 1;
  assign t_r29_c57_2 = p_29_57 << 2;
  assign t_r29_c57_3 = p_29_58 << 1;
  assign t_r29_c57_4 = p_30_57 << 1;
  assign t_r29_c57_5 = t_r29_c57_0 + p_28_56;
  assign t_r29_c57_6 = t_r29_c57_1 + p_28_58;
  assign t_r29_c57_7 = t_r29_c57_2 + t_r29_c57_3;
  assign t_r29_c57_8 = t_r29_c57_4 + p_30_56;
  assign t_r29_c57_9 = t_r29_c57_5 + t_r29_c57_6;
  assign t_r29_c57_10 = t_r29_c57_7 + t_r29_c57_8;
  assign t_r29_c57_11 = t_r29_c57_9 + t_r29_c57_10;
  assign t_r29_c57_12 = t_r29_c57_11 + p_30_58;
  assign out_29_57 = t_r29_c57_12 >> 4;

  assign t_r29_c58_0 = p_28_58 << 1;
  assign t_r29_c58_1 = p_29_57 << 1;
  assign t_r29_c58_2 = p_29_58 << 2;
  assign t_r29_c58_3 = p_29_59 << 1;
  assign t_r29_c58_4 = p_30_58 << 1;
  assign t_r29_c58_5 = t_r29_c58_0 + p_28_57;
  assign t_r29_c58_6 = t_r29_c58_1 + p_28_59;
  assign t_r29_c58_7 = t_r29_c58_2 + t_r29_c58_3;
  assign t_r29_c58_8 = t_r29_c58_4 + p_30_57;
  assign t_r29_c58_9 = t_r29_c58_5 + t_r29_c58_6;
  assign t_r29_c58_10 = t_r29_c58_7 + t_r29_c58_8;
  assign t_r29_c58_11 = t_r29_c58_9 + t_r29_c58_10;
  assign t_r29_c58_12 = t_r29_c58_11 + p_30_59;
  assign out_29_58 = t_r29_c58_12 >> 4;

  assign t_r29_c59_0 = p_28_59 << 1;
  assign t_r29_c59_1 = p_29_58 << 1;
  assign t_r29_c59_2 = p_29_59 << 2;
  assign t_r29_c59_3 = p_29_60 << 1;
  assign t_r29_c59_4 = p_30_59 << 1;
  assign t_r29_c59_5 = t_r29_c59_0 + p_28_58;
  assign t_r29_c59_6 = t_r29_c59_1 + p_28_60;
  assign t_r29_c59_7 = t_r29_c59_2 + t_r29_c59_3;
  assign t_r29_c59_8 = t_r29_c59_4 + p_30_58;
  assign t_r29_c59_9 = t_r29_c59_5 + t_r29_c59_6;
  assign t_r29_c59_10 = t_r29_c59_7 + t_r29_c59_8;
  assign t_r29_c59_11 = t_r29_c59_9 + t_r29_c59_10;
  assign t_r29_c59_12 = t_r29_c59_11 + p_30_60;
  assign out_29_59 = t_r29_c59_12 >> 4;

  assign t_r29_c60_0 = p_28_60 << 1;
  assign t_r29_c60_1 = p_29_59 << 1;
  assign t_r29_c60_2 = p_29_60 << 2;
  assign t_r29_c60_3 = p_29_61 << 1;
  assign t_r29_c60_4 = p_30_60 << 1;
  assign t_r29_c60_5 = t_r29_c60_0 + p_28_59;
  assign t_r29_c60_6 = t_r29_c60_1 + p_28_61;
  assign t_r29_c60_7 = t_r29_c60_2 + t_r29_c60_3;
  assign t_r29_c60_8 = t_r29_c60_4 + p_30_59;
  assign t_r29_c60_9 = t_r29_c60_5 + t_r29_c60_6;
  assign t_r29_c60_10 = t_r29_c60_7 + t_r29_c60_8;
  assign t_r29_c60_11 = t_r29_c60_9 + t_r29_c60_10;
  assign t_r29_c60_12 = t_r29_c60_11 + p_30_61;
  assign out_29_60 = t_r29_c60_12 >> 4;

  assign t_r29_c61_0 = p_28_61 << 1;
  assign t_r29_c61_1 = p_29_60 << 1;
  assign t_r29_c61_2 = p_29_61 << 2;
  assign t_r29_c61_3 = p_29_62 << 1;
  assign t_r29_c61_4 = p_30_61 << 1;
  assign t_r29_c61_5 = t_r29_c61_0 + p_28_60;
  assign t_r29_c61_6 = t_r29_c61_1 + p_28_62;
  assign t_r29_c61_7 = t_r29_c61_2 + t_r29_c61_3;
  assign t_r29_c61_8 = t_r29_c61_4 + p_30_60;
  assign t_r29_c61_9 = t_r29_c61_5 + t_r29_c61_6;
  assign t_r29_c61_10 = t_r29_c61_7 + t_r29_c61_8;
  assign t_r29_c61_11 = t_r29_c61_9 + t_r29_c61_10;
  assign t_r29_c61_12 = t_r29_c61_11 + p_30_62;
  assign out_29_61 = t_r29_c61_12 >> 4;

  assign t_r29_c62_0 = p_28_62 << 1;
  assign t_r29_c62_1 = p_29_61 << 1;
  assign t_r29_c62_2 = p_29_62 << 2;
  assign t_r29_c62_3 = p_29_63 << 1;
  assign t_r29_c62_4 = p_30_62 << 1;
  assign t_r29_c62_5 = t_r29_c62_0 + p_28_61;
  assign t_r29_c62_6 = t_r29_c62_1 + p_28_63;
  assign t_r29_c62_7 = t_r29_c62_2 + t_r29_c62_3;
  assign t_r29_c62_8 = t_r29_c62_4 + p_30_61;
  assign t_r29_c62_9 = t_r29_c62_5 + t_r29_c62_6;
  assign t_r29_c62_10 = t_r29_c62_7 + t_r29_c62_8;
  assign t_r29_c62_11 = t_r29_c62_9 + t_r29_c62_10;
  assign t_r29_c62_12 = t_r29_c62_11 + p_30_63;
  assign out_29_62 = t_r29_c62_12 >> 4;

  assign t_r29_c63_0 = p_28_63 << 1;
  assign t_r29_c63_1 = p_29_62 << 1;
  assign t_r29_c63_2 = p_29_63 << 2;
  assign t_r29_c63_3 = p_29_64 << 1;
  assign t_r29_c63_4 = p_30_63 << 1;
  assign t_r29_c63_5 = t_r29_c63_0 + p_28_62;
  assign t_r29_c63_6 = t_r29_c63_1 + p_28_64;
  assign t_r29_c63_7 = t_r29_c63_2 + t_r29_c63_3;
  assign t_r29_c63_8 = t_r29_c63_4 + p_30_62;
  assign t_r29_c63_9 = t_r29_c63_5 + t_r29_c63_6;
  assign t_r29_c63_10 = t_r29_c63_7 + t_r29_c63_8;
  assign t_r29_c63_11 = t_r29_c63_9 + t_r29_c63_10;
  assign t_r29_c63_12 = t_r29_c63_11 + p_30_64;
  assign out_29_63 = t_r29_c63_12 >> 4;

  assign t_r29_c64_0 = p_28_64 << 1;
  assign t_r29_c64_1 = p_29_63 << 1;
  assign t_r29_c64_2 = p_29_64 << 2;
  assign t_r29_c64_3 = p_29_65 << 1;
  assign t_r29_c64_4 = p_30_64 << 1;
  assign t_r29_c64_5 = t_r29_c64_0 + p_28_63;
  assign t_r29_c64_6 = t_r29_c64_1 + p_28_65;
  assign t_r29_c64_7 = t_r29_c64_2 + t_r29_c64_3;
  assign t_r29_c64_8 = t_r29_c64_4 + p_30_63;
  assign t_r29_c64_9 = t_r29_c64_5 + t_r29_c64_6;
  assign t_r29_c64_10 = t_r29_c64_7 + t_r29_c64_8;
  assign t_r29_c64_11 = t_r29_c64_9 + t_r29_c64_10;
  assign t_r29_c64_12 = t_r29_c64_11 + p_30_65;
  assign out_29_64 = t_r29_c64_12 >> 4;

  assign t_r30_c1_0 = p_29_1 << 1;
  assign t_r30_c1_1 = p_30_0 << 1;
  assign t_r30_c1_2 = p_30_1 << 2;
  assign t_r30_c1_3 = p_30_2 << 1;
  assign t_r30_c1_4 = p_31_1 << 1;
  assign t_r30_c1_5 = t_r30_c1_0 + p_29_0;
  assign t_r30_c1_6 = t_r30_c1_1 + p_29_2;
  assign t_r30_c1_7 = t_r30_c1_2 + t_r30_c1_3;
  assign t_r30_c1_8 = t_r30_c1_4 + p_31_0;
  assign t_r30_c1_9 = t_r30_c1_5 + t_r30_c1_6;
  assign t_r30_c1_10 = t_r30_c1_7 + t_r30_c1_8;
  assign t_r30_c1_11 = t_r30_c1_9 + t_r30_c1_10;
  assign t_r30_c1_12 = t_r30_c1_11 + p_31_2;
  assign out_30_1 = t_r30_c1_12 >> 4;

  assign t_r30_c2_0 = p_29_2 << 1;
  assign t_r30_c2_1 = p_30_1 << 1;
  assign t_r30_c2_2 = p_30_2 << 2;
  assign t_r30_c2_3 = p_30_3 << 1;
  assign t_r30_c2_4 = p_31_2 << 1;
  assign t_r30_c2_5 = t_r30_c2_0 + p_29_1;
  assign t_r30_c2_6 = t_r30_c2_1 + p_29_3;
  assign t_r30_c2_7 = t_r30_c2_2 + t_r30_c2_3;
  assign t_r30_c2_8 = t_r30_c2_4 + p_31_1;
  assign t_r30_c2_9 = t_r30_c2_5 + t_r30_c2_6;
  assign t_r30_c2_10 = t_r30_c2_7 + t_r30_c2_8;
  assign t_r30_c2_11 = t_r30_c2_9 + t_r30_c2_10;
  assign t_r30_c2_12 = t_r30_c2_11 + p_31_3;
  assign out_30_2 = t_r30_c2_12 >> 4;

  assign t_r30_c3_0 = p_29_3 << 1;
  assign t_r30_c3_1 = p_30_2 << 1;
  assign t_r30_c3_2 = p_30_3 << 2;
  assign t_r30_c3_3 = p_30_4 << 1;
  assign t_r30_c3_4 = p_31_3 << 1;
  assign t_r30_c3_5 = t_r30_c3_0 + p_29_2;
  assign t_r30_c3_6 = t_r30_c3_1 + p_29_4;
  assign t_r30_c3_7 = t_r30_c3_2 + t_r30_c3_3;
  assign t_r30_c3_8 = t_r30_c3_4 + p_31_2;
  assign t_r30_c3_9 = t_r30_c3_5 + t_r30_c3_6;
  assign t_r30_c3_10 = t_r30_c3_7 + t_r30_c3_8;
  assign t_r30_c3_11 = t_r30_c3_9 + t_r30_c3_10;
  assign t_r30_c3_12 = t_r30_c3_11 + p_31_4;
  assign out_30_3 = t_r30_c3_12 >> 4;

  assign t_r30_c4_0 = p_29_4 << 1;
  assign t_r30_c4_1 = p_30_3 << 1;
  assign t_r30_c4_2 = p_30_4 << 2;
  assign t_r30_c4_3 = p_30_5 << 1;
  assign t_r30_c4_4 = p_31_4 << 1;
  assign t_r30_c4_5 = t_r30_c4_0 + p_29_3;
  assign t_r30_c4_6 = t_r30_c4_1 + p_29_5;
  assign t_r30_c4_7 = t_r30_c4_2 + t_r30_c4_3;
  assign t_r30_c4_8 = t_r30_c4_4 + p_31_3;
  assign t_r30_c4_9 = t_r30_c4_5 + t_r30_c4_6;
  assign t_r30_c4_10 = t_r30_c4_7 + t_r30_c4_8;
  assign t_r30_c4_11 = t_r30_c4_9 + t_r30_c4_10;
  assign t_r30_c4_12 = t_r30_c4_11 + p_31_5;
  assign out_30_4 = t_r30_c4_12 >> 4;

  assign t_r30_c5_0 = p_29_5 << 1;
  assign t_r30_c5_1 = p_30_4 << 1;
  assign t_r30_c5_2 = p_30_5 << 2;
  assign t_r30_c5_3 = p_30_6 << 1;
  assign t_r30_c5_4 = p_31_5 << 1;
  assign t_r30_c5_5 = t_r30_c5_0 + p_29_4;
  assign t_r30_c5_6 = t_r30_c5_1 + p_29_6;
  assign t_r30_c5_7 = t_r30_c5_2 + t_r30_c5_3;
  assign t_r30_c5_8 = t_r30_c5_4 + p_31_4;
  assign t_r30_c5_9 = t_r30_c5_5 + t_r30_c5_6;
  assign t_r30_c5_10 = t_r30_c5_7 + t_r30_c5_8;
  assign t_r30_c5_11 = t_r30_c5_9 + t_r30_c5_10;
  assign t_r30_c5_12 = t_r30_c5_11 + p_31_6;
  assign out_30_5 = t_r30_c5_12 >> 4;

  assign t_r30_c6_0 = p_29_6 << 1;
  assign t_r30_c6_1 = p_30_5 << 1;
  assign t_r30_c6_2 = p_30_6 << 2;
  assign t_r30_c6_3 = p_30_7 << 1;
  assign t_r30_c6_4 = p_31_6 << 1;
  assign t_r30_c6_5 = t_r30_c6_0 + p_29_5;
  assign t_r30_c6_6 = t_r30_c6_1 + p_29_7;
  assign t_r30_c6_7 = t_r30_c6_2 + t_r30_c6_3;
  assign t_r30_c6_8 = t_r30_c6_4 + p_31_5;
  assign t_r30_c6_9 = t_r30_c6_5 + t_r30_c6_6;
  assign t_r30_c6_10 = t_r30_c6_7 + t_r30_c6_8;
  assign t_r30_c6_11 = t_r30_c6_9 + t_r30_c6_10;
  assign t_r30_c6_12 = t_r30_c6_11 + p_31_7;
  assign out_30_6 = t_r30_c6_12 >> 4;

  assign t_r30_c7_0 = p_29_7 << 1;
  assign t_r30_c7_1 = p_30_6 << 1;
  assign t_r30_c7_2 = p_30_7 << 2;
  assign t_r30_c7_3 = p_30_8 << 1;
  assign t_r30_c7_4 = p_31_7 << 1;
  assign t_r30_c7_5 = t_r30_c7_0 + p_29_6;
  assign t_r30_c7_6 = t_r30_c7_1 + p_29_8;
  assign t_r30_c7_7 = t_r30_c7_2 + t_r30_c7_3;
  assign t_r30_c7_8 = t_r30_c7_4 + p_31_6;
  assign t_r30_c7_9 = t_r30_c7_5 + t_r30_c7_6;
  assign t_r30_c7_10 = t_r30_c7_7 + t_r30_c7_8;
  assign t_r30_c7_11 = t_r30_c7_9 + t_r30_c7_10;
  assign t_r30_c7_12 = t_r30_c7_11 + p_31_8;
  assign out_30_7 = t_r30_c7_12 >> 4;

  assign t_r30_c8_0 = p_29_8 << 1;
  assign t_r30_c8_1 = p_30_7 << 1;
  assign t_r30_c8_2 = p_30_8 << 2;
  assign t_r30_c8_3 = p_30_9 << 1;
  assign t_r30_c8_4 = p_31_8 << 1;
  assign t_r30_c8_5 = t_r30_c8_0 + p_29_7;
  assign t_r30_c8_6 = t_r30_c8_1 + p_29_9;
  assign t_r30_c8_7 = t_r30_c8_2 + t_r30_c8_3;
  assign t_r30_c8_8 = t_r30_c8_4 + p_31_7;
  assign t_r30_c8_9 = t_r30_c8_5 + t_r30_c8_6;
  assign t_r30_c8_10 = t_r30_c8_7 + t_r30_c8_8;
  assign t_r30_c8_11 = t_r30_c8_9 + t_r30_c8_10;
  assign t_r30_c8_12 = t_r30_c8_11 + p_31_9;
  assign out_30_8 = t_r30_c8_12 >> 4;

  assign t_r30_c9_0 = p_29_9 << 1;
  assign t_r30_c9_1 = p_30_8 << 1;
  assign t_r30_c9_2 = p_30_9 << 2;
  assign t_r30_c9_3 = p_30_10 << 1;
  assign t_r30_c9_4 = p_31_9 << 1;
  assign t_r30_c9_5 = t_r30_c9_0 + p_29_8;
  assign t_r30_c9_6 = t_r30_c9_1 + p_29_10;
  assign t_r30_c9_7 = t_r30_c9_2 + t_r30_c9_3;
  assign t_r30_c9_8 = t_r30_c9_4 + p_31_8;
  assign t_r30_c9_9 = t_r30_c9_5 + t_r30_c9_6;
  assign t_r30_c9_10 = t_r30_c9_7 + t_r30_c9_8;
  assign t_r30_c9_11 = t_r30_c9_9 + t_r30_c9_10;
  assign t_r30_c9_12 = t_r30_c9_11 + p_31_10;
  assign out_30_9 = t_r30_c9_12 >> 4;

  assign t_r30_c10_0 = p_29_10 << 1;
  assign t_r30_c10_1 = p_30_9 << 1;
  assign t_r30_c10_2 = p_30_10 << 2;
  assign t_r30_c10_3 = p_30_11 << 1;
  assign t_r30_c10_4 = p_31_10 << 1;
  assign t_r30_c10_5 = t_r30_c10_0 + p_29_9;
  assign t_r30_c10_6 = t_r30_c10_1 + p_29_11;
  assign t_r30_c10_7 = t_r30_c10_2 + t_r30_c10_3;
  assign t_r30_c10_8 = t_r30_c10_4 + p_31_9;
  assign t_r30_c10_9 = t_r30_c10_5 + t_r30_c10_6;
  assign t_r30_c10_10 = t_r30_c10_7 + t_r30_c10_8;
  assign t_r30_c10_11 = t_r30_c10_9 + t_r30_c10_10;
  assign t_r30_c10_12 = t_r30_c10_11 + p_31_11;
  assign out_30_10 = t_r30_c10_12 >> 4;

  assign t_r30_c11_0 = p_29_11 << 1;
  assign t_r30_c11_1 = p_30_10 << 1;
  assign t_r30_c11_2 = p_30_11 << 2;
  assign t_r30_c11_3 = p_30_12 << 1;
  assign t_r30_c11_4 = p_31_11 << 1;
  assign t_r30_c11_5 = t_r30_c11_0 + p_29_10;
  assign t_r30_c11_6 = t_r30_c11_1 + p_29_12;
  assign t_r30_c11_7 = t_r30_c11_2 + t_r30_c11_3;
  assign t_r30_c11_8 = t_r30_c11_4 + p_31_10;
  assign t_r30_c11_9 = t_r30_c11_5 + t_r30_c11_6;
  assign t_r30_c11_10 = t_r30_c11_7 + t_r30_c11_8;
  assign t_r30_c11_11 = t_r30_c11_9 + t_r30_c11_10;
  assign t_r30_c11_12 = t_r30_c11_11 + p_31_12;
  assign out_30_11 = t_r30_c11_12 >> 4;

  assign t_r30_c12_0 = p_29_12 << 1;
  assign t_r30_c12_1 = p_30_11 << 1;
  assign t_r30_c12_2 = p_30_12 << 2;
  assign t_r30_c12_3 = p_30_13 << 1;
  assign t_r30_c12_4 = p_31_12 << 1;
  assign t_r30_c12_5 = t_r30_c12_0 + p_29_11;
  assign t_r30_c12_6 = t_r30_c12_1 + p_29_13;
  assign t_r30_c12_7 = t_r30_c12_2 + t_r30_c12_3;
  assign t_r30_c12_8 = t_r30_c12_4 + p_31_11;
  assign t_r30_c12_9 = t_r30_c12_5 + t_r30_c12_6;
  assign t_r30_c12_10 = t_r30_c12_7 + t_r30_c12_8;
  assign t_r30_c12_11 = t_r30_c12_9 + t_r30_c12_10;
  assign t_r30_c12_12 = t_r30_c12_11 + p_31_13;
  assign out_30_12 = t_r30_c12_12 >> 4;

  assign t_r30_c13_0 = p_29_13 << 1;
  assign t_r30_c13_1 = p_30_12 << 1;
  assign t_r30_c13_2 = p_30_13 << 2;
  assign t_r30_c13_3 = p_30_14 << 1;
  assign t_r30_c13_4 = p_31_13 << 1;
  assign t_r30_c13_5 = t_r30_c13_0 + p_29_12;
  assign t_r30_c13_6 = t_r30_c13_1 + p_29_14;
  assign t_r30_c13_7 = t_r30_c13_2 + t_r30_c13_3;
  assign t_r30_c13_8 = t_r30_c13_4 + p_31_12;
  assign t_r30_c13_9 = t_r30_c13_5 + t_r30_c13_6;
  assign t_r30_c13_10 = t_r30_c13_7 + t_r30_c13_8;
  assign t_r30_c13_11 = t_r30_c13_9 + t_r30_c13_10;
  assign t_r30_c13_12 = t_r30_c13_11 + p_31_14;
  assign out_30_13 = t_r30_c13_12 >> 4;

  assign t_r30_c14_0 = p_29_14 << 1;
  assign t_r30_c14_1 = p_30_13 << 1;
  assign t_r30_c14_2 = p_30_14 << 2;
  assign t_r30_c14_3 = p_30_15 << 1;
  assign t_r30_c14_4 = p_31_14 << 1;
  assign t_r30_c14_5 = t_r30_c14_0 + p_29_13;
  assign t_r30_c14_6 = t_r30_c14_1 + p_29_15;
  assign t_r30_c14_7 = t_r30_c14_2 + t_r30_c14_3;
  assign t_r30_c14_8 = t_r30_c14_4 + p_31_13;
  assign t_r30_c14_9 = t_r30_c14_5 + t_r30_c14_6;
  assign t_r30_c14_10 = t_r30_c14_7 + t_r30_c14_8;
  assign t_r30_c14_11 = t_r30_c14_9 + t_r30_c14_10;
  assign t_r30_c14_12 = t_r30_c14_11 + p_31_15;
  assign out_30_14 = t_r30_c14_12 >> 4;

  assign t_r30_c15_0 = p_29_15 << 1;
  assign t_r30_c15_1 = p_30_14 << 1;
  assign t_r30_c15_2 = p_30_15 << 2;
  assign t_r30_c15_3 = p_30_16 << 1;
  assign t_r30_c15_4 = p_31_15 << 1;
  assign t_r30_c15_5 = t_r30_c15_0 + p_29_14;
  assign t_r30_c15_6 = t_r30_c15_1 + p_29_16;
  assign t_r30_c15_7 = t_r30_c15_2 + t_r30_c15_3;
  assign t_r30_c15_8 = t_r30_c15_4 + p_31_14;
  assign t_r30_c15_9 = t_r30_c15_5 + t_r30_c15_6;
  assign t_r30_c15_10 = t_r30_c15_7 + t_r30_c15_8;
  assign t_r30_c15_11 = t_r30_c15_9 + t_r30_c15_10;
  assign t_r30_c15_12 = t_r30_c15_11 + p_31_16;
  assign out_30_15 = t_r30_c15_12 >> 4;

  assign t_r30_c16_0 = p_29_16 << 1;
  assign t_r30_c16_1 = p_30_15 << 1;
  assign t_r30_c16_2 = p_30_16 << 2;
  assign t_r30_c16_3 = p_30_17 << 1;
  assign t_r30_c16_4 = p_31_16 << 1;
  assign t_r30_c16_5 = t_r30_c16_0 + p_29_15;
  assign t_r30_c16_6 = t_r30_c16_1 + p_29_17;
  assign t_r30_c16_7 = t_r30_c16_2 + t_r30_c16_3;
  assign t_r30_c16_8 = t_r30_c16_4 + p_31_15;
  assign t_r30_c16_9 = t_r30_c16_5 + t_r30_c16_6;
  assign t_r30_c16_10 = t_r30_c16_7 + t_r30_c16_8;
  assign t_r30_c16_11 = t_r30_c16_9 + t_r30_c16_10;
  assign t_r30_c16_12 = t_r30_c16_11 + p_31_17;
  assign out_30_16 = t_r30_c16_12 >> 4;

  assign t_r30_c17_0 = p_29_17 << 1;
  assign t_r30_c17_1 = p_30_16 << 1;
  assign t_r30_c17_2 = p_30_17 << 2;
  assign t_r30_c17_3 = p_30_18 << 1;
  assign t_r30_c17_4 = p_31_17 << 1;
  assign t_r30_c17_5 = t_r30_c17_0 + p_29_16;
  assign t_r30_c17_6 = t_r30_c17_1 + p_29_18;
  assign t_r30_c17_7 = t_r30_c17_2 + t_r30_c17_3;
  assign t_r30_c17_8 = t_r30_c17_4 + p_31_16;
  assign t_r30_c17_9 = t_r30_c17_5 + t_r30_c17_6;
  assign t_r30_c17_10 = t_r30_c17_7 + t_r30_c17_8;
  assign t_r30_c17_11 = t_r30_c17_9 + t_r30_c17_10;
  assign t_r30_c17_12 = t_r30_c17_11 + p_31_18;
  assign out_30_17 = t_r30_c17_12 >> 4;

  assign t_r30_c18_0 = p_29_18 << 1;
  assign t_r30_c18_1 = p_30_17 << 1;
  assign t_r30_c18_2 = p_30_18 << 2;
  assign t_r30_c18_3 = p_30_19 << 1;
  assign t_r30_c18_4 = p_31_18 << 1;
  assign t_r30_c18_5 = t_r30_c18_0 + p_29_17;
  assign t_r30_c18_6 = t_r30_c18_1 + p_29_19;
  assign t_r30_c18_7 = t_r30_c18_2 + t_r30_c18_3;
  assign t_r30_c18_8 = t_r30_c18_4 + p_31_17;
  assign t_r30_c18_9 = t_r30_c18_5 + t_r30_c18_6;
  assign t_r30_c18_10 = t_r30_c18_7 + t_r30_c18_8;
  assign t_r30_c18_11 = t_r30_c18_9 + t_r30_c18_10;
  assign t_r30_c18_12 = t_r30_c18_11 + p_31_19;
  assign out_30_18 = t_r30_c18_12 >> 4;

  assign t_r30_c19_0 = p_29_19 << 1;
  assign t_r30_c19_1 = p_30_18 << 1;
  assign t_r30_c19_2 = p_30_19 << 2;
  assign t_r30_c19_3 = p_30_20 << 1;
  assign t_r30_c19_4 = p_31_19 << 1;
  assign t_r30_c19_5 = t_r30_c19_0 + p_29_18;
  assign t_r30_c19_6 = t_r30_c19_1 + p_29_20;
  assign t_r30_c19_7 = t_r30_c19_2 + t_r30_c19_3;
  assign t_r30_c19_8 = t_r30_c19_4 + p_31_18;
  assign t_r30_c19_9 = t_r30_c19_5 + t_r30_c19_6;
  assign t_r30_c19_10 = t_r30_c19_7 + t_r30_c19_8;
  assign t_r30_c19_11 = t_r30_c19_9 + t_r30_c19_10;
  assign t_r30_c19_12 = t_r30_c19_11 + p_31_20;
  assign out_30_19 = t_r30_c19_12 >> 4;

  assign t_r30_c20_0 = p_29_20 << 1;
  assign t_r30_c20_1 = p_30_19 << 1;
  assign t_r30_c20_2 = p_30_20 << 2;
  assign t_r30_c20_3 = p_30_21 << 1;
  assign t_r30_c20_4 = p_31_20 << 1;
  assign t_r30_c20_5 = t_r30_c20_0 + p_29_19;
  assign t_r30_c20_6 = t_r30_c20_1 + p_29_21;
  assign t_r30_c20_7 = t_r30_c20_2 + t_r30_c20_3;
  assign t_r30_c20_8 = t_r30_c20_4 + p_31_19;
  assign t_r30_c20_9 = t_r30_c20_5 + t_r30_c20_6;
  assign t_r30_c20_10 = t_r30_c20_7 + t_r30_c20_8;
  assign t_r30_c20_11 = t_r30_c20_9 + t_r30_c20_10;
  assign t_r30_c20_12 = t_r30_c20_11 + p_31_21;
  assign out_30_20 = t_r30_c20_12 >> 4;

  assign t_r30_c21_0 = p_29_21 << 1;
  assign t_r30_c21_1 = p_30_20 << 1;
  assign t_r30_c21_2 = p_30_21 << 2;
  assign t_r30_c21_3 = p_30_22 << 1;
  assign t_r30_c21_4 = p_31_21 << 1;
  assign t_r30_c21_5 = t_r30_c21_0 + p_29_20;
  assign t_r30_c21_6 = t_r30_c21_1 + p_29_22;
  assign t_r30_c21_7 = t_r30_c21_2 + t_r30_c21_3;
  assign t_r30_c21_8 = t_r30_c21_4 + p_31_20;
  assign t_r30_c21_9 = t_r30_c21_5 + t_r30_c21_6;
  assign t_r30_c21_10 = t_r30_c21_7 + t_r30_c21_8;
  assign t_r30_c21_11 = t_r30_c21_9 + t_r30_c21_10;
  assign t_r30_c21_12 = t_r30_c21_11 + p_31_22;
  assign out_30_21 = t_r30_c21_12 >> 4;

  assign t_r30_c22_0 = p_29_22 << 1;
  assign t_r30_c22_1 = p_30_21 << 1;
  assign t_r30_c22_2 = p_30_22 << 2;
  assign t_r30_c22_3 = p_30_23 << 1;
  assign t_r30_c22_4 = p_31_22 << 1;
  assign t_r30_c22_5 = t_r30_c22_0 + p_29_21;
  assign t_r30_c22_6 = t_r30_c22_1 + p_29_23;
  assign t_r30_c22_7 = t_r30_c22_2 + t_r30_c22_3;
  assign t_r30_c22_8 = t_r30_c22_4 + p_31_21;
  assign t_r30_c22_9 = t_r30_c22_5 + t_r30_c22_6;
  assign t_r30_c22_10 = t_r30_c22_7 + t_r30_c22_8;
  assign t_r30_c22_11 = t_r30_c22_9 + t_r30_c22_10;
  assign t_r30_c22_12 = t_r30_c22_11 + p_31_23;
  assign out_30_22 = t_r30_c22_12 >> 4;

  assign t_r30_c23_0 = p_29_23 << 1;
  assign t_r30_c23_1 = p_30_22 << 1;
  assign t_r30_c23_2 = p_30_23 << 2;
  assign t_r30_c23_3 = p_30_24 << 1;
  assign t_r30_c23_4 = p_31_23 << 1;
  assign t_r30_c23_5 = t_r30_c23_0 + p_29_22;
  assign t_r30_c23_6 = t_r30_c23_1 + p_29_24;
  assign t_r30_c23_7 = t_r30_c23_2 + t_r30_c23_3;
  assign t_r30_c23_8 = t_r30_c23_4 + p_31_22;
  assign t_r30_c23_9 = t_r30_c23_5 + t_r30_c23_6;
  assign t_r30_c23_10 = t_r30_c23_7 + t_r30_c23_8;
  assign t_r30_c23_11 = t_r30_c23_9 + t_r30_c23_10;
  assign t_r30_c23_12 = t_r30_c23_11 + p_31_24;
  assign out_30_23 = t_r30_c23_12 >> 4;

  assign t_r30_c24_0 = p_29_24 << 1;
  assign t_r30_c24_1 = p_30_23 << 1;
  assign t_r30_c24_2 = p_30_24 << 2;
  assign t_r30_c24_3 = p_30_25 << 1;
  assign t_r30_c24_4 = p_31_24 << 1;
  assign t_r30_c24_5 = t_r30_c24_0 + p_29_23;
  assign t_r30_c24_6 = t_r30_c24_1 + p_29_25;
  assign t_r30_c24_7 = t_r30_c24_2 + t_r30_c24_3;
  assign t_r30_c24_8 = t_r30_c24_4 + p_31_23;
  assign t_r30_c24_9 = t_r30_c24_5 + t_r30_c24_6;
  assign t_r30_c24_10 = t_r30_c24_7 + t_r30_c24_8;
  assign t_r30_c24_11 = t_r30_c24_9 + t_r30_c24_10;
  assign t_r30_c24_12 = t_r30_c24_11 + p_31_25;
  assign out_30_24 = t_r30_c24_12 >> 4;

  assign t_r30_c25_0 = p_29_25 << 1;
  assign t_r30_c25_1 = p_30_24 << 1;
  assign t_r30_c25_2 = p_30_25 << 2;
  assign t_r30_c25_3 = p_30_26 << 1;
  assign t_r30_c25_4 = p_31_25 << 1;
  assign t_r30_c25_5 = t_r30_c25_0 + p_29_24;
  assign t_r30_c25_6 = t_r30_c25_1 + p_29_26;
  assign t_r30_c25_7 = t_r30_c25_2 + t_r30_c25_3;
  assign t_r30_c25_8 = t_r30_c25_4 + p_31_24;
  assign t_r30_c25_9 = t_r30_c25_5 + t_r30_c25_6;
  assign t_r30_c25_10 = t_r30_c25_7 + t_r30_c25_8;
  assign t_r30_c25_11 = t_r30_c25_9 + t_r30_c25_10;
  assign t_r30_c25_12 = t_r30_c25_11 + p_31_26;
  assign out_30_25 = t_r30_c25_12 >> 4;

  assign t_r30_c26_0 = p_29_26 << 1;
  assign t_r30_c26_1 = p_30_25 << 1;
  assign t_r30_c26_2 = p_30_26 << 2;
  assign t_r30_c26_3 = p_30_27 << 1;
  assign t_r30_c26_4 = p_31_26 << 1;
  assign t_r30_c26_5 = t_r30_c26_0 + p_29_25;
  assign t_r30_c26_6 = t_r30_c26_1 + p_29_27;
  assign t_r30_c26_7 = t_r30_c26_2 + t_r30_c26_3;
  assign t_r30_c26_8 = t_r30_c26_4 + p_31_25;
  assign t_r30_c26_9 = t_r30_c26_5 + t_r30_c26_6;
  assign t_r30_c26_10 = t_r30_c26_7 + t_r30_c26_8;
  assign t_r30_c26_11 = t_r30_c26_9 + t_r30_c26_10;
  assign t_r30_c26_12 = t_r30_c26_11 + p_31_27;
  assign out_30_26 = t_r30_c26_12 >> 4;

  assign t_r30_c27_0 = p_29_27 << 1;
  assign t_r30_c27_1 = p_30_26 << 1;
  assign t_r30_c27_2 = p_30_27 << 2;
  assign t_r30_c27_3 = p_30_28 << 1;
  assign t_r30_c27_4 = p_31_27 << 1;
  assign t_r30_c27_5 = t_r30_c27_0 + p_29_26;
  assign t_r30_c27_6 = t_r30_c27_1 + p_29_28;
  assign t_r30_c27_7 = t_r30_c27_2 + t_r30_c27_3;
  assign t_r30_c27_8 = t_r30_c27_4 + p_31_26;
  assign t_r30_c27_9 = t_r30_c27_5 + t_r30_c27_6;
  assign t_r30_c27_10 = t_r30_c27_7 + t_r30_c27_8;
  assign t_r30_c27_11 = t_r30_c27_9 + t_r30_c27_10;
  assign t_r30_c27_12 = t_r30_c27_11 + p_31_28;
  assign out_30_27 = t_r30_c27_12 >> 4;

  assign t_r30_c28_0 = p_29_28 << 1;
  assign t_r30_c28_1 = p_30_27 << 1;
  assign t_r30_c28_2 = p_30_28 << 2;
  assign t_r30_c28_3 = p_30_29 << 1;
  assign t_r30_c28_4 = p_31_28 << 1;
  assign t_r30_c28_5 = t_r30_c28_0 + p_29_27;
  assign t_r30_c28_6 = t_r30_c28_1 + p_29_29;
  assign t_r30_c28_7 = t_r30_c28_2 + t_r30_c28_3;
  assign t_r30_c28_8 = t_r30_c28_4 + p_31_27;
  assign t_r30_c28_9 = t_r30_c28_5 + t_r30_c28_6;
  assign t_r30_c28_10 = t_r30_c28_7 + t_r30_c28_8;
  assign t_r30_c28_11 = t_r30_c28_9 + t_r30_c28_10;
  assign t_r30_c28_12 = t_r30_c28_11 + p_31_29;
  assign out_30_28 = t_r30_c28_12 >> 4;

  assign t_r30_c29_0 = p_29_29 << 1;
  assign t_r30_c29_1 = p_30_28 << 1;
  assign t_r30_c29_2 = p_30_29 << 2;
  assign t_r30_c29_3 = p_30_30 << 1;
  assign t_r30_c29_4 = p_31_29 << 1;
  assign t_r30_c29_5 = t_r30_c29_0 + p_29_28;
  assign t_r30_c29_6 = t_r30_c29_1 + p_29_30;
  assign t_r30_c29_7 = t_r30_c29_2 + t_r30_c29_3;
  assign t_r30_c29_8 = t_r30_c29_4 + p_31_28;
  assign t_r30_c29_9 = t_r30_c29_5 + t_r30_c29_6;
  assign t_r30_c29_10 = t_r30_c29_7 + t_r30_c29_8;
  assign t_r30_c29_11 = t_r30_c29_9 + t_r30_c29_10;
  assign t_r30_c29_12 = t_r30_c29_11 + p_31_30;
  assign out_30_29 = t_r30_c29_12 >> 4;

  assign t_r30_c30_0 = p_29_30 << 1;
  assign t_r30_c30_1 = p_30_29 << 1;
  assign t_r30_c30_2 = p_30_30 << 2;
  assign t_r30_c30_3 = p_30_31 << 1;
  assign t_r30_c30_4 = p_31_30 << 1;
  assign t_r30_c30_5 = t_r30_c30_0 + p_29_29;
  assign t_r30_c30_6 = t_r30_c30_1 + p_29_31;
  assign t_r30_c30_7 = t_r30_c30_2 + t_r30_c30_3;
  assign t_r30_c30_8 = t_r30_c30_4 + p_31_29;
  assign t_r30_c30_9 = t_r30_c30_5 + t_r30_c30_6;
  assign t_r30_c30_10 = t_r30_c30_7 + t_r30_c30_8;
  assign t_r30_c30_11 = t_r30_c30_9 + t_r30_c30_10;
  assign t_r30_c30_12 = t_r30_c30_11 + p_31_31;
  assign out_30_30 = t_r30_c30_12 >> 4;

  assign t_r30_c31_0 = p_29_31 << 1;
  assign t_r30_c31_1 = p_30_30 << 1;
  assign t_r30_c31_2 = p_30_31 << 2;
  assign t_r30_c31_3 = p_30_32 << 1;
  assign t_r30_c31_4 = p_31_31 << 1;
  assign t_r30_c31_5 = t_r30_c31_0 + p_29_30;
  assign t_r30_c31_6 = t_r30_c31_1 + p_29_32;
  assign t_r30_c31_7 = t_r30_c31_2 + t_r30_c31_3;
  assign t_r30_c31_8 = t_r30_c31_4 + p_31_30;
  assign t_r30_c31_9 = t_r30_c31_5 + t_r30_c31_6;
  assign t_r30_c31_10 = t_r30_c31_7 + t_r30_c31_8;
  assign t_r30_c31_11 = t_r30_c31_9 + t_r30_c31_10;
  assign t_r30_c31_12 = t_r30_c31_11 + p_31_32;
  assign out_30_31 = t_r30_c31_12 >> 4;

  assign t_r30_c32_0 = p_29_32 << 1;
  assign t_r30_c32_1 = p_30_31 << 1;
  assign t_r30_c32_2 = p_30_32 << 2;
  assign t_r30_c32_3 = p_30_33 << 1;
  assign t_r30_c32_4 = p_31_32 << 1;
  assign t_r30_c32_5 = t_r30_c32_0 + p_29_31;
  assign t_r30_c32_6 = t_r30_c32_1 + p_29_33;
  assign t_r30_c32_7 = t_r30_c32_2 + t_r30_c32_3;
  assign t_r30_c32_8 = t_r30_c32_4 + p_31_31;
  assign t_r30_c32_9 = t_r30_c32_5 + t_r30_c32_6;
  assign t_r30_c32_10 = t_r30_c32_7 + t_r30_c32_8;
  assign t_r30_c32_11 = t_r30_c32_9 + t_r30_c32_10;
  assign t_r30_c32_12 = t_r30_c32_11 + p_31_33;
  assign out_30_32 = t_r30_c32_12 >> 4;

  assign t_r30_c33_0 = p_29_33 << 1;
  assign t_r30_c33_1 = p_30_32 << 1;
  assign t_r30_c33_2 = p_30_33 << 2;
  assign t_r30_c33_3 = p_30_34 << 1;
  assign t_r30_c33_4 = p_31_33 << 1;
  assign t_r30_c33_5 = t_r30_c33_0 + p_29_32;
  assign t_r30_c33_6 = t_r30_c33_1 + p_29_34;
  assign t_r30_c33_7 = t_r30_c33_2 + t_r30_c33_3;
  assign t_r30_c33_8 = t_r30_c33_4 + p_31_32;
  assign t_r30_c33_9 = t_r30_c33_5 + t_r30_c33_6;
  assign t_r30_c33_10 = t_r30_c33_7 + t_r30_c33_8;
  assign t_r30_c33_11 = t_r30_c33_9 + t_r30_c33_10;
  assign t_r30_c33_12 = t_r30_c33_11 + p_31_34;
  assign out_30_33 = t_r30_c33_12 >> 4;

  assign t_r30_c34_0 = p_29_34 << 1;
  assign t_r30_c34_1 = p_30_33 << 1;
  assign t_r30_c34_2 = p_30_34 << 2;
  assign t_r30_c34_3 = p_30_35 << 1;
  assign t_r30_c34_4 = p_31_34 << 1;
  assign t_r30_c34_5 = t_r30_c34_0 + p_29_33;
  assign t_r30_c34_6 = t_r30_c34_1 + p_29_35;
  assign t_r30_c34_7 = t_r30_c34_2 + t_r30_c34_3;
  assign t_r30_c34_8 = t_r30_c34_4 + p_31_33;
  assign t_r30_c34_9 = t_r30_c34_5 + t_r30_c34_6;
  assign t_r30_c34_10 = t_r30_c34_7 + t_r30_c34_8;
  assign t_r30_c34_11 = t_r30_c34_9 + t_r30_c34_10;
  assign t_r30_c34_12 = t_r30_c34_11 + p_31_35;
  assign out_30_34 = t_r30_c34_12 >> 4;

  assign t_r30_c35_0 = p_29_35 << 1;
  assign t_r30_c35_1 = p_30_34 << 1;
  assign t_r30_c35_2 = p_30_35 << 2;
  assign t_r30_c35_3 = p_30_36 << 1;
  assign t_r30_c35_4 = p_31_35 << 1;
  assign t_r30_c35_5 = t_r30_c35_0 + p_29_34;
  assign t_r30_c35_6 = t_r30_c35_1 + p_29_36;
  assign t_r30_c35_7 = t_r30_c35_2 + t_r30_c35_3;
  assign t_r30_c35_8 = t_r30_c35_4 + p_31_34;
  assign t_r30_c35_9 = t_r30_c35_5 + t_r30_c35_6;
  assign t_r30_c35_10 = t_r30_c35_7 + t_r30_c35_8;
  assign t_r30_c35_11 = t_r30_c35_9 + t_r30_c35_10;
  assign t_r30_c35_12 = t_r30_c35_11 + p_31_36;
  assign out_30_35 = t_r30_c35_12 >> 4;

  assign t_r30_c36_0 = p_29_36 << 1;
  assign t_r30_c36_1 = p_30_35 << 1;
  assign t_r30_c36_2 = p_30_36 << 2;
  assign t_r30_c36_3 = p_30_37 << 1;
  assign t_r30_c36_4 = p_31_36 << 1;
  assign t_r30_c36_5 = t_r30_c36_0 + p_29_35;
  assign t_r30_c36_6 = t_r30_c36_1 + p_29_37;
  assign t_r30_c36_7 = t_r30_c36_2 + t_r30_c36_3;
  assign t_r30_c36_8 = t_r30_c36_4 + p_31_35;
  assign t_r30_c36_9 = t_r30_c36_5 + t_r30_c36_6;
  assign t_r30_c36_10 = t_r30_c36_7 + t_r30_c36_8;
  assign t_r30_c36_11 = t_r30_c36_9 + t_r30_c36_10;
  assign t_r30_c36_12 = t_r30_c36_11 + p_31_37;
  assign out_30_36 = t_r30_c36_12 >> 4;

  assign t_r30_c37_0 = p_29_37 << 1;
  assign t_r30_c37_1 = p_30_36 << 1;
  assign t_r30_c37_2 = p_30_37 << 2;
  assign t_r30_c37_3 = p_30_38 << 1;
  assign t_r30_c37_4 = p_31_37 << 1;
  assign t_r30_c37_5 = t_r30_c37_0 + p_29_36;
  assign t_r30_c37_6 = t_r30_c37_1 + p_29_38;
  assign t_r30_c37_7 = t_r30_c37_2 + t_r30_c37_3;
  assign t_r30_c37_8 = t_r30_c37_4 + p_31_36;
  assign t_r30_c37_9 = t_r30_c37_5 + t_r30_c37_6;
  assign t_r30_c37_10 = t_r30_c37_7 + t_r30_c37_8;
  assign t_r30_c37_11 = t_r30_c37_9 + t_r30_c37_10;
  assign t_r30_c37_12 = t_r30_c37_11 + p_31_38;
  assign out_30_37 = t_r30_c37_12 >> 4;

  assign t_r30_c38_0 = p_29_38 << 1;
  assign t_r30_c38_1 = p_30_37 << 1;
  assign t_r30_c38_2 = p_30_38 << 2;
  assign t_r30_c38_3 = p_30_39 << 1;
  assign t_r30_c38_4 = p_31_38 << 1;
  assign t_r30_c38_5 = t_r30_c38_0 + p_29_37;
  assign t_r30_c38_6 = t_r30_c38_1 + p_29_39;
  assign t_r30_c38_7 = t_r30_c38_2 + t_r30_c38_3;
  assign t_r30_c38_8 = t_r30_c38_4 + p_31_37;
  assign t_r30_c38_9 = t_r30_c38_5 + t_r30_c38_6;
  assign t_r30_c38_10 = t_r30_c38_7 + t_r30_c38_8;
  assign t_r30_c38_11 = t_r30_c38_9 + t_r30_c38_10;
  assign t_r30_c38_12 = t_r30_c38_11 + p_31_39;
  assign out_30_38 = t_r30_c38_12 >> 4;

  assign t_r30_c39_0 = p_29_39 << 1;
  assign t_r30_c39_1 = p_30_38 << 1;
  assign t_r30_c39_2 = p_30_39 << 2;
  assign t_r30_c39_3 = p_30_40 << 1;
  assign t_r30_c39_4 = p_31_39 << 1;
  assign t_r30_c39_5 = t_r30_c39_0 + p_29_38;
  assign t_r30_c39_6 = t_r30_c39_1 + p_29_40;
  assign t_r30_c39_7 = t_r30_c39_2 + t_r30_c39_3;
  assign t_r30_c39_8 = t_r30_c39_4 + p_31_38;
  assign t_r30_c39_9 = t_r30_c39_5 + t_r30_c39_6;
  assign t_r30_c39_10 = t_r30_c39_7 + t_r30_c39_8;
  assign t_r30_c39_11 = t_r30_c39_9 + t_r30_c39_10;
  assign t_r30_c39_12 = t_r30_c39_11 + p_31_40;
  assign out_30_39 = t_r30_c39_12 >> 4;

  assign t_r30_c40_0 = p_29_40 << 1;
  assign t_r30_c40_1 = p_30_39 << 1;
  assign t_r30_c40_2 = p_30_40 << 2;
  assign t_r30_c40_3 = p_30_41 << 1;
  assign t_r30_c40_4 = p_31_40 << 1;
  assign t_r30_c40_5 = t_r30_c40_0 + p_29_39;
  assign t_r30_c40_6 = t_r30_c40_1 + p_29_41;
  assign t_r30_c40_7 = t_r30_c40_2 + t_r30_c40_3;
  assign t_r30_c40_8 = t_r30_c40_4 + p_31_39;
  assign t_r30_c40_9 = t_r30_c40_5 + t_r30_c40_6;
  assign t_r30_c40_10 = t_r30_c40_7 + t_r30_c40_8;
  assign t_r30_c40_11 = t_r30_c40_9 + t_r30_c40_10;
  assign t_r30_c40_12 = t_r30_c40_11 + p_31_41;
  assign out_30_40 = t_r30_c40_12 >> 4;

  assign t_r30_c41_0 = p_29_41 << 1;
  assign t_r30_c41_1 = p_30_40 << 1;
  assign t_r30_c41_2 = p_30_41 << 2;
  assign t_r30_c41_3 = p_30_42 << 1;
  assign t_r30_c41_4 = p_31_41 << 1;
  assign t_r30_c41_5 = t_r30_c41_0 + p_29_40;
  assign t_r30_c41_6 = t_r30_c41_1 + p_29_42;
  assign t_r30_c41_7 = t_r30_c41_2 + t_r30_c41_3;
  assign t_r30_c41_8 = t_r30_c41_4 + p_31_40;
  assign t_r30_c41_9 = t_r30_c41_5 + t_r30_c41_6;
  assign t_r30_c41_10 = t_r30_c41_7 + t_r30_c41_8;
  assign t_r30_c41_11 = t_r30_c41_9 + t_r30_c41_10;
  assign t_r30_c41_12 = t_r30_c41_11 + p_31_42;
  assign out_30_41 = t_r30_c41_12 >> 4;

  assign t_r30_c42_0 = p_29_42 << 1;
  assign t_r30_c42_1 = p_30_41 << 1;
  assign t_r30_c42_2 = p_30_42 << 2;
  assign t_r30_c42_3 = p_30_43 << 1;
  assign t_r30_c42_4 = p_31_42 << 1;
  assign t_r30_c42_5 = t_r30_c42_0 + p_29_41;
  assign t_r30_c42_6 = t_r30_c42_1 + p_29_43;
  assign t_r30_c42_7 = t_r30_c42_2 + t_r30_c42_3;
  assign t_r30_c42_8 = t_r30_c42_4 + p_31_41;
  assign t_r30_c42_9 = t_r30_c42_5 + t_r30_c42_6;
  assign t_r30_c42_10 = t_r30_c42_7 + t_r30_c42_8;
  assign t_r30_c42_11 = t_r30_c42_9 + t_r30_c42_10;
  assign t_r30_c42_12 = t_r30_c42_11 + p_31_43;
  assign out_30_42 = t_r30_c42_12 >> 4;

  assign t_r30_c43_0 = p_29_43 << 1;
  assign t_r30_c43_1 = p_30_42 << 1;
  assign t_r30_c43_2 = p_30_43 << 2;
  assign t_r30_c43_3 = p_30_44 << 1;
  assign t_r30_c43_4 = p_31_43 << 1;
  assign t_r30_c43_5 = t_r30_c43_0 + p_29_42;
  assign t_r30_c43_6 = t_r30_c43_1 + p_29_44;
  assign t_r30_c43_7 = t_r30_c43_2 + t_r30_c43_3;
  assign t_r30_c43_8 = t_r30_c43_4 + p_31_42;
  assign t_r30_c43_9 = t_r30_c43_5 + t_r30_c43_6;
  assign t_r30_c43_10 = t_r30_c43_7 + t_r30_c43_8;
  assign t_r30_c43_11 = t_r30_c43_9 + t_r30_c43_10;
  assign t_r30_c43_12 = t_r30_c43_11 + p_31_44;
  assign out_30_43 = t_r30_c43_12 >> 4;

  assign t_r30_c44_0 = p_29_44 << 1;
  assign t_r30_c44_1 = p_30_43 << 1;
  assign t_r30_c44_2 = p_30_44 << 2;
  assign t_r30_c44_3 = p_30_45 << 1;
  assign t_r30_c44_4 = p_31_44 << 1;
  assign t_r30_c44_5 = t_r30_c44_0 + p_29_43;
  assign t_r30_c44_6 = t_r30_c44_1 + p_29_45;
  assign t_r30_c44_7 = t_r30_c44_2 + t_r30_c44_3;
  assign t_r30_c44_8 = t_r30_c44_4 + p_31_43;
  assign t_r30_c44_9 = t_r30_c44_5 + t_r30_c44_6;
  assign t_r30_c44_10 = t_r30_c44_7 + t_r30_c44_8;
  assign t_r30_c44_11 = t_r30_c44_9 + t_r30_c44_10;
  assign t_r30_c44_12 = t_r30_c44_11 + p_31_45;
  assign out_30_44 = t_r30_c44_12 >> 4;

  assign t_r30_c45_0 = p_29_45 << 1;
  assign t_r30_c45_1 = p_30_44 << 1;
  assign t_r30_c45_2 = p_30_45 << 2;
  assign t_r30_c45_3 = p_30_46 << 1;
  assign t_r30_c45_4 = p_31_45 << 1;
  assign t_r30_c45_5 = t_r30_c45_0 + p_29_44;
  assign t_r30_c45_6 = t_r30_c45_1 + p_29_46;
  assign t_r30_c45_7 = t_r30_c45_2 + t_r30_c45_3;
  assign t_r30_c45_8 = t_r30_c45_4 + p_31_44;
  assign t_r30_c45_9 = t_r30_c45_5 + t_r30_c45_6;
  assign t_r30_c45_10 = t_r30_c45_7 + t_r30_c45_8;
  assign t_r30_c45_11 = t_r30_c45_9 + t_r30_c45_10;
  assign t_r30_c45_12 = t_r30_c45_11 + p_31_46;
  assign out_30_45 = t_r30_c45_12 >> 4;

  assign t_r30_c46_0 = p_29_46 << 1;
  assign t_r30_c46_1 = p_30_45 << 1;
  assign t_r30_c46_2 = p_30_46 << 2;
  assign t_r30_c46_3 = p_30_47 << 1;
  assign t_r30_c46_4 = p_31_46 << 1;
  assign t_r30_c46_5 = t_r30_c46_0 + p_29_45;
  assign t_r30_c46_6 = t_r30_c46_1 + p_29_47;
  assign t_r30_c46_7 = t_r30_c46_2 + t_r30_c46_3;
  assign t_r30_c46_8 = t_r30_c46_4 + p_31_45;
  assign t_r30_c46_9 = t_r30_c46_5 + t_r30_c46_6;
  assign t_r30_c46_10 = t_r30_c46_7 + t_r30_c46_8;
  assign t_r30_c46_11 = t_r30_c46_9 + t_r30_c46_10;
  assign t_r30_c46_12 = t_r30_c46_11 + p_31_47;
  assign out_30_46 = t_r30_c46_12 >> 4;

  assign t_r30_c47_0 = p_29_47 << 1;
  assign t_r30_c47_1 = p_30_46 << 1;
  assign t_r30_c47_2 = p_30_47 << 2;
  assign t_r30_c47_3 = p_30_48 << 1;
  assign t_r30_c47_4 = p_31_47 << 1;
  assign t_r30_c47_5 = t_r30_c47_0 + p_29_46;
  assign t_r30_c47_6 = t_r30_c47_1 + p_29_48;
  assign t_r30_c47_7 = t_r30_c47_2 + t_r30_c47_3;
  assign t_r30_c47_8 = t_r30_c47_4 + p_31_46;
  assign t_r30_c47_9 = t_r30_c47_5 + t_r30_c47_6;
  assign t_r30_c47_10 = t_r30_c47_7 + t_r30_c47_8;
  assign t_r30_c47_11 = t_r30_c47_9 + t_r30_c47_10;
  assign t_r30_c47_12 = t_r30_c47_11 + p_31_48;
  assign out_30_47 = t_r30_c47_12 >> 4;

  assign t_r30_c48_0 = p_29_48 << 1;
  assign t_r30_c48_1 = p_30_47 << 1;
  assign t_r30_c48_2 = p_30_48 << 2;
  assign t_r30_c48_3 = p_30_49 << 1;
  assign t_r30_c48_4 = p_31_48 << 1;
  assign t_r30_c48_5 = t_r30_c48_0 + p_29_47;
  assign t_r30_c48_6 = t_r30_c48_1 + p_29_49;
  assign t_r30_c48_7 = t_r30_c48_2 + t_r30_c48_3;
  assign t_r30_c48_8 = t_r30_c48_4 + p_31_47;
  assign t_r30_c48_9 = t_r30_c48_5 + t_r30_c48_6;
  assign t_r30_c48_10 = t_r30_c48_7 + t_r30_c48_8;
  assign t_r30_c48_11 = t_r30_c48_9 + t_r30_c48_10;
  assign t_r30_c48_12 = t_r30_c48_11 + p_31_49;
  assign out_30_48 = t_r30_c48_12 >> 4;

  assign t_r30_c49_0 = p_29_49 << 1;
  assign t_r30_c49_1 = p_30_48 << 1;
  assign t_r30_c49_2 = p_30_49 << 2;
  assign t_r30_c49_3 = p_30_50 << 1;
  assign t_r30_c49_4 = p_31_49 << 1;
  assign t_r30_c49_5 = t_r30_c49_0 + p_29_48;
  assign t_r30_c49_6 = t_r30_c49_1 + p_29_50;
  assign t_r30_c49_7 = t_r30_c49_2 + t_r30_c49_3;
  assign t_r30_c49_8 = t_r30_c49_4 + p_31_48;
  assign t_r30_c49_9 = t_r30_c49_5 + t_r30_c49_6;
  assign t_r30_c49_10 = t_r30_c49_7 + t_r30_c49_8;
  assign t_r30_c49_11 = t_r30_c49_9 + t_r30_c49_10;
  assign t_r30_c49_12 = t_r30_c49_11 + p_31_50;
  assign out_30_49 = t_r30_c49_12 >> 4;

  assign t_r30_c50_0 = p_29_50 << 1;
  assign t_r30_c50_1 = p_30_49 << 1;
  assign t_r30_c50_2 = p_30_50 << 2;
  assign t_r30_c50_3 = p_30_51 << 1;
  assign t_r30_c50_4 = p_31_50 << 1;
  assign t_r30_c50_5 = t_r30_c50_0 + p_29_49;
  assign t_r30_c50_6 = t_r30_c50_1 + p_29_51;
  assign t_r30_c50_7 = t_r30_c50_2 + t_r30_c50_3;
  assign t_r30_c50_8 = t_r30_c50_4 + p_31_49;
  assign t_r30_c50_9 = t_r30_c50_5 + t_r30_c50_6;
  assign t_r30_c50_10 = t_r30_c50_7 + t_r30_c50_8;
  assign t_r30_c50_11 = t_r30_c50_9 + t_r30_c50_10;
  assign t_r30_c50_12 = t_r30_c50_11 + p_31_51;
  assign out_30_50 = t_r30_c50_12 >> 4;

  assign t_r30_c51_0 = p_29_51 << 1;
  assign t_r30_c51_1 = p_30_50 << 1;
  assign t_r30_c51_2 = p_30_51 << 2;
  assign t_r30_c51_3 = p_30_52 << 1;
  assign t_r30_c51_4 = p_31_51 << 1;
  assign t_r30_c51_5 = t_r30_c51_0 + p_29_50;
  assign t_r30_c51_6 = t_r30_c51_1 + p_29_52;
  assign t_r30_c51_7 = t_r30_c51_2 + t_r30_c51_3;
  assign t_r30_c51_8 = t_r30_c51_4 + p_31_50;
  assign t_r30_c51_9 = t_r30_c51_5 + t_r30_c51_6;
  assign t_r30_c51_10 = t_r30_c51_7 + t_r30_c51_8;
  assign t_r30_c51_11 = t_r30_c51_9 + t_r30_c51_10;
  assign t_r30_c51_12 = t_r30_c51_11 + p_31_52;
  assign out_30_51 = t_r30_c51_12 >> 4;

  assign t_r30_c52_0 = p_29_52 << 1;
  assign t_r30_c52_1 = p_30_51 << 1;
  assign t_r30_c52_2 = p_30_52 << 2;
  assign t_r30_c52_3 = p_30_53 << 1;
  assign t_r30_c52_4 = p_31_52 << 1;
  assign t_r30_c52_5 = t_r30_c52_0 + p_29_51;
  assign t_r30_c52_6 = t_r30_c52_1 + p_29_53;
  assign t_r30_c52_7 = t_r30_c52_2 + t_r30_c52_3;
  assign t_r30_c52_8 = t_r30_c52_4 + p_31_51;
  assign t_r30_c52_9 = t_r30_c52_5 + t_r30_c52_6;
  assign t_r30_c52_10 = t_r30_c52_7 + t_r30_c52_8;
  assign t_r30_c52_11 = t_r30_c52_9 + t_r30_c52_10;
  assign t_r30_c52_12 = t_r30_c52_11 + p_31_53;
  assign out_30_52 = t_r30_c52_12 >> 4;

  assign t_r30_c53_0 = p_29_53 << 1;
  assign t_r30_c53_1 = p_30_52 << 1;
  assign t_r30_c53_2 = p_30_53 << 2;
  assign t_r30_c53_3 = p_30_54 << 1;
  assign t_r30_c53_4 = p_31_53 << 1;
  assign t_r30_c53_5 = t_r30_c53_0 + p_29_52;
  assign t_r30_c53_6 = t_r30_c53_1 + p_29_54;
  assign t_r30_c53_7 = t_r30_c53_2 + t_r30_c53_3;
  assign t_r30_c53_8 = t_r30_c53_4 + p_31_52;
  assign t_r30_c53_9 = t_r30_c53_5 + t_r30_c53_6;
  assign t_r30_c53_10 = t_r30_c53_7 + t_r30_c53_8;
  assign t_r30_c53_11 = t_r30_c53_9 + t_r30_c53_10;
  assign t_r30_c53_12 = t_r30_c53_11 + p_31_54;
  assign out_30_53 = t_r30_c53_12 >> 4;

  assign t_r30_c54_0 = p_29_54 << 1;
  assign t_r30_c54_1 = p_30_53 << 1;
  assign t_r30_c54_2 = p_30_54 << 2;
  assign t_r30_c54_3 = p_30_55 << 1;
  assign t_r30_c54_4 = p_31_54 << 1;
  assign t_r30_c54_5 = t_r30_c54_0 + p_29_53;
  assign t_r30_c54_6 = t_r30_c54_1 + p_29_55;
  assign t_r30_c54_7 = t_r30_c54_2 + t_r30_c54_3;
  assign t_r30_c54_8 = t_r30_c54_4 + p_31_53;
  assign t_r30_c54_9 = t_r30_c54_5 + t_r30_c54_6;
  assign t_r30_c54_10 = t_r30_c54_7 + t_r30_c54_8;
  assign t_r30_c54_11 = t_r30_c54_9 + t_r30_c54_10;
  assign t_r30_c54_12 = t_r30_c54_11 + p_31_55;
  assign out_30_54 = t_r30_c54_12 >> 4;

  assign t_r30_c55_0 = p_29_55 << 1;
  assign t_r30_c55_1 = p_30_54 << 1;
  assign t_r30_c55_2 = p_30_55 << 2;
  assign t_r30_c55_3 = p_30_56 << 1;
  assign t_r30_c55_4 = p_31_55 << 1;
  assign t_r30_c55_5 = t_r30_c55_0 + p_29_54;
  assign t_r30_c55_6 = t_r30_c55_1 + p_29_56;
  assign t_r30_c55_7 = t_r30_c55_2 + t_r30_c55_3;
  assign t_r30_c55_8 = t_r30_c55_4 + p_31_54;
  assign t_r30_c55_9 = t_r30_c55_5 + t_r30_c55_6;
  assign t_r30_c55_10 = t_r30_c55_7 + t_r30_c55_8;
  assign t_r30_c55_11 = t_r30_c55_9 + t_r30_c55_10;
  assign t_r30_c55_12 = t_r30_c55_11 + p_31_56;
  assign out_30_55 = t_r30_c55_12 >> 4;

  assign t_r30_c56_0 = p_29_56 << 1;
  assign t_r30_c56_1 = p_30_55 << 1;
  assign t_r30_c56_2 = p_30_56 << 2;
  assign t_r30_c56_3 = p_30_57 << 1;
  assign t_r30_c56_4 = p_31_56 << 1;
  assign t_r30_c56_5 = t_r30_c56_0 + p_29_55;
  assign t_r30_c56_6 = t_r30_c56_1 + p_29_57;
  assign t_r30_c56_7 = t_r30_c56_2 + t_r30_c56_3;
  assign t_r30_c56_8 = t_r30_c56_4 + p_31_55;
  assign t_r30_c56_9 = t_r30_c56_5 + t_r30_c56_6;
  assign t_r30_c56_10 = t_r30_c56_7 + t_r30_c56_8;
  assign t_r30_c56_11 = t_r30_c56_9 + t_r30_c56_10;
  assign t_r30_c56_12 = t_r30_c56_11 + p_31_57;
  assign out_30_56 = t_r30_c56_12 >> 4;

  assign t_r30_c57_0 = p_29_57 << 1;
  assign t_r30_c57_1 = p_30_56 << 1;
  assign t_r30_c57_2 = p_30_57 << 2;
  assign t_r30_c57_3 = p_30_58 << 1;
  assign t_r30_c57_4 = p_31_57 << 1;
  assign t_r30_c57_5 = t_r30_c57_0 + p_29_56;
  assign t_r30_c57_6 = t_r30_c57_1 + p_29_58;
  assign t_r30_c57_7 = t_r30_c57_2 + t_r30_c57_3;
  assign t_r30_c57_8 = t_r30_c57_4 + p_31_56;
  assign t_r30_c57_9 = t_r30_c57_5 + t_r30_c57_6;
  assign t_r30_c57_10 = t_r30_c57_7 + t_r30_c57_8;
  assign t_r30_c57_11 = t_r30_c57_9 + t_r30_c57_10;
  assign t_r30_c57_12 = t_r30_c57_11 + p_31_58;
  assign out_30_57 = t_r30_c57_12 >> 4;

  assign t_r30_c58_0 = p_29_58 << 1;
  assign t_r30_c58_1 = p_30_57 << 1;
  assign t_r30_c58_2 = p_30_58 << 2;
  assign t_r30_c58_3 = p_30_59 << 1;
  assign t_r30_c58_4 = p_31_58 << 1;
  assign t_r30_c58_5 = t_r30_c58_0 + p_29_57;
  assign t_r30_c58_6 = t_r30_c58_1 + p_29_59;
  assign t_r30_c58_7 = t_r30_c58_2 + t_r30_c58_3;
  assign t_r30_c58_8 = t_r30_c58_4 + p_31_57;
  assign t_r30_c58_9 = t_r30_c58_5 + t_r30_c58_6;
  assign t_r30_c58_10 = t_r30_c58_7 + t_r30_c58_8;
  assign t_r30_c58_11 = t_r30_c58_9 + t_r30_c58_10;
  assign t_r30_c58_12 = t_r30_c58_11 + p_31_59;
  assign out_30_58 = t_r30_c58_12 >> 4;

  assign t_r30_c59_0 = p_29_59 << 1;
  assign t_r30_c59_1 = p_30_58 << 1;
  assign t_r30_c59_2 = p_30_59 << 2;
  assign t_r30_c59_3 = p_30_60 << 1;
  assign t_r30_c59_4 = p_31_59 << 1;
  assign t_r30_c59_5 = t_r30_c59_0 + p_29_58;
  assign t_r30_c59_6 = t_r30_c59_1 + p_29_60;
  assign t_r30_c59_7 = t_r30_c59_2 + t_r30_c59_3;
  assign t_r30_c59_8 = t_r30_c59_4 + p_31_58;
  assign t_r30_c59_9 = t_r30_c59_5 + t_r30_c59_6;
  assign t_r30_c59_10 = t_r30_c59_7 + t_r30_c59_8;
  assign t_r30_c59_11 = t_r30_c59_9 + t_r30_c59_10;
  assign t_r30_c59_12 = t_r30_c59_11 + p_31_60;
  assign out_30_59 = t_r30_c59_12 >> 4;

  assign t_r30_c60_0 = p_29_60 << 1;
  assign t_r30_c60_1 = p_30_59 << 1;
  assign t_r30_c60_2 = p_30_60 << 2;
  assign t_r30_c60_3 = p_30_61 << 1;
  assign t_r30_c60_4 = p_31_60 << 1;
  assign t_r30_c60_5 = t_r30_c60_0 + p_29_59;
  assign t_r30_c60_6 = t_r30_c60_1 + p_29_61;
  assign t_r30_c60_7 = t_r30_c60_2 + t_r30_c60_3;
  assign t_r30_c60_8 = t_r30_c60_4 + p_31_59;
  assign t_r30_c60_9 = t_r30_c60_5 + t_r30_c60_6;
  assign t_r30_c60_10 = t_r30_c60_7 + t_r30_c60_8;
  assign t_r30_c60_11 = t_r30_c60_9 + t_r30_c60_10;
  assign t_r30_c60_12 = t_r30_c60_11 + p_31_61;
  assign out_30_60 = t_r30_c60_12 >> 4;

  assign t_r30_c61_0 = p_29_61 << 1;
  assign t_r30_c61_1 = p_30_60 << 1;
  assign t_r30_c61_2 = p_30_61 << 2;
  assign t_r30_c61_3 = p_30_62 << 1;
  assign t_r30_c61_4 = p_31_61 << 1;
  assign t_r30_c61_5 = t_r30_c61_0 + p_29_60;
  assign t_r30_c61_6 = t_r30_c61_1 + p_29_62;
  assign t_r30_c61_7 = t_r30_c61_2 + t_r30_c61_3;
  assign t_r30_c61_8 = t_r30_c61_4 + p_31_60;
  assign t_r30_c61_9 = t_r30_c61_5 + t_r30_c61_6;
  assign t_r30_c61_10 = t_r30_c61_7 + t_r30_c61_8;
  assign t_r30_c61_11 = t_r30_c61_9 + t_r30_c61_10;
  assign t_r30_c61_12 = t_r30_c61_11 + p_31_62;
  assign out_30_61 = t_r30_c61_12 >> 4;

  assign t_r30_c62_0 = p_29_62 << 1;
  assign t_r30_c62_1 = p_30_61 << 1;
  assign t_r30_c62_2 = p_30_62 << 2;
  assign t_r30_c62_3 = p_30_63 << 1;
  assign t_r30_c62_4 = p_31_62 << 1;
  assign t_r30_c62_5 = t_r30_c62_0 + p_29_61;
  assign t_r30_c62_6 = t_r30_c62_1 + p_29_63;
  assign t_r30_c62_7 = t_r30_c62_2 + t_r30_c62_3;
  assign t_r30_c62_8 = t_r30_c62_4 + p_31_61;
  assign t_r30_c62_9 = t_r30_c62_5 + t_r30_c62_6;
  assign t_r30_c62_10 = t_r30_c62_7 + t_r30_c62_8;
  assign t_r30_c62_11 = t_r30_c62_9 + t_r30_c62_10;
  assign t_r30_c62_12 = t_r30_c62_11 + p_31_63;
  assign out_30_62 = t_r30_c62_12 >> 4;

  assign t_r30_c63_0 = p_29_63 << 1;
  assign t_r30_c63_1 = p_30_62 << 1;
  assign t_r30_c63_2 = p_30_63 << 2;
  assign t_r30_c63_3 = p_30_64 << 1;
  assign t_r30_c63_4 = p_31_63 << 1;
  assign t_r30_c63_5 = t_r30_c63_0 + p_29_62;
  assign t_r30_c63_6 = t_r30_c63_1 + p_29_64;
  assign t_r30_c63_7 = t_r30_c63_2 + t_r30_c63_3;
  assign t_r30_c63_8 = t_r30_c63_4 + p_31_62;
  assign t_r30_c63_9 = t_r30_c63_5 + t_r30_c63_6;
  assign t_r30_c63_10 = t_r30_c63_7 + t_r30_c63_8;
  assign t_r30_c63_11 = t_r30_c63_9 + t_r30_c63_10;
  assign t_r30_c63_12 = t_r30_c63_11 + p_31_64;
  assign out_30_63 = t_r30_c63_12 >> 4;

  assign t_r30_c64_0 = p_29_64 << 1;
  assign t_r30_c64_1 = p_30_63 << 1;
  assign t_r30_c64_2 = p_30_64 << 2;
  assign t_r30_c64_3 = p_30_65 << 1;
  assign t_r30_c64_4 = p_31_64 << 1;
  assign t_r30_c64_5 = t_r30_c64_0 + p_29_63;
  assign t_r30_c64_6 = t_r30_c64_1 + p_29_65;
  assign t_r30_c64_7 = t_r30_c64_2 + t_r30_c64_3;
  assign t_r30_c64_8 = t_r30_c64_4 + p_31_63;
  assign t_r30_c64_9 = t_r30_c64_5 + t_r30_c64_6;
  assign t_r30_c64_10 = t_r30_c64_7 + t_r30_c64_8;
  assign t_r30_c64_11 = t_r30_c64_9 + t_r30_c64_10;
  assign t_r30_c64_12 = t_r30_c64_11 + p_31_65;
  assign out_30_64 = t_r30_c64_12 >> 4;

  assign t_r31_c1_0 = p_30_1 << 1;
  assign t_r31_c1_1 = p_31_0 << 1;
  assign t_r31_c1_2 = p_31_1 << 2;
  assign t_r31_c1_3 = p_31_2 << 1;
  assign t_r31_c1_4 = p_32_1 << 1;
  assign t_r31_c1_5 = t_r31_c1_0 + p_30_0;
  assign t_r31_c1_6 = t_r31_c1_1 + p_30_2;
  assign t_r31_c1_7 = t_r31_c1_2 + t_r31_c1_3;
  assign t_r31_c1_8 = t_r31_c1_4 + p_32_0;
  assign t_r31_c1_9 = t_r31_c1_5 + t_r31_c1_6;
  assign t_r31_c1_10 = t_r31_c1_7 + t_r31_c1_8;
  assign t_r31_c1_11 = t_r31_c1_9 + t_r31_c1_10;
  assign t_r31_c1_12 = t_r31_c1_11 + p_32_2;
  assign out_31_1 = t_r31_c1_12 >> 4;

  assign t_r31_c2_0 = p_30_2 << 1;
  assign t_r31_c2_1 = p_31_1 << 1;
  assign t_r31_c2_2 = p_31_2 << 2;
  assign t_r31_c2_3 = p_31_3 << 1;
  assign t_r31_c2_4 = p_32_2 << 1;
  assign t_r31_c2_5 = t_r31_c2_0 + p_30_1;
  assign t_r31_c2_6 = t_r31_c2_1 + p_30_3;
  assign t_r31_c2_7 = t_r31_c2_2 + t_r31_c2_3;
  assign t_r31_c2_8 = t_r31_c2_4 + p_32_1;
  assign t_r31_c2_9 = t_r31_c2_5 + t_r31_c2_6;
  assign t_r31_c2_10 = t_r31_c2_7 + t_r31_c2_8;
  assign t_r31_c2_11 = t_r31_c2_9 + t_r31_c2_10;
  assign t_r31_c2_12 = t_r31_c2_11 + p_32_3;
  assign out_31_2 = t_r31_c2_12 >> 4;

  assign t_r31_c3_0 = p_30_3 << 1;
  assign t_r31_c3_1 = p_31_2 << 1;
  assign t_r31_c3_2 = p_31_3 << 2;
  assign t_r31_c3_3 = p_31_4 << 1;
  assign t_r31_c3_4 = p_32_3 << 1;
  assign t_r31_c3_5 = t_r31_c3_0 + p_30_2;
  assign t_r31_c3_6 = t_r31_c3_1 + p_30_4;
  assign t_r31_c3_7 = t_r31_c3_2 + t_r31_c3_3;
  assign t_r31_c3_8 = t_r31_c3_4 + p_32_2;
  assign t_r31_c3_9 = t_r31_c3_5 + t_r31_c3_6;
  assign t_r31_c3_10 = t_r31_c3_7 + t_r31_c3_8;
  assign t_r31_c3_11 = t_r31_c3_9 + t_r31_c3_10;
  assign t_r31_c3_12 = t_r31_c3_11 + p_32_4;
  assign out_31_3 = t_r31_c3_12 >> 4;

  assign t_r31_c4_0 = p_30_4 << 1;
  assign t_r31_c4_1 = p_31_3 << 1;
  assign t_r31_c4_2 = p_31_4 << 2;
  assign t_r31_c4_3 = p_31_5 << 1;
  assign t_r31_c4_4 = p_32_4 << 1;
  assign t_r31_c4_5 = t_r31_c4_0 + p_30_3;
  assign t_r31_c4_6 = t_r31_c4_1 + p_30_5;
  assign t_r31_c4_7 = t_r31_c4_2 + t_r31_c4_3;
  assign t_r31_c4_8 = t_r31_c4_4 + p_32_3;
  assign t_r31_c4_9 = t_r31_c4_5 + t_r31_c4_6;
  assign t_r31_c4_10 = t_r31_c4_7 + t_r31_c4_8;
  assign t_r31_c4_11 = t_r31_c4_9 + t_r31_c4_10;
  assign t_r31_c4_12 = t_r31_c4_11 + p_32_5;
  assign out_31_4 = t_r31_c4_12 >> 4;

  assign t_r31_c5_0 = p_30_5 << 1;
  assign t_r31_c5_1 = p_31_4 << 1;
  assign t_r31_c5_2 = p_31_5 << 2;
  assign t_r31_c5_3 = p_31_6 << 1;
  assign t_r31_c5_4 = p_32_5 << 1;
  assign t_r31_c5_5 = t_r31_c5_0 + p_30_4;
  assign t_r31_c5_6 = t_r31_c5_1 + p_30_6;
  assign t_r31_c5_7 = t_r31_c5_2 + t_r31_c5_3;
  assign t_r31_c5_8 = t_r31_c5_4 + p_32_4;
  assign t_r31_c5_9 = t_r31_c5_5 + t_r31_c5_6;
  assign t_r31_c5_10 = t_r31_c5_7 + t_r31_c5_8;
  assign t_r31_c5_11 = t_r31_c5_9 + t_r31_c5_10;
  assign t_r31_c5_12 = t_r31_c5_11 + p_32_6;
  assign out_31_5 = t_r31_c5_12 >> 4;

  assign t_r31_c6_0 = p_30_6 << 1;
  assign t_r31_c6_1 = p_31_5 << 1;
  assign t_r31_c6_2 = p_31_6 << 2;
  assign t_r31_c6_3 = p_31_7 << 1;
  assign t_r31_c6_4 = p_32_6 << 1;
  assign t_r31_c6_5 = t_r31_c6_0 + p_30_5;
  assign t_r31_c6_6 = t_r31_c6_1 + p_30_7;
  assign t_r31_c6_7 = t_r31_c6_2 + t_r31_c6_3;
  assign t_r31_c6_8 = t_r31_c6_4 + p_32_5;
  assign t_r31_c6_9 = t_r31_c6_5 + t_r31_c6_6;
  assign t_r31_c6_10 = t_r31_c6_7 + t_r31_c6_8;
  assign t_r31_c6_11 = t_r31_c6_9 + t_r31_c6_10;
  assign t_r31_c6_12 = t_r31_c6_11 + p_32_7;
  assign out_31_6 = t_r31_c6_12 >> 4;

  assign t_r31_c7_0 = p_30_7 << 1;
  assign t_r31_c7_1 = p_31_6 << 1;
  assign t_r31_c7_2 = p_31_7 << 2;
  assign t_r31_c7_3 = p_31_8 << 1;
  assign t_r31_c7_4 = p_32_7 << 1;
  assign t_r31_c7_5 = t_r31_c7_0 + p_30_6;
  assign t_r31_c7_6 = t_r31_c7_1 + p_30_8;
  assign t_r31_c7_7 = t_r31_c7_2 + t_r31_c7_3;
  assign t_r31_c7_8 = t_r31_c7_4 + p_32_6;
  assign t_r31_c7_9 = t_r31_c7_5 + t_r31_c7_6;
  assign t_r31_c7_10 = t_r31_c7_7 + t_r31_c7_8;
  assign t_r31_c7_11 = t_r31_c7_9 + t_r31_c7_10;
  assign t_r31_c7_12 = t_r31_c7_11 + p_32_8;
  assign out_31_7 = t_r31_c7_12 >> 4;

  assign t_r31_c8_0 = p_30_8 << 1;
  assign t_r31_c8_1 = p_31_7 << 1;
  assign t_r31_c8_2 = p_31_8 << 2;
  assign t_r31_c8_3 = p_31_9 << 1;
  assign t_r31_c8_4 = p_32_8 << 1;
  assign t_r31_c8_5 = t_r31_c8_0 + p_30_7;
  assign t_r31_c8_6 = t_r31_c8_1 + p_30_9;
  assign t_r31_c8_7 = t_r31_c8_2 + t_r31_c8_3;
  assign t_r31_c8_8 = t_r31_c8_4 + p_32_7;
  assign t_r31_c8_9 = t_r31_c8_5 + t_r31_c8_6;
  assign t_r31_c8_10 = t_r31_c8_7 + t_r31_c8_8;
  assign t_r31_c8_11 = t_r31_c8_9 + t_r31_c8_10;
  assign t_r31_c8_12 = t_r31_c8_11 + p_32_9;
  assign out_31_8 = t_r31_c8_12 >> 4;

  assign t_r31_c9_0 = p_30_9 << 1;
  assign t_r31_c9_1 = p_31_8 << 1;
  assign t_r31_c9_2 = p_31_9 << 2;
  assign t_r31_c9_3 = p_31_10 << 1;
  assign t_r31_c9_4 = p_32_9 << 1;
  assign t_r31_c9_5 = t_r31_c9_0 + p_30_8;
  assign t_r31_c9_6 = t_r31_c9_1 + p_30_10;
  assign t_r31_c9_7 = t_r31_c9_2 + t_r31_c9_3;
  assign t_r31_c9_8 = t_r31_c9_4 + p_32_8;
  assign t_r31_c9_9 = t_r31_c9_5 + t_r31_c9_6;
  assign t_r31_c9_10 = t_r31_c9_7 + t_r31_c9_8;
  assign t_r31_c9_11 = t_r31_c9_9 + t_r31_c9_10;
  assign t_r31_c9_12 = t_r31_c9_11 + p_32_10;
  assign out_31_9 = t_r31_c9_12 >> 4;

  assign t_r31_c10_0 = p_30_10 << 1;
  assign t_r31_c10_1 = p_31_9 << 1;
  assign t_r31_c10_2 = p_31_10 << 2;
  assign t_r31_c10_3 = p_31_11 << 1;
  assign t_r31_c10_4 = p_32_10 << 1;
  assign t_r31_c10_5 = t_r31_c10_0 + p_30_9;
  assign t_r31_c10_6 = t_r31_c10_1 + p_30_11;
  assign t_r31_c10_7 = t_r31_c10_2 + t_r31_c10_3;
  assign t_r31_c10_8 = t_r31_c10_4 + p_32_9;
  assign t_r31_c10_9 = t_r31_c10_5 + t_r31_c10_6;
  assign t_r31_c10_10 = t_r31_c10_7 + t_r31_c10_8;
  assign t_r31_c10_11 = t_r31_c10_9 + t_r31_c10_10;
  assign t_r31_c10_12 = t_r31_c10_11 + p_32_11;
  assign out_31_10 = t_r31_c10_12 >> 4;

  assign t_r31_c11_0 = p_30_11 << 1;
  assign t_r31_c11_1 = p_31_10 << 1;
  assign t_r31_c11_2 = p_31_11 << 2;
  assign t_r31_c11_3 = p_31_12 << 1;
  assign t_r31_c11_4 = p_32_11 << 1;
  assign t_r31_c11_5 = t_r31_c11_0 + p_30_10;
  assign t_r31_c11_6 = t_r31_c11_1 + p_30_12;
  assign t_r31_c11_7 = t_r31_c11_2 + t_r31_c11_3;
  assign t_r31_c11_8 = t_r31_c11_4 + p_32_10;
  assign t_r31_c11_9 = t_r31_c11_5 + t_r31_c11_6;
  assign t_r31_c11_10 = t_r31_c11_7 + t_r31_c11_8;
  assign t_r31_c11_11 = t_r31_c11_9 + t_r31_c11_10;
  assign t_r31_c11_12 = t_r31_c11_11 + p_32_12;
  assign out_31_11 = t_r31_c11_12 >> 4;

  assign t_r31_c12_0 = p_30_12 << 1;
  assign t_r31_c12_1 = p_31_11 << 1;
  assign t_r31_c12_2 = p_31_12 << 2;
  assign t_r31_c12_3 = p_31_13 << 1;
  assign t_r31_c12_4 = p_32_12 << 1;
  assign t_r31_c12_5 = t_r31_c12_0 + p_30_11;
  assign t_r31_c12_6 = t_r31_c12_1 + p_30_13;
  assign t_r31_c12_7 = t_r31_c12_2 + t_r31_c12_3;
  assign t_r31_c12_8 = t_r31_c12_4 + p_32_11;
  assign t_r31_c12_9 = t_r31_c12_5 + t_r31_c12_6;
  assign t_r31_c12_10 = t_r31_c12_7 + t_r31_c12_8;
  assign t_r31_c12_11 = t_r31_c12_9 + t_r31_c12_10;
  assign t_r31_c12_12 = t_r31_c12_11 + p_32_13;
  assign out_31_12 = t_r31_c12_12 >> 4;

  assign t_r31_c13_0 = p_30_13 << 1;
  assign t_r31_c13_1 = p_31_12 << 1;
  assign t_r31_c13_2 = p_31_13 << 2;
  assign t_r31_c13_3 = p_31_14 << 1;
  assign t_r31_c13_4 = p_32_13 << 1;
  assign t_r31_c13_5 = t_r31_c13_0 + p_30_12;
  assign t_r31_c13_6 = t_r31_c13_1 + p_30_14;
  assign t_r31_c13_7 = t_r31_c13_2 + t_r31_c13_3;
  assign t_r31_c13_8 = t_r31_c13_4 + p_32_12;
  assign t_r31_c13_9 = t_r31_c13_5 + t_r31_c13_6;
  assign t_r31_c13_10 = t_r31_c13_7 + t_r31_c13_8;
  assign t_r31_c13_11 = t_r31_c13_9 + t_r31_c13_10;
  assign t_r31_c13_12 = t_r31_c13_11 + p_32_14;
  assign out_31_13 = t_r31_c13_12 >> 4;

  assign t_r31_c14_0 = p_30_14 << 1;
  assign t_r31_c14_1 = p_31_13 << 1;
  assign t_r31_c14_2 = p_31_14 << 2;
  assign t_r31_c14_3 = p_31_15 << 1;
  assign t_r31_c14_4 = p_32_14 << 1;
  assign t_r31_c14_5 = t_r31_c14_0 + p_30_13;
  assign t_r31_c14_6 = t_r31_c14_1 + p_30_15;
  assign t_r31_c14_7 = t_r31_c14_2 + t_r31_c14_3;
  assign t_r31_c14_8 = t_r31_c14_4 + p_32_13;
  assign t_r31_c14_9 = t_r31_c14_5 + t_r31_c14_6;
  assign t_r31_c14_10 = t_r31_c14_7 + t_r31_c14_8;
  assign t_r31_c14_11 = t_r31_c14_9 + t_r31_c14_10;
  assign t_r31_c14_12 = t_r31_c14_11 + p_32_15;
  assign out_31_14 = t_r31_c14_12 >> 4;

  assign t_r31_c15_0 = p_30_15 << 1;
  assign t_r31_c15_1 = p_31_14 << 1;
  assign t_r31_c15_2 = p_31_15 << 2;
  assign t_r31_c15_3 = p_31_16 << 1;
  assign t_r31_c15_4 = p_32_15 << 1;
  assign t_r31_c15_5 = t_r31_c15_0 + p_30_14;
  assign t_r31_c15_6 = t_r31_c15_1 + p_30_16;
  assign t_r31_c15_7 = t_r31_c15_2 + t_r31_c15_3;
  assign t_r31_c15_8 = t_r31_c15_4 + p_32_14;
  assign t_r31_c15_9 = t_r31_c15_5 + t_r31_c15_6;
  assign t_r31_c15_10 = t_r31_c15_7 + t_r31_c15_8;
  assign t_r31_c15_11 = t_r31_c15_9 + t_r31_c15_10;
  assign t_r31_c15_12 = t_r31_c15_11 + p_32_16;
  assign out_31_15 = t_r31_c15_12 >> 4;

  assign t_r31_c16_0 = p_30_16 << 1;
  assign t_r31_c16_1 = p_31_15 << 1;
  assign t_r31_c16_2 = p_31_16 << 2;
  assign t_r31_c16_3 = p_31_17 << 1;
  assign t_r31_c16_4 = p_32_16 << 1;
  assign t_r31_c16_5 = t_r31_c16_0 + p_30_15;
  assign t_r31_c16_6 = t_r31_c16_1 + p_30_17;
  assign t_r31_c16_7 = t_r31_c16_2 + t_r31_c16_3;
  assign t_r31_c16_8 = t_r31_c16_4 + p_32_15;
  assign t_r31_c16_9 = t_r31_c16_5 + t_r31_c16_6;
  assign t_r31_c16_10 = t_r31_c16_7 + t_r31_c16_8;
  assign t_r31_c16_11 = t_r31_c16_9 + t_r31_c16_10;
  assign t_r31_c16_12 = t_r31_c16_11 + p_32_17;
  assign out_31_16 = t_r31_c16_12 >> 4;

  assign t_r31_c17_0 = p_30_17 << 1;
  assign t_r31_c17_1 = p_31_16 << 1;
  assign t_r31_c17_2 = p_31_17 << 2;
  assign t_r31_c17_3 = p_31_18 << 1;
  assign t_r31_c17_4 = p_32_17 << 1;
  assign t_r31_c17_5 = t_r31_c17_0 + p_30_16;
  assign t_r31_c17_6 = t_r31_c17_1 + p_30_18;
  assign t_r31_c17_7 = t_r31_c17_2 + t_r31_c17_3;
  assign t_r31_c17_8 = t_r31_c17_4 + p_32_16;
  assign t_r31_c17_9 = t_r31_c17_5 + t_r31_c17_6;
  assign t_r31_c17_10 = t_r31_c17_7 + t_r31_c17_8;
  assign t_r31_c17_11 = t_r31_c17_9 + t_r31_c17_10;
  assign t_r31_c17_12 = t_r31_c17_11 + p_32_18;
  assign out_31_17 = t_r31_c17_12 >> 4;

  assign t_r31_c18_0 = p_30_18 << 1;
  assign t_r31_c18_1 = p_31_17 << 1;
  assign t_r31_c18_2 = p_31_18 << 2;
  assign t_r31_c18_3 = p_31_19 << 1;
  assign t_r31_c18_4 = p_32_18 << 1;
  assign t_r31_c18_5 = t_r31_c18_0 + p_30_17;
  assign t_r31_c18_6 = t_r31_c18_1 + p_30_19;
  assign t_r31_c18_7 = t_r31_c18_2 + t_r31_c18_3;
  assign t_r31_c18_8 = t_r31_c18_4 + p_32_17;
  assign t_r31_c18_9 = t_r31_c18_5 + t_r31_c18_6;
  assign t_r31_c18_10 = t_r31_c18_7 + t_r31_c18_8;
  assign t_r31_c18_11 = t_r31_c18_9 + t_r31_c18_10;
  assign t_r31_c18_12 = t_r31_c18_11 + p_32_19;
  assign out_31_18 = t_r31_c18_12 >> 4;

  assign t_r31_c19_0 = p_30_19 << 1;
  assign t_r31_c19_1 = p_31_18 << 1;
  assign t_r31_c19_2 = p_31_19 << 2;
  assign t_r31_c19_3 = p_31_20 << 1;
  assign t_r31_c19_4 = p_32_19 << 1;
  assign t_r31_c19_5 = t_r31_c19_0 + p_30_18;
  assign t_r31_c19_6 = t_r31_c19_1 + p_30_20;
  assign t_r31_c19_7 = t_r31_c19_2 + t_r31_c19_3;
  assign t_r31_c19_8 = t_r31_c19_4 + p_32_18;
  assign t_r31_c19_9 = t_r31_c19_5 + t_r31_c19_6;
  assign t_r31_c19_10 = t_r31_c19_7 + t_r31_c19_8;
  assign t_r31_c19_11 = t_r31_c19_9 + t_r31_c19_10;
  assign t_r31_c19_12 = t_r31_c19_11 + p_32_20;
  assign out_31_19 = t_r31_c19_12 >> 4;

  assign t_r31_c20_0 = p_30_20 << 1;
  assign t_r31_c20_1 = p_31_19 << 1;
  assign t_r31_c20_2 = p_31_20 << 2;
  assign t_r31_c20_3 = p_31_21 << 1;
  assign t_r31_c20_4 = p_32_20 << 1;
  assign t_r31_c20_5 = t_r31_c20_0 + p_30_19;
  assign t_r31_c20_6 = t_r31_c20_1 + p_30_21;
  assign t_r31_c20_7 = t_r31_c20_2 + t_r31_c20_3;
  assign t_r31_c20_8 = t_r31_c20_4 + p_32_19;
  assign t_r31_c20_9 = t_r31_c20_5 + t_r31_c20_6;
  assign t_r31_c20_10 = t_r31_c20_7 + t_r31_c20_8;
  assign t_r31_c20_11 = t_r31_c20_9 + t_r31_c20_10;
  assign t_r31_c20_12 = t_r31_c20_11 + p_32_21;
  assign out_31_20 = t_r31_c20_12 >> 4;

  assign t_r31_c21_0 = p_30_21 << 1;
  assign t_r31_c21_1 = p_31_20 << 1;
  assign t_r31_c21_2 = p_31_21 << 2;
  assign t_r31_c21_3 = p_31_22 << 1;
  assign t_r31_c21_4 = p_32_21 << 1;
  assign t_r31_c21_5 = t_r31_c21_0 + p_30_20;
  assign t_r31_c21_6 = t_r31_c21_1 + p_30_22;
  assign t_r31_c21_7 = t_r31_c21_2 + t_r31_c21_3;
  assign t_r31_c21_8 = t_r31_c21_4 + p_32_20;
  assign t_r31_c21_9 = t_r31_c21_5 + t_r31_c21_6;
  assign t_r31_c21_10 = t_r31_c21_7 + t_r31_c21_8;
  assign t_r31_c21_11 = t_r31_c21_9 + t_r31_c21_10;
  assign t_r31_c21_12 = t_r31_c21_11 + p_32_22;
  assign out_31_21 = t_r31_c21_12 >> 4;

  assign t_r31_c22_0 = p_30_22 << 1;
  assign t_r31_c22_1 = p_31_21 << 1;
  assign t_r31_c22_2 = p_31_22 << 2;
  assign t_r31_c22_3 = p_31_23 << 1;
  assign t_r31_c22_4 = p_32_22 << 1;
  assign t_r31_c22_5 = t_r31_c22_0 + p_30_21;
  assign t_r31_c22_6 = t_r31_c22_1 + p_30_23;
  assign t_r31_c22_7 = t_r31_c22_2 + t_r31_c22_3;
  assign t_r31_c22_8 = t_r31_c22_4 + p_32_21;
  assign t_r31_c22_9 = t_r31_c22_5 + t_r31_c22_6;
  assign t_r31_c22_10 = t_r31_c22_7 + t_r31_c22_8;
  assign t_r31_c22_11 = t_r31_c22_9 + t_r31_c22_10;
  assign t_r31_c22_12 = t_r31_c22_11 + p_32_23;
  assign out_31_22 = t_r31_c22_12 >> 4;

  assign t_r31_c23_0 = p_30_23 << 1;
  assign t_r31_c23_1 = p_31_22 << 1;
  assign t_r31_c23_2 = p_31_23 << 2;
  assign t_r31_c23_3 = p_31_24 << 1;
  assign t_r31_c23_4 = p_32_23 << 1;
  assign t_r31_c23_5 = t_r31_c23_0 + p_30_22;
  assign t_r31_c23_6 = t_r31_c23_1 + p_30_24;
  assign t_r31_c23_7 = t_r31_c23_2 + t_r31_c23_3;
  assign t_r31_c23_8 = t_r31_c23_4 + p_32_22;
  assign t_r31_c23_9 = t_r31_c23_5 + t_r31_c23_6;
  assign t_r31_c23_10 = t_r31_c23_7 + t_r31_c23_8;
  assign t_r31_c23_11 = t_r31_c23_9 + t_r31_c23_10;
  assign t_r31_c23_12 = t_r31_c23_11 + p_32_24;
  assign out_31_23 = t_r31_c23_12 >> 4;

  assign t_r31_c24_0 = p_30_24 << 1;
  assign t_r31_c24_1 = p_31_23 << 1;
  assign t_r31_c24_2 = p_31_24 << 2;
  assign t_r31_c24_3 = p_31_25 << 1;
  assign t_r31_c24_4 = p_32_24 << 1;
  assign t_r31_c24_5 = t_r31_c24_0 + p_30_23;
  assign t_r31_c24_6 = t_r31_c24_1 + p_30_25;
  assign t_r31_c24_7 = t_r31_c24_2 + t_r31_c24_3;
  assign t_r31_c24_8 = t_r31_c24_4 + p_32_23;
  assign t_r31_c24_9 = t_r31_c24_5 + t_r31_c24_6;
  assign t_r31_c24_10 = t_r31_c24_7 + t_r31_c24_8;
  assign t_r31_c24_11 = t_r31_c24_9 + t_r31_c24_10;
  assign t_r31_c24_12 = t_r31_c24_11 + p_32_25;
  assign out_31_24 = t_r31_c24_12 >> 4;

  assign t_r31_c25_0 = p_30_25 << 1;
  assign t_r31_c25_1 = p_31_24 << 1;
  assign t_r31_c25_2 = p_31_25 << 2;
  assign t_r31_c25_3 = p_31_26 << 1;
  assign t_r31_c25_4 = p_32_25 << 1;
  assign t_r31_c25_5 = t_r31_c25_0 + p_30_24;
  assign t_r31_c25_6 = t_r31_c25_1 + p_30_26;
  assign t_r31_c25_7 = t_r31_c25_2 + t_r31_c25_3;
  assign t_r31_c25_8 = t_r31_c25_4 + p_32_24;
  assign t_r31_c25_9 = t_r31_c25_5 + t_r31_c25_6;
  assign t_r31_c25_10 = t_r31_c25_7 + t_r31_c25_8;
  assign t_r31_c25_11 = t_r31_c25_9 + t_r31_c25_10;
  assign t_r31_c25_12 = t_r31_c25_11 + p_32_26;
  assign out_31_25 = t_r31_c25_12 >> 4;

  assign t_r31_c26_0 = p_30_26 << 1;
  assign t_r31_c26_1 = p_31_25 << 1;
  assign t_r31_c26_2 = p_31_26 << 2;
  assign t_r31_c26_3 = p_31_27 << 1;
  assign t_r31_c26_4 = p_32_26 << 1;
  assign t_r31_c26_5 = t_r31_c26_0 + p_30_25;
  assign t_r31_c26_6 = t_r31_c26_1 + p_30_27;
  assign t_r31_c26_7 = t_r31_c26_2 + t_r31_c26_3;
  assign t_r31_c26_8 = t_r31_c26_4 + p_32_25;
  assign t_r31_c26_9 = t_r31_c26_5 + t_r31_c26_6;
  assign t_r31_c26_10 = t_r31_c26_7 + t_r31_c26_8;
  assign t_r31_c26_11 = t_r31_c26_9 + t_r31_c26_10;
  assign t_r31_c26_12 = t_r31_c26_11 + p_32_27;
  assign out_31_26 = t_r31_c26_12 >> 4;

  assign t_r31_c27_0 = p_30_27 << 1;
  assign t_r31_c27_1 = p_31_26 << 1;
  assign t_r31_c27_2 = p_31_27 << 2;
  assign t_r31_c27_3 = p_31_28 << 1;
  assign t_r31_c27_4 = p_32_27 << 1;
  assign t_r31_c27_5 = t_r31_c27_0 + p_30_26;
  assign t_r31_c27_6 = t_r31_c27_1 + p_30_28;
  assign t_r31_c27_7 = t_r31_c27_2 + t_r31_c27_3;
  assign t_r31_c27_8 = t_r31_c27_4 + p_32_26;
  assign t_r31_c27_9 = t_r31_c27_5 + t_r31_c27_6;
  assign t_r31_c27_10 = t_r31_c27_7 + t_r31_c27_8;
  assign t_r31_c27_11 = t_r31_c27_9 + t_r31_c27_10;
  assign t_r31_c27_12 = t_r31_c27_11 + p_32_28;
  assign out_31_27 = t_r31_c27_12 >> 4;

  assign t_r31_c28_0 = p_30_28 << 1;
  assign t_r31_c28_1 = p_31_27 << 1;
  assign t_r31_c28_2 = p_31_28 << 2;
  assign t_r31_c28_3 = p_31_29 << 1;
  assign t_r31_c28_4 = p_32_28 << 1;
  assign t_r31_c28_5 = t_r31_c28_0 + p_30_27;
  assign t_r31_c28_6 = t_r31_c28_1 + p_30_29;
  assign t_r31_c28_7 = t_r31_c28_2 + t_r31_c28_3;
  assign t_r31_c28_8 = t_r31_c28_4 + p_32_27;
  assign t_r31_c28_9 = t_r31_c28_5 + t_r31_c28_6;
  assign t_r31_c28_10 = t_r31_c28_7 + t_r31_c28_8;
  assign t_r31_c28_11 = t_r31_c28_9 + t_r31_c28_10;
  assign t_r31_c28_12 = t_r31_c28_11 + p_32_29;
  assign out_31_28 = t_r31_c28_12 >> 4;

  assign t_r31_c29_0 = p_30_29 << 1;
  assign t_r31_c29_1 = p_31_28 << 1;
  assign t_r31_c29_2 = p_31_29 << 2;
  assign t_r31_c29_3 = p_31_30 << 1;
  assign t_r31_c29_4 = p_32_29 << 1;
  assign t_r31_c29_5 = t_r31_c29_0 + p_30_28;
  assign t_r31_c29_6 = t_r31_c29_1 + p_30_30;
  assign t_r31_c29_7 = t_r31_c29_2 + t_r31_c29_3;
  assign t_r31_c29_8 = t_r31_c29_4 + p_32_28;
  assign t_r31_c29_9 = t_r31_c29_5 + t_r31_c29_6;
  assign t_r31_c29_10 = t_r31_c29_7 + t_r31_c29_8;
  assign t_r31_c29_11 = t_r31_c29_9 + t_r31_c29_10;
  assign t_r31_c29_12 = t_r31_c29_11 + p_32_30;
  assign out_31_29 = t_r31_c29_12 >> 4;

  assign t_r31_c30_0 = p_30_30 << 1;
  assign t_r31_c30_1 = p_31_29 << 1;
  assign t_r31_c30_2 = p_31_30 << 2;
  assign t_r31_c30_3 = p_31_31 << 1;
  assign t_r31_c30_4 = p_32_30 << 1;
  assign t_r31_c30_5 = t_r31_c30_0 + p_30_29;
  assign t_r31_c30_6 = t_r31_c30_1 + p_30_31;
  assign t_r31_c30_7 = t_r31_c30_2 + t_r31_c30_3;
  assign t_r31_c30_8 = t_r31_c30_4 + p_32_29;
  assign t_r31_c30_9 = t_r31_c30_5 + t_r31_c30_6;
  assign t_r31_c30_10 = t_r31_c30_7 + t_r31_c30_8;
  assign t_r31_c30_11 = t_r31_c30_9 + t_r31_c30_10;
  assign t_r31_c30_12 = t_r31_c30_11 + p_32_31;
  assign out_31_30 = t_r31_c30_12 >> 4;

  assign t_r31_c31_0 = p_30_31 << 1;
  assign t_r31_c31_1 = p_31_30 << 1;
  assign t_r31_c31_2 = p_31_31 << 2;
  assign t_r31_c31_3 = p_31_32 << 1;
  assign t_r31_c31_4 = p_32_31 << 1;
  assign t_r31_c31_5 = t_r31_c31_0 + p_30_30;
  assign t_r31_c31_6 = t_r31_c31_1 + p_30_32;
  assign t_r31_c31_7 = t_r31_c31_2 + t_r31_c31_3;
  assign t_r31_c31_8 = t_r31_c31_4 + p_32_30;
  assign t_r31_c31_9 = t_r31_c31_5 + t_r31_c31_6;
  assign t_r31_c31_10 = t_r31_c31_7 + t_r31_c31_8;
  assign t_r31_c31_11 = t_r31_c31_9 + t_r31_c31_10;
  assign t_r31_c31_12 = t_r31_c31_11 + p_32_32;
  assign out_31_31 = t_r31_c31_12 >> 4;

  assign t_r31_c32_0 = p_30_32 << 1;
  assign t_r31_c32_1 = p_31_31 << 1;
  assign t_r31_c32_2 = p_31_32 << 2;
  assign t_r31_c32_3 = p_31_33 << 1;
  assign t_r31_c32_4 = p_32_32 << 1;
  assign t_r31_c32_5 = t_r31_c32_0 + p_30_31;
  assign t_r31_c32_6 = t_r31_c32_1 + p_30_33;
  assign t_r31_c32_7 = t_r31_c32_2 + t_r31_c32_3;
  assign t_r31_c32_8 = t_r31_c32_4 + p_32_31;
  assign t_r31_c32_9 = t_r31_c32_5 + t_r31_c32_6;
  assign t_r31_c32_10 = t_r31_c32_7 + t_r31_c32_8;
  assign t_r31_c32_11 = t_r31_c32_9 + t_r31_c32_10;
  assign t_r31_c32_12 = t_r31_c32_11 + p_32_33;
  assign out_31_32 = t_r31_c32_12 >> 4;

  assign t_r31_c33_0 = p_30_33 << 1;
  assign t_r31_c33_1 = p_31_32 << 1;
  assign t_r31_c33_2 = p_31_33 << 2;
  assign t_r31_c33_3 = p_31_34 << 1;
  assign t_r31_c33_4 = p_32_33 << 1;
  assign t_r31_c33_5 = t_r31_c33_0 + p_30_32;
  assign t_r31_c33_6 = t_r31_c33_1 + p_30_34;
  assign t_r31_c33_7 = t_r31_c33_2 + t_r31_c33_3;
  assign t_r31_c33_8 = t_r31_c33_4 + p_32_32;
  assign t_r31_c33_9 = t_r31_c33_5 + t_r31_c33_6;
  assign t_r31_c33_10 = t_r31_c33_7 + t_r31_c33_8;
  assign t_r31_c33_11 = t_r31_c33_9 + t_r31_c33_10;
  assign t_r31_c33_12 = t_r31_c33_11 + p_32_34;
  assign out_31_33 = t_r31_c33_12 >> 4;

  assign t_r31_c34_0 = p_30_34 << 1;
  assign t_r31_c34_1 = p_31_33 << 1;
  assign t_r31_c34_2 = p_31_34 << 2;
  assign t_r31_c34_3 = p_31_35 << 1;
  assign t_r31_c34_4 = p_32_34 << 1;
  assign t_r31_c34_5 = t_r31_c34_0 + p_30_33;
  assign t_r31_c34_6 = t_r31_c34_1 + p_30_35;
  assign t_r31_c34_7 = t_r31_c34_2 + t_r31_c34_3;
  assign t_r31_c34_8 = t_r31_c34_4 + p_32_33;
  assign t_r31_c34_9 = t_r31_c34_5 + t_r31_c34_6;
  assign t_r31_c34_10 = t_r31_c34_7 + t_r31_c34_8;
  assign t_r31_c34_11 = t_r31_c34_9 + t_r31_c34_10;
  assign t_r31_c34_12 = t_r31_c34_11 + p_32_35;
  assign out_31_34 = t_r31_c34_12 >> 4;

  assign t_r31_c35_0 = p_30_35 << 1;
  assign t_r31_c35_1 = p_31_34 << 1;
  assign t_r31_c35_2 = p_31_35 << 2;
  assign t_r31_c35_3 = p_31_36 << 1;
  assign t_r31_c35_4 = p_32_35 << 1;
  assign t_r31_c35_5 = t_r31_c35_0 + p_30_34;
  assign t_r31_c35_6 = t_r31_c35_1 + p_30_36;
  assign t_r31_c35_7 = t_r31_c35_2 + t_r31_c35_3;
  assign t_r31_c35_8 = t_r31_c35_4 + p_32_34;
  assign t_r31_c35_9 = t_r31_c35_5 + t_r31_c35_6;
  assign t_r31_c35_10 = t_r31_c35_7 + t_r31_c35_8;
  assign t_r31_c35_11 = t_r31_c35_9 + t_r31_c35_10;
  assign t_r31_c35_12 = t_r31_c35_11 + p_32_36;
  assign out_31_35 = t_r31_c35_12 >> 4;

  assign t_r31_c36_0 = p_30_36 << 1;
  assign t_r31_c36_1 = p_31_35 << 1;
  assign t_r31_c36_2 = p_31_36 << 2;
  assign t_r31_c36_3 = p_31_37 << 1;
  assign t_r31_c36_4 = p_32_36 << 1;
  assign t_r31_c36_5 = t_r31_c36_0 + p_30_35;
  assign t_r31_c36_6 = t_r31_c36_1 + p_30_37;
  assign t_r31_c36_7 = t_r31_c36_2 + t_r31_c36_3;
  assign t_r31_c36_8 = t_r31_c36_4 + p_32_35;
  assign t_r31_c36_9 = t_r31_c36_5 + t_r31_c36_6;
  assign t_r31_c36_10 = t_r31_c36_7 + t_r31_c36_8;
  assign t_r31_c36_11 = t_r31_c36_9 + t_r31_c36_10;
  assign t_r31_c36_12 = t_r31_c36_11 + p_32_37;
  assign out_31_36 = t_r31_c36_12 >> 4;

  assign t_r31_c37_0 = p_30_37 << 1;
  assign t_r31_c37_1 = p_31_36 << 1;
  assign t_r31_c37_2 = p_31_37 << 2;
  assign t_r31_c37_3 = p_31_38 << 1;
  assign t_r31_c37_4 = p_32_37 << 1;
  assign t_r31_c37_5 = t_r31_c37_0 + p_30_36;
  assign t_r31_c37_6 = t_r31_c37_1 + p_30_38;
  assign t_r31_c37_7 = t_r31_c37_2 + t_r31_c37_3;
  assign t_r31_c37_8 = t_r31_c37_4 + p_32_36;
  assign t_r31_c37_9 = t_r31_c37_5 + t_r31_c37_6;
  assign t_r31_c37_10 = t_r31_c37_7 + t_r31_c37_8;
  assign t_r31_c37_11 = t_r31_c37_9 + t_r31_c37_10;
  assign t_r31_c37_12 = t_r31_c37_11 + p_32_38;
  assign out_31_37 = t_r31_c37_12 >> 4;

  assign t_r31_c38_0 = p_30_38 << 1;
  assign t_r31_c38_1 = p_31_37 << 1;
  assign t_r31_c38_2 = p_31_38 << 2;
  assign t_r31_c38_3 = p_31_39 << 1;
  assign t_r31_c38_4 = p_32_38 << 1;
  assign t_r31_c38_5 = t_r31_c38_0 + p_30_37;
  assign t_r31_c38_6 = t_r31_c38_1 + p_30_39;
  assign t_r31_c38_7 = t_r31_c38_2 + t_r31_c38_3;
  assign t_r31_c38_8 = t_r31_c38_4 + p_32_37;
  assign t_r31_c38_9 = t_r31_c38_5 + t_r31_c38_6;
  assign t_r31_c38_10 = t_r31_c38_7 + t_r31_c38_8;
  assign t_r31_c38_11 = t_r31_c38_9 + t_r31_c38_10;
  assign t_r31_c38_12 = t_r31_c38_11 + p_32_39;
  assign out_31_38 = t_r31_c38_12 >> 4;

  assign t_r31_c39_0 = p_30_39 << 1;
  assign t_r31_c39_1 = p_31_38 << 1;
  assign t_r31_c39_2 = p_31_39 << 2;
  assign t_r31_c39_3 = p_31_40 << 1;
  assign t_r31_c39_4 = p_32_39 << 1;
  assign t_r31_c39_5 = t_r31_c39_0 + p_30_38;
  assign t_r31_c39_6 = t_r31_c39_1 + p_30_40;
  assign t_r31_c39_7 = t_r31_c39_2 + t_r31_c39_3;
  assign t_r31_c39_8 = t_r31_c39_4 + p_32_38;
  assign t_r31_c39_9 = t_r31_c39_5 + t_r31_c39_6;
  assign t_r31_c39_10 = t_r31_c39_7 + t_r31_c39_8;
  assign t_r31_c39_11 = t_r31_c39_9 + t_r31_c39_10;
  assign t_r31_c39_12 = t_r31_c39_11 + p_32_40;
  assign out_31_39 = t_r31_c39_12 >> 4;

  assign t_r31_c40_0 = p_30_40 << 1;
  assign t_r31_c40_1 = p_31_39 << 1;
  assign t_r31_c40_2 = p_31_40 << 2;
  assign t_r31_c40_3 = p_31_41 << 1;
  assign t_r31_c40_4 = p_32_40 << 1;
  assign t_r31_c40_5 = t_r31_c40_0 + p_30_39;
  assign t_r31_c40_6 = t_r31_c40_1 + p_30_41;
  assign t_r31_c40_7 = t_r31_c40_2 + t_r31_c40_3;
  assign t_r31_c40_8 = t_r31_c40_4 + p_32_39;
  assign t_r31_c40_9 = t_r31_c40_5 + t_r31_c40_6;
  assign t_r31_c40_10 = t_r31_c40_7 + t_r31_c40_8;
  assign t_r31_c40_11 = t_r31_c40_9 + t_r31_c40_10;
  assign t_r31_c40_12 = t_r31_c40_11 + p_32_41;
  assign out_31_40 = t_r31_c40_12 >> 4;

  assign t_r31_c41_0 = p_30_41 << 1;
  assign t_r31_c41_1 = p_31_40 << 1;
  assign t_r31_c41_2 = p_31_41 << 2;
  assign t_r31_c41_3 = p_31_42 << 1;
  assign t_r31_c41_4 = p_32_41 << 1;
  assign t_r31_c41_5 = t_r31_c41_0 + p_30_40;
  assign t_r31_c41_6 = t_r31_c41_1 + p_30_42;
  assign t_r31_c41_7 = t_r31_c41_2 + t_r31_c41_3;
  assign t_r31_c41_8 = t_r31_c41_4 + p_32_40;
  assign t_r31_c41_9 = t_r31_c41_5 + t_r31_c41_6;
  assign t_r31_c41_10 = t_r31_c41_7 + t_r31_c41_8;
  assign t_r31_c41_11 = t_r31_c41_9 + t_r31_c41_10;
  assign t_r31_c41_12 = t_r31_c41_11 + p_32_42;
  assign out_31_41 = t_r31_c41_12 >> 4;

  assign t_r31_c42_0 = p_30_42 << 1;
  assign t_r31_c42_1 = p_31_41 << 1;
  assign t_r31_c42_2 = p_31_42 << 2;
  assign t_r31_c42_3 = p_31_43 << 1;
  assign t_r31_c42_4 = p_32_42 << 1;
  assign t_r31_c42_5 = t_r31_c42_0 + p_30_41;
  assign t_r31_c42_6 = t_r31_c42_1 + p_30_43;
  assign t_r31_c42_7 = t_r31_c42_2 + t_r31_c42_3;
  assign t_r31_c42_8 = t_r31_c42_4 + p_32_41;
  assign t_r31_c42_9 = t_r31_c42_5 + t_r31_c42_6;
  assign t_r31_c42_10 = t_r31_c42_7 + t_r31_c42_8;
  assign t_r31_c42_11 = t_r31_c42_9 + t_r31_c42_10;
  assign t_r31_c42_12 = t_r31_c42_11 + p_32_43;
  assign out_31_42 = t_r31_c42_12 >> 4;

  assign t_r31_c43_0 = p_30_43 << 1;
  assign t_r31_c43_1 = p_31_42 << 1;
  assign t_r31_c43_2 = p_31_43 << 2;
  assign t_r31_c43_3 = p_31_44 << 1;
  assign t_r31_c43_4 = p_32_43 << 1;
  assign t_r31_c43_5 = t_r31_c43_0 + p_30_42;
  assign t_r31_c43_6 = t_r31_c43_1 + p_30_44;
  assign t_r31_c43_7 = t_r31_c43_2 + t_r31_c43_3;
  assign t_r31_c43_8 = t_r31_c43_4 + p_32_42;
  assign t_r31_c43_9 = t_r31_c43_5 + t_r31_c43_6;
  assign t_r31_c43_10 = t_r31_c43_7 + t_r31_c43_8;
  assign t_r31_c43_11 = t_r31_c43_9 + t_r31_c43_10;
  assign t_r31_c43_12 = t_r31_c43_11 + p_32_44;
  assign out_31_43 = t_r31_c43_12 >> 4;

  assign t_r31_c44_0 = p_30_44 << 1;
  assign t_r31_c44_1 = p_31_43 << 1;
  assign t_r31_c44_2 = p_31_44 << 2;
  assign t_r31_c44_3 = p_31_45 << 1;
  assign t_r31_c44_4 = p_32_44 << 1;
  assign t_r31_c44_5 = t_r31_c44_0 + p_30_43;
  assign t_r31_c44_6 = t_r31_c44_1 + p_30_45;
  assign t_r31_c44_7 = t_r31_c44_2 + t_r31_c44_3;
  assign t_r31_c44_8 = t_r31_c44_4 + p_32_43;
  assign t_r31_c44_9 = t_r31_c44_5 + t_r31_c44_6;
  assign t_r31_c44_10 = t_r31_c44_7 + t_r31_c44_8;
  assign t_r31_c44_11 = t_r31_c44_9 + t_r31_c44_10;
  assign t_r31_c44_12 = t_r31_c44_11 + p_32_45;
  assign out_31_44 = t_r31_c44_12 >> 4;

  assign t_r31_c45_0 = p_30_45 << 1;
  assign t_r31_c45_1 = p_31_44 << 1;
  assign t_r31_c45_2 = p_31_45 << 2;
  assign t_r31_c45_3 = p_31_46 << 1;
  assign t_r31_c45_4 = p_32_45 << 1;
  assign t_r31_c45_5 = t_r31_c45_0 + p_30_44;
  assign t_r31_c45_6 = t_r31_c45_1 + p_30_46;
  assign t_r31_c45_7 = t_r31_c45_2 + t_r31_c45_3;
  assign t_r31_c45_8 = t_r31_c45_4 + p_32_44;
  assign t_r31_c45_9 = t_r31_c45_5 + t_r31_c45_6;
  assign t_r31_c45_10 = t_r31_c45_7 + t_r31_c45_8;
  assign t_r31_c45_11 = t_r31_c45_9 + t_r31_c45_10;
  assign t_r31_c45_12 = t_r31_c45_11 + p_32_46;
  assign out_31_45 = t_r31_c45_12 >> 4;

  assign t_r31_c46_0 = p_30_46 << 1;
  assign t_r31_c46_1 = p_31_45 << 1;
  assign t_r31_c46_2 = p_31_46 << 2;
  assign t_r31_c46_3 = p_31_47 << 1;
  assign t_r31_c46_4 = p_32_46 << 1;
  assign t_r31_c46_5 = t_r31_c46_0 + p_30_45;
  assign t_r31_c46_6 = t_r31_c46_1 + p_30_47;
  assign t_r31_c46_7 = t_r31_c46_2 + t_r31_c46_3;
  assign t_r31_c46_8 = t_r31_c46_4 + p_32_45;
  assign t_r31_c46_9 = t_r31_c46_5 + t_r31_c46_6;
  assign t_r31_c46_10 = t_r31_c46_7 + t_r31_c46_8;
  assign t_r31_c46_11 = t_r31_c46_9 + t_r31_c46_10;
  assign t_r31_c46_12 = t_r31_c46_11 + p_32_47;
  assign out_31_46 = t_r31_c46_12 >> 4;

  assign t_r31_c47_0 = p_30_47 << 1;
  assign t_r31_c47_1 = p_31_46 << 1;
  assign t_r31_c47_2 = p_31_47 << 2;
  assign t_r31_c47_3 = p_31_48 << 1;
  assign t_r31_c47_4 = p_32_47 << 1;
  assign t_r31_c47_5 = t_r31_c47_0 + p_30_46;
  assign t_r31_c47_6 = t_r31_c47_1 + p_30_48;
  assign t_r31_c47_7 = t_r31_c47_2 + t_r31_c47_3;
  assign t_r31_c47_8 = t_r31_c47_4 + p_32_46;
  assign t_r31_c47_9 = t_r31_c47_5 + t_r31_c47_6;
  assign t_r31_c47_10 = t_r31_c47_7 + t_r31_c47_8;
  assign t_r31_c47_11 = t_r31_c47_9 + t_r31_c47_10;
  assign t_r31_c47_12 = t_r31_c47_11 + p_32_48;
  assign out_31_47 = t_r31_c47_12 >> 4;

  assign t_r31_c48_0 = p_30_48 << 1;
  assign t_r31_c48_1 = p_31_47 << 1;
  assign t_r31_c48_2 = p_31_48 << 2;
  assign t_r31_c48_3 = p_31_49 << 1;
  assign t_r31_c48_4 = p_32_48 << 1;
  assign t_r31_c48_5 = t_r31_c48_0 + p_30_47;
  assign t_r31_c48_6 = t_r31_c48_1 + p_30_49;
  assign t_r31_c48_7 = t_r31_c48_2 + t_r31_c48_3;
  assign t_r31_c48_8 = t_r31_c48_4 + p_32_47;
  assign t_r31_c48_9 = t_r31_c48_5 + t_r31_c48_6;
  assign t_r31_c48_10 = t_r31_c48_7 + t_r31_c48_8;
  assign t_r31_c48_11 = t_r31_c48_9 + t_r31_c48_10;
  assign t_r31_c48_12 = t_r31_c48_11 + p_32_49;
  assign out_31_48 = t_r31_c48_12 >> 4;

  assign t_r31_c49_0 = p_30_49 << 1;
  assign t_r31_c49_1 = p_31_48 << 1;
  assign t_r31_c49_2 = p_31_49 << 2;
  assign t_r31_c49_3 = p_31_50 << 1;
  assign t_r31_c49_4 = p_32_49 << 1;
  assign t_r31_c49_5 = t_r31_c49_0 + p_30_48;
  assign t_r31_c49_6 = t_r31_c49_1 + p_30_50;
  assign t_r31_c49_7 = t_r31_c49_2 + t_r31_c49_3;
  assign t_r31_c49_8 = t_r31_c49_4 + p_32_48;
  assign t_r31_c49_9 = t_r31_c49_5 + t_r31_c49_6;
  assign t_r31_c49_10 = t_r31_c49_7 + t_r31_c49_8;
  assign t_r31_c49_11 = t_r31_c49_9 + t_r31_c49_10;
  assign t_r31_c49_12 = t_r31_c49_11 + p_32_50;
  assign out_31_49 = t_r31_c49_12 >> 4;

  assign t_r31_c50_0 = p_30_50 << 1;
  assign t_r31_c50_1 = p_31_49 << 1;
  assign t_r31_c50_2 = p_31_50 << 2;
  assign t_r31_c50_3 = p_31_51 << 1;
  assign t_r31_c50_4 = p_32_50 << 1;
  assign t_r31_c50_5 = t_r31_c50_0 + p_30_49;
  assign t_r31_c50_6 = t_r31_c50_1 + p_30_51;
  assign t_r31_c50_7 = t_r31_c50_2 + t_r31_c50_3;
  assign t_r31_c50_8 = t_r31_c50_4 + p_32_49;
  assign t_r31_c50_9 = t_r31_c50_5 + t_r31_c50_6;
  assign t_r31_c50_10 = t_r31_c50_7 + t_r31_c50_8;
  assign t_r31_c50_11 = t_r31_c50_9 + t_r31_c50_10;
  assign t_r31_c50_12 = t_r31_c50_11 + p_32_51;
  assign out_31_50 = t_r31_c50_12 >> 4;

  assign t_r31_c51_0 = p_30_51 << 1;
  assign t_r31_c51_1 = p_31_50 << 1;
  assign t_r31_c51_2 = p_31_51 << 2;
  assign t_r31_c51_3 = p_31_52 << 1;
  assign t_r31_c51_4 = p_32_51 << 1;
  assign t_r31_c51_5 = t_r31_c51_0 + p_30_50;
  assign t_r31_c51_6 = t_r31_c51_1 + p_30_52;
  assign t_r31_c51_7 = t_r31_c51_2 + t_r31_c51_3;
  assign t_r31_c51_8 = t_r31_c51_4 + p_32_50;
  assign t_r31_c51_9 = t_r31_c51_5 + t_r31_c51_6;
  assign t_r31_c51_10 = t_r31_c51_7 + t_r31_c51_8;
  assign t_r31_c51_11 = t_r31_c51_9 + t_r31_c51_10;
  assign t_r31_c51_12 = t_r31_c51_11 + p_32_52;
  assign out_31_51 = t_r31_c51_12 >> 4;

  assign t_r31_c52_0 = p_30_52 << 1;
  assign t_r31_c52_1 = p_31_51 << 1;
  assign t_r31_c52_2 = p_31_52 << 2;
  assign t_r31_c52_3 = p_31_53 << 1;
  assign t_r31_c52_4 = p_32_52 << 1;
  assign t_r31_c52_5 = t_r31_c52_0 + p_30_51;
  assign t_r31_c52_6 = t_r31_c52_1 + p_30_53;
  assign t_r31_c52_7 = t_r31_c52_2 + t_r31_c52_3;
  assign t_r31_c52_8 = t_r31_c52_4 + p_32_51;
  assign t_r31_c52_9 = t_r31_c52_5 + t_r31_c52_6;
  assign t_r31_c52_10 = t_r31_c52_7 + t_r31_c52_8;
  assign t_r31_c52_11 = t_r31_c52_9 + t_r31_c52_10;
  assign t_r31_c52_12 = t_r31_c52_11 + p_32_53;
  assign out_31_52 = t_r31_c52_12 >> 4;

  assign t_r31_c53_0 = p_30_53 << 1;
  assign t_r31_c53_1 = p_31_52 << 1;
  assign t_r31_c53_2 = p_31_53 << 2;
  assign t_r31_c53_3 = p_31_54 << 1;
  assign t_r31_c53_4 = p_32_53 << 1;
  assign t_r31_c53_5 = t_r31_c53_0 + p_30_52;
  assign t_r31_c53_6 = t_r31_c53_1 + p_30_54;
  assign t_r31_c53_7 = t_r31_c53_2 + t_r31_c53_3;
  assign t_r31_c53_8 = t_r31_c53_4 + p_32_52;
  assign t_r31_c53_9 = t_r31_c53_5 + t_r31_c53_6;
  assign t_r31_c53_10 = t_r31_c53_7 + t_r31_c53_8;
  assign t_r31_c53_11 = t_r31_c53_9 + t_r31_c53_10;
  assign t_r31_c53_12 = t_r31_c53_11 + p_32_54;
  assign out_31_53 = t_r31_c53_12 >> 4;

  assign t_r31_c54_0 = p_30_54 << 1;
  assign t_r31_c54_1 = p_31_53 << 1;
  assign t_r31_c54_2 = p_31_54 << 2;
  assign t_r31_c54_3 = p_31_55 << 1;
  assign t_r31_c54_4 = p_32_54 << 1;
  assign t_r31_c54_5 = t_r31_c54_0 + p_30_53;
  assign t_r31_c54_6 = t_r31_c54_1 + p_30_55;
  assign t_r31_c54_7 = t_r31_c54_2 + t_r31_c54_3;
  assign t_r31_c54_8 = t_r31_c54_4 + p_32_53;
  assign t_r31_c54_9 = t_r31_c54_5 + t_r31_c54_6;
  assign t_r31_c54_10 = t_r31_c54_7 + t_r31_c54_8;
  assign t_r31_c54_11 = t_r31_c54_9 + t_r31_c54_10;
  assign t_r31_c54_12 = t_r31_c54_11 + p_32_55;
  assign out_31_54 = t_r31_c54_12 >> 4;

  assign t_r31_c55_0 = p_30_55 << 1;
  assign t_r31_c55_1 = p_31_54 << 1;
  assign t_r31_c55_2 = p_31_55 << 2;
  assign t_r31_c55_3 = p_31_56 << 1;
  assign t_r31_c55_4 = p_32_55 << 1;
  assign t_r31_c55_5 = t_r31_c55_0 + p_30_54;
  assign t_r31_c55_6 = t_r31_c55_1 + p_30_56;
  assign t_r31_c55_7 = t_r31_c55_2 + t_r31_c55_3;
  assign t_r31_c55_8 = t_r31_c55_4 + p_32_54;
  assign t_r31_c55_9 = t_r31_c55_5 + t_r31_c55_6;
  assign t_r31_c55_10 = t_r31_c55_7 + t_r31_c55_8;
  assign t_r31_c55_11 = t_r31_c55_9 + t_r31_c55_10;
  assign t_r31_c55_12 = t_r31_c55_11 + p_32_56;
  assign out_31_55 = t_r31_c55_12 >> 4;

  assign t_r31_c56_0 = p_30_56 << 1;
  assign t_r31_c56_1 = p_31_55 << 1;
  assign t_r31_c56_2 = p_31_56 << 2;
  assign t_r31_c56_3 = p_31_57 << 1;
  assign t_r31_c56_4 = p_32_56 << 1;
  assign t_r31_c56_5 = t_r31_c56_0 + p_30_55;
  assign t_r31_c56_6 = t_r31_c56_1 + p_30_57;
  assign t_r31_c56_7 = t_r31_c56_2 + t_r31_c56_3;
  assign t_r31_c56_8 = t_r31_c56_4 + p_32_55;
  assign t_r31_c56_9 = t_r31_c56_5 + t_r31_c56_6;
  assign t_r31_c56_10 = t_r31_c56_7 + t_r31_c56_8;
  assign t_r31_c56_11 = t_r31_c56_9 + t_r31_c56_10;
  assign t_r31_c56_12 = t_r31_c56_11 + p_32_57;
  assign out_31_56 = t_r31_c56_12 >> 4;

  assign t_r31_c57_0 = p_30_57 << 1;
  assign t_r31_c57_1 = p_31_56 << 1;
  assign t_r31_c57_2 = p_31_57 << 2;
  assign t_r31_c57_3 = p_31_58 << 1;
  assign t_r31_c57_4 = p_32_57 << 1;
  assign t_r31_c57_5 = t_r31_c57_0 + p_30_56;
  assign t_r31_c57_6 = t_r31_c57_1 + p_30_58;
  assign t_r31_c57_7 = t_r31_c57_2 + t_r31_c57_3;
  assign t_r31_c57_8 = t_r31_c57_4 + p_32_56;
  assign t_r31_c57_9 = t_r31_c57_5 + t_r31_c57_6;
  assign t_r31_c57_10 = t_r31_c57_7 + t_r31_c57_8;
  assign t_r31_c57_11 = t_r31_c57_9 + t_r31_c57_10;
  assign t_r31_c57_12 = t_r31_c57_11 + p_32_58;
  assign out_31_57 = t_r31_c57_12 >> 4;

  assign t_r31_c58_0 = p_30_58 << 1;
  assign t_r31_c58_1 = p_31_57 << 1;
  assign t_r31_c58_2 = p_31_58 << 2;
  assign t_r31_c58_3 = p_31_59 << 1;
  assign t_r31_c58_4 = p_32_58 << 1;
  assign t_r31_c58_5 = t_r31_c58_0 + p_30_57;
  assign t_r31_c58_6 = t_r31_c58_1 + p_30_59;
  assign t_r31_c58_7 = t_r31_c58_2 + t_r31_c58_3;
  assign t_r31_c58_8 = t_r31_c58_4 + p_32_57;
  assign t_r31_c58_9 = t_r31_c58_5 + t_r31_c58_6;
  assign t_r31_c58_10 = t_r31_c58_7 + t_r31_c58_8;
  assign t_r31_c58_11 = t_r31_c58_9 + t_r31_c58_10;
  assign t_r31_c58_12 = t_r31_c58_11 + p_32_59;
  assign out_31_58 = t_r31_c58_12 >> 4;

  assign t_r31_c59_0 = p_30_59 << 1;
  assign t_r31_c59_1 = p_31_58 << 1;
  assign t_r31_c59_2 = p_31_59 << 2;
  assign t_r31_c59_3 = p_31_60 << 1;
  assign t_r31_c59_4 = p_32_59 << 1;
  assign t_r31_c59_5 = t_r31_c59_0 + p_30_58;
  assign t_r31_c59_6 = t_r31_c59_1 + p_30_60;
  assign t_r31_c59_7 = t_r31_c59_2 + t_r31_c59_3;
  assign t_r31_c59_8 = t_r31_c59_4 + p_32_58;
  assign t_r31_c59_9 = t_r31_c59_5 + t_r31_c59_6;
  assign t_r31_c59_10 = t_r31_c59_7 + t_r31_c59_8;
  assign t_r31_c59_11 = t_r31_c59_9 + t_r31_c59_10;
  assign t_r31_c59_12 = t_r31_c59_11 + p_32_60;
  assign out_31_59 = t_r31_c59_12 >> 4;

  assign t_r31_c60_0 = p_30_60 << 1;
  assign t_r31_c60_1 = p_31_59 << 1;
  assign t_r31_c60_2 = p_31_60 << 2;
  assign t_r31_c60_3 = p_31_61 << 1;
  assign t_r31_c60_4 = p_32_60 << 1;
  assign t_r31_c60_5 = t_r31_c60_0 + p_30_59;
  assign t_r31_c60_6 = t_r31_c60_1 + p_30_61;
  assign t_r31_c60_7 = t_r31_c60_2 + t_r31_c60_3;
  assign t_r31_c60_8 = t_r31_c60_4 + p_32_59;
  assign t_r31_c60_9 = t_r31_c60_5 + t_r31_c60_6;
  assign t_r31_c60_10 = t_r31_c60_7 + t_r31_c60_8;
  assign t_r31_c60_11 = t_r31_c60_9 + t_r31_c60_10;
  assign t_r31_c60_12 = t_r31_c60_11 + p_32_61;
  assign out_31_60 = t_r31_c60_12 >> 4;

  assign t_r31_c61_0 = p_30_61 << 1;
  assign t_r31_c61_1 = p_31_60 << 1;
  assign t_r31_c61_2 = p_31_61 << 2;
  assign t_r31_c61_3 = p_31_62 << 1;
  assign t_r31_c61_4 = p_32_61 << 1;
  assign t_r31_c61_5 = t_r31_c61_0 + p_30_60;
  assign t_r31_c61_6 = t_r31_c61_1 + p_30_62;
  assign t_r31_c61_7 = t_r31_c61_2 + t_r31_c61_3;
  assign t_r31_c61_8 = t_r31_c61_4 + p_32_60;
  assign t_r31_c61_9 = t_r31_c61_5 + t_r31_c61_6;
  assign t_r31_c61_10 = t_r31_c61_7 + t_r31_c61_8;
  assign t_r31_c61_11 = t_r31_c61_9 + t_r31_c61_10;
  assign t_r31_c61_12 = t_r31_c61_11 + p_32_62;
  assign out_31_61 = t_r31_c61_12 >> 4;

  assign t_r31_c62_0 = p_30_62 << 1;
  assign t_r31_c62_1 = p_31_61 << 1;
  assign t_r31_c62_2 = p_31_62 << 2;
  assign t_r31_c62_3 = p_31_63 << 1;
  assign t_r31_c62_4 = p_32_62 << 1;
  assign t_r31_c62_5 = t_r31_c62_0 + p_30_61;
  assign t_r31_c62_6 = t_r31_c62_1 + p_30_63;
  assign t_r31_c62_7 = t_r31_c62_2 + t_r31_c62_3;
  assign t_r31_c62_8 = t_r31_c62_4 + p_32_61;
  assign t_r31_c62_9 = t_r31_c62_5 + t_r31_c62_6;
  assign t_r31_c62_10 = t_r31_c62_7 + t_r31_c62_8;
  assign t_r31_c62_11 = t_r31_c62_9 + t_r31_c62_10;
  assign t_r31_c62_12 = t_r31_c62_11 + p_32_63;
  assign out_31_62 = t_r31_c62_12 >> 4;

  assign t_r31_c63_0 = p_30_63 << 1;
  assign t_r31_c63_1 = p_31_62 << 1;
  assign t_r31_c63_2 = p_31_63 << 2;
  assign t_r31_c63_3 = p_31_64 << 1;
  assign t_r31_c63_4 = p_32_63 << 1;
  assign t_r31_c63_5 = t_r31_c63_0 + p_30_62;
  assign t_r31_c63_6 = t_r31_c63_1 + p_30_64;
  assign t_r31_c63_7 = t_r31_c63_2 + t_r31_c63_3;
  assign t_r31_c63_8 = t_r31_c63_4 + p_32_62;
  assign t_r31_c63_9 = t_r31_c63_5 + t_r31_c63_6;
  assign t_r31_c63_10 = t_r31_c63_7 + t_r31_c63_8;
  assign t_r31_c63_11 = t_r31_c63_9 + t_r31_c63_10;
  assign t_r31_c63_12 = t_r31_c63_11 + p_32_64;
  assign out_31_63 = t_r31_c63_12 >> 4;

  assign t_r31_c64_0 = p_30_64 << 1;
  assign t_r31_c64_1 = p_31_63 << 1;
  assign t_r31_c64_2 = p_31_64 << 2;
  assign t_r31_c64_3 = p_31_65 << 1;
  assign t_r31_c64_4 = p_32_64 << 1;
  assign t_r31_c64_5 = t_r31_c64_0 + p_30_63;
  assign t_r31_c64_6 = t_r31_c64_1 + p_30_65;
  assign t_r31_c64_7 = t_r31_c64_2 + t_r31_c64_3;
  assign t_r31_c64_8 = t_r31_c64_4 + p_32_63;
  assign t_r31_c64_9 = t_r31_c64_5 + t_r31_c64_6;
  assign t_r31_c64_10 = t_r31_c64_7 + t_r31_c64_8;
  assign t_r31_c64_11 = t_r31_c64_9 + t_r31_c64_10;
  assign t_r31_c64_12 = t_r31_c64_11 + p_32_65;
  assign out_31_64 = t_r31_c64_12 >> 4;

  assign t_r32_c1_0 = p_31_1 << 1;
  assign t_r32_c1_1 = p_32_0 << 1;
  assign t_r32_c1_2 = p_32_1 << 2;
  assign t_r32_c1_3 = p_32_2 << 1;
  assign t_r32_c1_4 = p_33_1 << 1;
  assign t_r32_c1_5 = t_r32_c1_0 + p_31_0;
  assign t_r32_c1_6 = t_r32_c1_1 + p_31_2;
  assign t_r32_c1_7 = t_r32_c1_2 + t_r32_c1_3;
  assign t_r32_c1_8 = t_r32_c1_4 + p_33_0;
  assign t_r32_c1_9 = t_r32_c1_5 + t_r32_c1_6;
  assign t_r32_c1_10 = t_r32_c1_7 + t_r32_c1_8;
  assign t_r32_c1_11 = t_r32_c1_9 + t_r32_c1_10;
  assign t_r32_c1_12 = t_r32_c1_11 + p_33_2;
  assign out_32_1 = t_r32_c1_12 >> 4;

  assign t_r32_c2_0 = p_31_2 << 1;
  assign t_r32_c2_1 = p_32_1 << 1;
  assign t_r32_c2_2 = p_32_2 << 2;
  assign t_r32_c2_3 = p_32_3 << 1;
  assign t_r32_c2_4 = p_33_2 << 1;
  assign t_r32_c2_5 = t_r32_c2_0 + p_31_1;
  assign t_r32_c2_6 = t_r32_c2_1 + p_31_3;
  assign t_r32_c2_7 = t_r32_c2_2 + t_r32_c2_3;
  assign t_r32_c2_8 = t_r32_c2_4 + p_33_1;
  assign t_r32_c2_9 = t_r32_c2_5 + t_r32_c2_6;
  assign t_r32_c2_10 = t_r32_c2_7 + t_r32_c2_8;
  assign t_r32_c2_11 = t_r32_c2_9 + t_r32_c2_10;
  assign t_r32_c2_12 = t_r32_c2_11 + p_33_3;
  assign out_32_2 = t_r32_c2_12 >> 4;

  assign t_r32_c3_0 = p_31_3 << 1;
  assign t_r32_c3_1 = p_32_2 << 1;
  assign t_r32_c3_2 = p_32_3 << 2;
  assign t_r32_c3_3 = p_32_4 << 1;
  assign t_r32_c3_4 = p_33_3 << 1;
  assign t_r32_c3_5 = t_r32_c3_0 + p_31_2;
  assign t_r32_c3_6 = t_r32_c3_1 + p_31_4;
  assign t_r32_c3_7 = t_r32_c3_2 + t_r32_c3_3;
  assign t_r32_c3_8 = t_r32_c3_4 + p_33_2;
  assign t_r32_c3_9 = t_r32_c3_5 + t_r32_c3_6;
  assign t_r32_c3_10 = t_r32_c3_7 + t_r32_c3_8;
  assign t_r32_c3_11 = t_r32_c3_9 + t_r32_c3_10;
  assign t_r32_c3_12 = t_r32_c3_11 + p_33_4;
  assign out_32_3 = t_r32_c3_12 >> 4;

  assign t_r32_c4_0 = p_31_4 << 1;
  assign t_r32_c4_1 = p_32_3 << 1;
  assign t_r32_c4_2 = p_32_4 << 2;
  assign t_r32_c4_3 = p_32_5 << 1;
  assign t_r32_c4_4 = p_33_4 << 1;
  assign t_r32_c4_5 = t_r32_c4_0 + p_31_3;
  assign t_r32_c4_6 = t_r32_c4_1 + p_31_5;
  assign t_r32_c4_7 = t_r32_c4_2 + t_r32_c4_3;
  assign t_r32_c4_8 = t_r32_c4_4 + p_33_3;
  assign t_r32_c4_9 = t_r32_c4_5 + t_r32_c4_6;
  assign t_r32_c4_10 = t_r32_c4_7 + t_r32_c4_8;
  assign t_r32_c4_11 = t_r32_c4_9 + t_r32_c4_10;
  assign t_r32_c4_12 = t_r32_c4_11 + p_33_5;
  assign out_32_4 = t_r32_c4_12 >> 4;

  assign t_r32_c5_0 = p_31_5 << 1;
  assign t_r32_c5_1 = p_32_4 << 1;
  assign t_r32_c5_2 = p_32_5 << 2;
  assign t_r32_c5_3 = p_32_6 << 1;
  assign t_r32_c5_4 = p_33_5 << 1;
  assign t_r32_c5_5 = t_r32_c5_0 + p_31_4;
  assign t_r32_c5_6 = t_r32_c5_1 + p_31_6;
  assign t_r32_c5_7 = t_r32_c5_2 + t_r32_c5_3;
  assign t_r32_c5_8 = t_r32_c5_4 + p_33_4;
  assign t_r32_c5_9 = t_r32_c5_5 + t_r32_c5_6;
  assign t_r32_c5_10 = t_r32_c5_7 + t_r32_c5_8;
  assign t_r32_c5_11 = t_r32_c5_9 + t_r32_c5_10;
  assign t_r32_c5_12 = t_r32_c5_11 + p_33_6;
  assign out_32_5 = t_r32_c5_12 >> 4;

  assign t_r32_c6_0 = p_31_6 << 1;
  assign t_r32_c6_1 = p_32_5 << 1;
  assign t_r32_c6_2 = p_32_6 << 2;
  assign t_r32_c6_3 = p_32_7 << 1;
  assign t_r32_c6_4 = p_33_6 << 1;
  assign t_r32_c6_5 = t_r32_c6_0 + p_31_5;
  assign t_r32_c6_6 = t_r32_c6_1 + p_31_7;
  assign t_r32_c6_7 = t_r32_c6_2 + t_r32_c6_3;
  assign t_r32_c6_8 = t_r32_c6_4 + p_33_5;
  assign t_r32_c6_9 = t_r32_c6_5 + t_r32_c6_6;
  assign t_r32_c6_10 = t_r32_c6_7 + t_r32_c6_8;
  assign t_r32_c6_11 = t_r32_c6_9 + t_r32_c6_10;
  assign t_r32_c6_12 = t_r32_c6_11 + p_33_7;
  assign out_32_6 = t_r32_c6_12 >> 4;

  assign t_r32_c7_0 = p_31_7 << 1;
  assign t_r32_c7_1 = p_32_6 << 1;
  assign t_r32_c7_2 = p_32_7 << 2;
  assign t_r32_c7_3 = p_32_8 << 1;
  assign t_r32_c7_4 = p_33_7 << 1;
  assign t_r32_c7_5 = t_r32_c7_0 + p_31_6;
  assign t_r32_c7_6 = t_r32_c7_1 + p_31_8;
  assign t_r32_c7_7 = t_r32_c7_2 + t_r32_c7_3;
  assign t_r32_c7_8 = t_r32_c7_4 + p_33_6;
  assign t_r32_c7_9 = t_r32_c7_5 + t_r32_c7_6;
  assign t_r32_c7_10 = t_r32_c7_7 + t_r32_c7_8;
  assign t_r32_c7_11 = t_r32_c7_9 + t_r32_c7_10;
  assign t_r32_c7_12 = t_r32_c7_11 + p_33_8;
  assign out_32_7 = t_r32_c7_12 >> 4;

  assign t_r32_c8_0 = p_31_8 << 1;
  assign t_r32_c8_1 = p_32_7 << 1;
  assign t_r32_c8_2 = p_32_8 << 2;
  assign t_r32_c8_3 = p_32_9 << 1;
  assign t_r32_c8_4 = p_33_8 << 1;
  assign t_r32_c8_5 = t_r32_c8_0 + p_31_7;
  assign t_r32_c8_6 = t_r32_c8_1 + p_31_9;
  assign t_r32_c8_7 = t_r32_c8_2 + t_r32_c8_3;
  assign t_r32_c8_8 = t_r32_c8_4 + p_33_7;
  assign t_r32_c8_9 = t_r32_c8_5 + t_r32_c8_6;
  assign t_r32_c8_10 = t_r32_c8_7 + t_r32_c8_8;
  assign t_r32_c8_11 = t_r32_c8_9 + t_r32_c8_10;
  assign t_r32_c8_12 = t_r32_c8_11 + p_33_9;
  assign out_32_8 = t_r32_c8_12 >> 4;

  assign t_r32_c9_0 = p_31_9 << 1;
  assign t_r32_c9_1 = p_32_8 << 1;
  assign t_r32_c9_2 = p_32_9 << 2;
  assign t_r32_c9_3 = p_32_10 << 1;
  assign t_r32_c9_4 = p_33_9 << 1;
  assign t_r32_c9_5 = t_r32_c9_0 + p_31_8;
  assign t_r32_c9_6 = t_r32_c9_1 + p_31_10;
  assign t_r32_c9_7 = t_r32_c9_2 + t_r32_c9_3;
  assign t_r32_c9_8 = t_r32_c9_4 + p_33_8;
  assign t_r32_c9_9 = t_r32_c9_5 + t_r32_c9_6;
  assign t_r32_c9_10 = t_r32_c9_7 + t_r32_c9_8;
  assign t_r32_c9_11 = t_r32_c9_9 + t_r32_c9_10;
  assign t_r32_c9_12 = t_r32_c9_11 + p_33_10;
  assign out_32_9 = t_r32_c9_12 >> 4;

  assign t_r32_c10_0 = p_31_10 << 1;
  assign t_r32_c10_1 = p_32_9 << 1;
  assign t_r32_c10_2 = p_32_10 << 2;
  assign t_r32_c10_3 = p_32_11 << 1;
  assign t_r32_c10_4 = p_33_10 << 1;
  assign t_r32_c10_5 = t_r32_c10_0 + p_31_9;
  assign t_r32_c10_6 = t_r32_c10_1 + p_31_11;
  assign t_r32_c10_7 = t_r32_c10_2 + t_r32_c10_3;
  assign t_r32_c10_8 = t_r32_c10_4 + p_33_9;
  assign t_r32_c10_9 = t_r32_c10_5 + t_r32_c10_6;
  assign t_r32_c10_10 = t_r32_c10_7 + t_r32_c10_8;
  assign t_r32_c10_11 = t_r32_c10_9 + t_r32_c10_10;
  assign t_r32_c10_12 = t_r32_c10_11 + p_33_11;
  assign out_32_10 = t_r32_c10_12 >> 4;

  assign t_r32_c11_0 = p_31_11 << 1;
  assign t_r32_c11_1 = p_32_10 << 1;
  assign t_r32_c11_2 = p_32_11 << 2;
  assign t_r32_c11_3 = p_32_12 << 1;
  assign t_r32_c11_4 = p_33_11 << 1;
  assign t_r32_c11_5 = t_r32_c11_0 + p_31_10;
  assign t_r32_c11_6 = t_r32_c11_1 + p_31_12;
  assign t_r32_c11_7 = t_r32_c11_2 + t_r32_c11_3;
  assign t_r32_c11_8 = t_r32_c11_4 + p_33_10;
  assign t_r32_c11_9 = t_r32_c11_5 + t_r32_c11_6;
  assign t_r32_c11_10 = t_r32_c11_7 + t_r32_c11_8;
  assign t_r32_c11_11 = t_r32_c11_9 + t_r32_c11_10;
  assign t_r32_c11_12 = t_r32_c11_11 + p_33_12;
  assign out_32_11 = t_r32_c11_12 >> 4;

  assign t_r32_c12_0 = p_31_12 << 1;
  assign t_r32_c12_1 = p_32_11 << 1;
  assign t_r32_c12_2 = p_32_12 << 2;
  assign t_r32_c12_3 = p_32_13 << 1;
  assign t_r32_c12_4 = p_33_12 << 1;
  assign t_r32_c12_5 = t_r32_c12_0 + p_31_11;
  assign t_r32_c12_6 = t_r32_c12_1 + p_31_13;
  assign t_r32_c12_7 = t_r32_c12_2 + t_r32_c12_3;
  assign t_r32_c12_8 = t_r32_c12_4 + p_33_11;
  assign t_r32_c12_9 = t_r32_c12_5 + t_r32_c12_6;
  assign t_r32_c12_10 = t_r32_c12_7 + t_r32_c12_8;
  assign t_r32_c12_11 = t_r32_c12_9 + t_r32_c12_10;
  assign t_r32_c12_12 = t_r32_c12_11 + p_33_13;
  assign out_32_12 = t_r32_c12_12 >> 4;

  assign t_r32_c13_0 = p_31_13 << 1;
  assign t_r32_c13_1 = p_32_12 << 1;
  assign t_r32_c13_2 = p_32_13 << 2;
  assign t_r32_c13_3 = p_32_14 << 1;
  assign t_r32_c13_4 = p_33_13 << 1;
  assign t_r32_c13_5 = t_r32_c13_0 + p_31_12;
  assign t_r32_c13_6 = t_r32_c13_1 + p_31_14;
  assign t_r32_c13_7 = t_r32_c13_2 + t_r32_c13_3;
  assign t_r32_c13_8 = t_r32_c13_4 + p_33_12;
  assign t_r32_c13_9 = t_r32_c13_5 + t_r32_c13_6;
  assign t_r32_c13_10 = t_r32_c13_7 + t_r32_c13_8;
  assign t_r32_c13_11 = t_r32_c13_9 + t_r32_c13_10;
  assign t_r32_c13_12 = t_r32_c13_11 + p_33_14;
  assign out_32_13 = t_r32_c13_12 >> 4;

  assign t_r32_c14_0 = p_31_14 << 1;
  assign t_r32_c14_1 = p_32_13 << 1;
  assign t_r32_c14_2 = p_32_14 << 2;
  assign t_r32_c14_3 = p_32_15 << 1;
  assign t_r32_c14_4 = p_33_14 << 1;
  assign t_r32_c14_5 = t_r32_c14_0 + p_31_13;
  assign t_r32_c14_6 = t_r32_c14_1 + p_31_15;
  assign t_r32_c14_7 = t_r32_c14_2 + t_r32_c14_3;
  assign t_r32_c14_8 = t_r32_c14_4 + p_33_13;
  assign t_r32_c14_9 = t_r32_c14_5 + t_r32_c14_6;
  assign t_r32_c14_10 = t_r32_c14_7 + t_r32_c14_8;
  assign t_r32_c14_11 = t_r32_c14_9 + t_r32_c14_10;
  assign t_r32_c14_12 = t_r32_c14_11 + p_33_15;
  assign out_32_14 = t_r32_c14_12 >> 4;

  assign t_r32_c15_0 = p_31_15 << 1;
  assign t_r32_c15_1 = p_32_14 << 1;
  assign t_r32_c15_2 = p_32_15 << 2;
  assign t_r32_c15_3 = p_32_16 << 1;
  assign t_r32_c15_4 = p_33_15 << 1;
  assign t_r32_c15_5 = t_r32_c15_0 + p_31_14;
  assign t_r32_c15_6 = t_r32_c15_1 + p_31_16;
  assign t_r32_c15_7 = t_r32_c15_2 + t_r32_c15_3;
  assign t_r32_c15_8 = t_r32_c15_4 + p_33_14;
  assign t_r32_c15_9 = t_r32_c15_5 + t_r32_c15_6;
  assign t_r32_c15_10 = t_r32_c15_7 + t_r32_c15_8;
  assign t_r32_c15_11 = t_r32_c15_9 + t_r32_c15_10;
  assign t_r32_c15_12 = t_r32_c15_11 + p_33_16;
  assign out_32_15 = t_r32_c15_12 >> 4;

  assign t_r32_c16_0 = p_31_16 << 1;
  assign t_r32_c16_1 = p_32_15 << 1;
  assign t_r32_c16_2 = p_32_16 << 2;
  assign t_r32_c16_3 = p_32_17 << 1;
  assign t_r32_c16_4 = p_33_16 << 1;
  assign t_r32_c16_5 = t_r32_c16_0 + p_31_15;
  assign t_r32_c16_6 = t_r32_c16_1 + p_31_17;
  assign t_r32_c16_7 = t_r32_c16_2 + t_r32_c16_3;
  assign t_r32_c16_8 = t_r32_c16_4 + p_33_15;
  assign t_r32_c16_9 = t_r32_c16_5 + t_r32_c16_6;
  assign t_r32_c16_10 = t_r32_c16_7 + t_r32_c16_8;
  assign t_r32_c16_11 = t_r32_c16_9 + t_r32_c16_10;
  assign t_r32_c16_12 = t_r32_c16_11 + p_33_17;
  assign out_32_16 = t_r32_c16_12 >> 4;

  assign t_r32_c17_0 = p_31_17 << 1;
  assign t_r32_c17_1 = p_32_16 << 1;
  assign t_r32_c17_2 = p_32_17 << 2;
  assign t_r32_c17_3 = p_32_18 << 1;
  assign t_r32_c17_4 = p_33_17 << 1;
  assign t_r32_c17_5 = t_r32_c17_0 + p_31_16;
  assign t_r32_c17_6 = t_r32_c17_1 + p_31_18;
  assign t_r32_c17_7 = t_r32_c17_2 + t_r32_c17_3;
  assign t_r32_c17_8 = t_r32_c17_4 + p_33_16;
  assign t_r32_c17_9 = t_r32_c17_5 + t_r32_c17_6;
  assign t_r32_c17_10 = t_r32_c17_7 + t_r32_c17_8;
  assign t_r32_c17_11 = t_r32_c17_9 + t_r32_c17_10;
  assign t_r32_c17_12 = t_r32_c17_11 + p_33_18;
  assign out_32_17 = t_r32_c17_12 >> 4;

  assign t_r32_c18_0 = p_31_18 << 1;
  assign t_r32_c18_1 = p_32_17 << 1;
  assign t_r32_c18_2 = p_32_18 << 2;
  assign t_r32_c18_3 = p_32_19 << 1;
  assign t_r32_c18_4 = p_33_18 << 1;
  assign t_r32_c18_5 = t_r32_c18_0 + p_31_17;
  assign t_r32_c18_6 = t_r32_c18_1 + p_31_19;
  assign t_r32_c18_7 = t_r32_c18_2 + t_r32_c18_3;
  assign t_r32_c18_8 = t_r32_c18_4 + p_33_17;
  assign t_r32_c18_9 = t_r32_c18_5 + t_r32_c18_6;
  assign t_r32_c18_10 = t_r32_c18_7 + t_r32_c18_8;
  assign t_r32_c18_11 = t_r32_c18_9 + t_r32_c18_10;
  assign t_r32_c18_12 = t_r32_c18_11 + p_33_19;
  assign out_32_18 = t_r32_c18_12 >> 4;

  assign t_r32_c19_0 = p_31_19 << 1;
  assign t_r32_c19_1 = p_32_18 << 1;
  assign t_r32_c19_2 = p_32_19 << 2;
  assign t_r32_c19_3 = p_32_20 << 1;
  assign t_r32_c19_4 = p_33_19 << 1;
  assign t_r32_c19_5 = t_r32_c19_0 + p_31_18;
  assign t_r32_c19_6 = t_r32_c19_1 + p_31_20;
  assign t_r32_c19_7 = t_r32_c19_2 + t_r32_c19_3;
  assign t_r32_c19_8 = t_r32_c19_4 + p_33_18;
  assign t_r32_c19_9 = t_r32_c19_5 + t_r32_c19_6;
  assign t_r32_c19_10 = t_r32_c19_7 + t_r32_c19_8;
  assign t_r32_c19_11 = t_r32_c19_9 + t_r32_c19_10;
  assign t_r32_c19_12 = t_r32_c19_11 + p_33_20;
  assign out_32_19 = t_r32_c19_12 >> 4;

  assign t_r32_c20_0 = p_31_20 << 1;
  assign t_r32_c20_1 = p_32_19 << 1;
  assign t_r32_c20_2 = p_32_20 << 2;
  assign t_r32_c20_3 = p_32_21 << 1;
  assign t_r32_c20_4 = p_33_20 << 1;
  assign t_r32_c20_5 = t_r32_c20_0 + p_31_19;
  assign t_r32_c20_6 = t_r32_c20_1 + p_31_21;
  assign t_r32_c20_7 = t_r32_c20_2 + t_r32_c20_3;
  assign t_r32_c20_8 = t_r32_c20_4 + p_33_19;
  assign t_r32_c20_9 = t_r32_c20_5 + t_r32_c20_6;
  assign t_r32_c20_10 = t_r32_c20_7 + t_r32_c20_8;
  assign t_r32_c20_11 = t_r32_c20_9 + t_r32_c20_10;
  assign t_r32_c20_12 = t_r32_c20_11 + p_33_21;
  assign out_32_20 = t_r32_c20_12 >> 4;

  assign t_r32_c21_0 = p_31_21 << 1;
  assign t_r32_c21_1 = p_32_20 << 1;
  assign t_r32_c21_2 = p_32_21 << 2;
  assign t_r32_c21_3 = p_32_22 << 1;
  assign t_r32_c21_4 = p_33_21 << 1;
  assign t_r32_c21_5 = t_r32_c21_0 + p_31_20;
  assign t_r32_c21_6 = t_r32_c21_1 + p_31_22;
  assign t_r32_c21_7 = t_r32_c21_2 + t_r32_c21_3;
  assign t_r32_c21_8 = t_r32_c21_4 + p_33_20;
  assign t_r32_c21_9 = t_r32_c21_5 + t_r32_c21_6;
  assign t_r32_c21_10 = t_r32_c21_7 + t_r32_c21_8;
  assign t_r32_c21_11 = t_r32_c21_9 + t_r32_c21_10;
  assign t_r32_c21_12 = t_r32_c21_11 + p_33_22;
  assign out_32_21 = t_r32_c21_12 >> 4;

  assign t_r32_c22_0 = p_31_22 << 1;
  assign t_r32_c22_1 = p_32_21 << 1;
  assign t_r32_c22_2 = p_32_22 << 2;
  assign t_r32_c22_3 = p_32_23 << 1;
  assign t_r32_c22_4 = p_33_22 << 1;
  assign t_r32_c22_5 = t_r32_c22_0 + p_31_21;
  assign t_r32_c22_6 = t_r32_c22_1 + p_31_23;
  assign t_r32_c22_7 = t_r32_c22_2 + t_r32_c22_3;
  assign t_r32_c22_8 = t_r32_c22_4 + p_33_21;
  assign t_r32_c22_9 = t_r32_c22_5 + t_r32_c22_6;
  assign t_r32_c22_10 = t_r32_c22_7 + t_r32_c22_8;
  assign t_r32_c22_11 = t_r32_c22_9 + t_r32_c22_10;
  assign t_r32_c22_12 = t_r32_c22_11 + p_33_23;
  assign out_32_22 = t_r32_c22_12 >> 4;

  assign t_r32_c23_0 = p_31_23 << 1;
  assign t_r32_c23_1 = p_32_22 << 1;
  assign t_r32_c23_2 = p_32_23 << 2;
  assign t_r32_c23_3 = p_32_24 << 1;
  assign t_r32_c23_4 = p_33_23 << 1;
  assign t_r32_c23_5 = t_r32_c23_0 + p_31_22;
  assign t_r32_c23_6 = t_r32_c23_1 + p_31_24;
  assign t_r32_c23_7 = t_r32_c23_2 + t_r32_c23_3;
  assign t_r32_c23_8 = t_r32_c23_4 + p_33_22;
  assign t_r32_c23_9 = t_r32_c23_5 + t_r32_c23_6;
  assign t_r32_c23_10 = t_r32_c23_7 + t_r32_c23_8;
  assign t_r32_c23_11 = t_r32_c23_9 + t_r32_c23_10;
  assign t_r32_c23_12 = t_r32_c23_11 + p_33_24;
  assign out_32_23 = t_r32_c23_12 >> 4;

  assign t_r32_c24_0 = p_31_24 << 1;
  assign t_r32_c24_1 = p_32_23 << 1;
  assign t_r32_c24_2 = p_32_24 << 2;
  assign t_r32_c24_3 = p_32_25 << 1;
  assign t_r32_c24_4 = p_33_24 << 1;
  assign t_r32_c24_5 = t_r32_c24_0 + p_31_23;
  assign t_r32_c24_6 = t_r32_c24_1 + p_31_25;
  assign t_r32_c24_7 = t_r32_c24_2 + t_r32_c24_3;
  assign t_r32_c24_8 = t_r32_c24_4 + p_33_23;
  assign t_r32_c24_9 = t_r32_c24_5 + t_r32_c24_6;
  assign t_r32_c24_10 = t_r32_c24_7 + t_r32_c24_8;
  assign t_r32_c24_11 = t_r32_c24_9 + t_r32_c24_10;
  assign t_r32_c24_12 = t_r32_c24_11 + p_33_25;
  assign out_32_24 = t_r32_c24_12 >> 4;

  assign t_r32_c25_0 = p_31_25 << 1;
  assign t_r32_c25_1 = p_32_24 << 1;
  assign t_r32_c25_2 = p_32_25 << 2;
  assign t_r32_c25_3 = p_32_26 << 1;
  assign t_r32_c25_4 = p_33_25 << 1;
  assign t_r32_c25_5 = t_r32_c25_0 + p_31_24;
  assign t_r32_c25_6 = t_r32_c25_1 + p_31_26;
  assign t_r32_c25_7 = t_r32_c25_2 + t_r32_c25_3;
  assign t_r32_c25_8 = t_r32_c25_4 + p_33_24;
  assign t_r32_c25_9 = t_r32_c25_5 + t_r32_c25_6;
  assign t_r32_c25_10 = t_r32_c25_7 + t_r32_c25_8;
  assign t_r32_c25_11 = t_r32_c25_9 + t_r32_c25_10;
  assign t_r32_c25_12 = t_r32_c25_11 + p_33_26;
  assign out_32_25 = t_r32_c25_12 >> 4;

  assign t_r32_c26_0 = p_31_26 << 1;
  assign t_r32_c26_1 = p_32_25 << 1;
  assign t_r32_c26_2 = p_32_26 << 2;
  assign t_r32_c26_3 = p_32_27 << 1;
  assign t_r32_c26_4 = p_33_26 << 1;
  assign t_r32_c26_5 = t_r32_c26_0 + p_31_25;
  assign t_r32_c26_6 = t_r32_c26_1 + p_31_27;
  assign t_r32_c26_7 = t_r32_c26_2 + t_r32_c26_3;
  assign t_r32_c26_8 = t_r32_c26_4 + p_33_25;
  assign t_r32_c26_9 = t_r32_c26_5 + t_r32_c26_6;
  assign t_r32_c26_10 = t_r32_c26_7 + t_r32_c26_8;
  assign t_r32_c26_11 = t_r32_c26_9 + t_r32_c26_10;
  assign t_r32_c26_12 = t_r32_c26_11 + p_33_27;
  assign out_32_26 = t_r32_c26_12 >> 4;

  assign t_r32_c27_0 = p_31_27 << 1;
  assign t_r32_c27_1 = p_32_26 << 1;
  assign t_r32_c27_2 = p_32_27 << 2;
  assign t_r32_c27_3 = p_32_28 << 1;
  assign t_r32_c27_4 = p_33_27 << 1;
  assign t_r32_c27_5 = t_r32_c27_0 + p_31_26;
  assign t_r32_c27_6 = t_r32_c27_1 + p_31_28;
  assign t_r32_c27_7 = t_r32_c27_2 + t_r32_c27_3;
  assign t_r32_c27_8 = t_r32_c27_4 + p_33_26;
  assign t_r32_c27_9 = t_r32_c27_5 + t_r32_c27_6;
  assign t_r32_c27_10 = t_r32_c27_7 + t_r32_c27_8;
  assign t_r32_c27_11 = t_r32_c27_9 + t_r32_c27_10;
  assign t_r32_c27_12 = t_r32_c27_11 + p_33_28;
  assign out_32_27 = t_r32_c27_12 >> 4;

  assign t_r32_c28_0 = p_31_28 << 1;
  assign t_r32_c28_1 = p_32_27 << 1;
  assign t_r32_c28_2 = p_32_28 << 2;
  assign t_r32_c28_3 = p_32_29 << 1;
  assign t_r32_c28_4 = p_33_28 << 1;
  assign t_r32_c28_5 = t_r32_c28_0 + p_31_27;
  assign t_r32_c28_6 = t_r32_c28_1 + p_31_29;
  assign t_r32_c28_7 = t_r32_c28_2 + t_r32_c28_3;
  assign t_r32_c28_8 = t_r32_c28_4 + p_33_27;
  assign t_r32_c28_9 = t_r32_c28_5 + t_r32_c28_6;
  assign t_r32_c28_10 = t_r32_c28_7 + t_r32_c28_8;
  assign t_r32_c28_11 = t_r32_c28_9 + t_r32_c28_10;
  assign t_r32_c28_12 = t_r32_c28_11 + p_33_29;
  assign out_32_28 = t_r32_c28_12 >> 4;

  assign t_r32_c29_0 = p_31_29 << 1;
  assign t_r32_c29_1 = p_32_28 << 1;
  assign t_r32_c29_2 = p_32_29 << 2;
  assign t_r32_c29_3 = p_32_30 << 1;
  assign t_r32_c29_4 = p_33_29 << 1;
  assign t_r32_c29_5 = t_r32_c29_0 + p_31_28;
  assign t_r32_c29_6 = t_r32_c29_1 + p_31_30;
  assign t_r32_c29_7 = t_r32_c29_2 + t_r32_c29_3;
  assign t_r32_c29_8 = t_r32_c29_4 + p_33_28;
  assign t_r32_c29_9 = t_r32_c29_5 + t_r32_c29_6;
  assign t_r32_c29_10 = t_r32_c29_7 + t_r32_c29_8;
  assign t_r32_c29_11 = t_r32_c29_9 + t_r32_c29_10;
  assign t_r32_c29_12 = t_r32_c29_11 + p_33_30;
  assign out_32_29 = t_r32_c29_12 >> 4;

  assign t_r32_c30_0 = p_31_30 << 1;
  assign t_r32_c30_1 = p_32_29 << 1;
  assign t_r32_c30_2 = p_32_30 << 2;
  assign t_r32_c30_3 = p_32_31 << 1;
  assign t_r32_c30_4 = p_33_30 << 1;
  assign t_r32_c30_5 = t_r32_c30_0 + p_31_29;
  assign t_r32_c30_6 = t_r32_c30_1 + p_31_31;
  assign t_r32_c30_7 = t_r32_c30_2 + t_r32_c30_3;
  assign t_r32_c30_8 = t_r32_c30_4 + p_33_29;
  assign t_r32_c30_9 = t_r32_c30_5 + t_r32_c30_6;
  assign t_r32_c30_10 = t_r32_c30_7 + t_r32_c30_8;
  assign t_r32_c30_11 = t_r32_c30_9 + t_r32_c30_10;
  assign t_r32_c30_12 = t_r32_c30_11 + p_33_31;
  assign out_32_30 = t_r32_c30_12 >> 4;

  assign t_r32_c31_0 = p_31_31 << 1;
  assign t_r32_c31_1 = p_32_30 << 1;
  assign t_r32_c31_2 = p_32_31 << 2;
  assign t_r32_c31_3 = p_32_32 << 1;
  assign t_r32_c31_4 = p_33_31 << 1;
  assign t_r32_c31_5 = t_r32_c31_0 + p_31_30;
  assign t_r32_c31_6 = t_r32_c31_1 + p_31_32;
  assign t_r32_c31_7 = t_r32_c31_2 + t_r32_c31_3;
  assign t_r32_c31_8 = t_r32_c31_4 + p_33_30;
  assign t_r32_c31_9 = t_r32_c31_5 + t_r32_c31_6;
  assign t_r32_c31_10 = t_r32_c31_7 + t_r32_c31_8;
  assign t_r32_c31_11 = t_r32_c31_9 + t_r32_c31_10;
  assign t_r32_c31_12 = t_r32_c31_11 + p_33_32;
  assign out_32_31 = t_r32_c31_12 >> 4;

  assign t_r32_c32_0 = p_31_32 << 1;
  assign t_r32_c32_1 = p_32_31 << 1;
  assign t_r32_c32_2 = p_32_32 << 2;
  assign t_r32_c32_3 = p_32_33 << 1;
  assign t_r32_c32_4 = p_33_32 << 1;
  assign t_r32_c32_5 = t_r32_c32_0 + p_31_31;
  assign t_r32_c32_6 = t_r32_c32_1 + p_31_33;
  assign t_r32_c32_7 = t_r32_c32_2 + t_r32_c32_3;
  assign t_r32_c32_8 = t_r32_c32_4 + p_33_31;
  assign t_r32_c32_9 = t_r32_c32_5 + t_r32_c32_6;
  assign t_r32_c32_10 = t_r32_c32_7 + t_r32_c32_8;
  assign t_r32_c32_11 = t_r32_c32_9 + t_r32_c32_10;
  assign t_r32_c32_12 = t_r32_c32_11 + p_33_33;
  assign out_32_32 = t_r32_c32_12 >> 4;

  assign t_r32_c33_0 = p_31_33 << 1;
  assign t_r32_c33_1 = p_32_32 << 1;
  assign t_r32_c33_2 = p_32_33 << 2;
  assign t_r32_c33_3 = p_32_34 << 1;
  assign t_r32_c33_4 = p_33_33 << 1;
  assign t_r32_c33_5 = t_r32_c33_0 + p_31_32;
  assign t_r32_c33_6 = t_r32_c33_1 + p_31_34;
  assign t_r32_c33_7 = t_r32_c33_2 + t_r32_c33_3;
  assign t_r32_c33_8 = t_r32_c33_4 + p_33_32;
  assign t_r32_c33_9 = t_r32_c33_5 + t_r32_c33_6;
  assign t_r32_c33_10 = t_r32_c33_7 + t_r32_c33_8;
  assign t_r32_c33_11 = t_r32_c33_9 + t_r32_c33_10;
  assign t_r32_c33_12 = t_r32_c33_11 + p_33_34;
  assign out_32_33 = t_r32_c33_12 >> 4;

  assign t_r32_c34_0 = p_31_34 << 1;
  assign t_r32_c34_1 = p_32_33 << 1;
  assign t_r32_c34_2 = p_32_34 << 2;
  assign t_r32_c34_3 = p_32_35 << 1;
  assign t_r32_c34_4 = p_33_34 << 1;
  assign t_r32_c34_5 = t_r32_c34_0 + p_31_33;
  assign t_r32_c34_6 = t_r32_c34_1 + p_31_35;
  assign t_r32_c34_7 = t_r32_c34_2 + t_r32_c34_3;
  assign t_r32_c34_8 = t_r32_c34_4 + p_33_33;
  assign t_r32_c34_9 = t_r32_c34_5 + t_r32_c34_6;
  assign t_r32_c34_10 = t_r32_c34_7 + t_r32_c34_8;
  assign t_r32_c34_11 = t_r32_c34_9 + t_r32_c34_10;
  assign t_r32_c34_12 = t_r32_c34_11 + p_33_35;
  assign out_32_34 = t_r32_c34_12 >> 4;

  assign t_r32_c35_0 = p_31_35 << 1;
  assign t_r32_c35_1 = p_32_34 << 1;
  assign t_r32_c35_2 = p_32_35 << 2;
  assign t_r32_c35_3 = p_32_36 << 1;
  assign t_r32_c35_4 = p_33_35 << 1;
  assign t_r32_c35_5 = t_r32_c35_0 + p_31_34;
  assign t_r32_c35_6 = t_r32_c35_1 + p_31_36;
  assign t_r32_c35_7 = t_r32_c35_2 + t_r32_c35_3;
  assign t_r32_c35_8 = t_r32_c35_4 + p_33_34;
  assign t_r32_c35_9 = t_r32_c35_5 + t_r32_c35_6;
  assign t_r32_c35_10 = t_r32_c35_7 + t_r32_c35_8;
  assign t_r32_c35_11 = t_r32_c35_9 + t_r32_c35_10;
  assign t_r32_c35_12 = t_r32_c35_11 + p_33_36;
  assign out_32_35 = t_r32_c35_12 >> 4;

  assign t_r32_c36_0 = p_31_36 << 1;
  assign t_r32_c36_1 = p_32_35 << 1;
  assign t_r32_c36_2 = p_32_36 << 2;
  assign t_r32_c36_3 = p_32_37 << 1;
  assign t_r32_c36_4 = p_33_36 << 1;
  assign t_r32_c36_5 = t_r32_c36_0 + p_31_35;
  assign t_r32_c36_6 = t_r32_c36_1 + p_31_37;
  assign t_r32_c36_7 = t_r32_c36_2 + t_r32_c36_3;
  assign t_r32_c36_8 = t_r32_c36_4 + p_33_35;
  assign t_r32_c36_9 = t_r32_c36_5 + t_r32_c36_6;
  assign t_r32_c36_10 = t_r32_c36_7 + t_r32_c36_8;
  assign t_r32_c36_11 = t_r32_c36_9 + t_r32_c36_10;
  assign t_r32_c36_12 = t_r32_c36_11 + p_33_37;
  assign out_32_36 = t_r32_c36_12 >> 4;

  assign t_r32_c37_0 = p_31_37 << 1;
  assign t_r32_c37_1 = p_32_36 << 1;
  assign t_r32_c37_2 = p_32_37 << 2;
  assign t_r32_c37_3 = p_32_38 << 1;
  assign t_r32_c37_4 = p_33_37 << 1;
  assign t_r32_c37_5 = t_r32_c37_0 + p_31_36;
  assign t_r32_c37_6 = t_r32_c37_1 + p_31_38;
  assign t_r32_c37_7 = t_r32_c37_2 + t_r32_c37_3;
  assign t_r32_c37_8 = t_r32_c37_4 + p_33_36;
  assign t_r32_c37_9 = t_r32_c37_5 + t_r32_c37_6;
  assign t_r32_c37_10 = t_r32_c37_7 + t_r32_c37_8;
  assign t_r32_c37_11 = t_r32_c37_9 + t_r32_c37_10;
  assign t_r32_c37_12 = t_r32_c37_11 + p_33_38;
  assign out_32_37 = t_r32_c37_12 >> 4;

  assign t_r32_c38_0 = p_31_38 << 1;
  assign t_r32_c38_1 = p_32_37 << 1;
  assign t_r32_c38_2 = p_32_38 << 2;
  assign t_r32_c38_3 = p_32_39 << 1;
  assign t_r32_c38_4 = p_33_38 << 1;
  assign t_r32_c38_5 = t_r32_c38_0 + p_31_37;
  assign t_r32_c38_6 = t_r32_c38_1 + p_31_39;
  assign t_r32_c38_7 = t_r32_c38_2 + t_r32_c38_3;
  assign t_r32_c38_8 = t_r32_c38_4 + p_33_37;
  assign t_r32_c38_9 = t_r32_c38_5 + t_r32_c38_6;
  assign t_r32_c38_10 = t_r32_c38_7 + t_r32_c38_8;
  assign t_r32_c38_11 = t_r32_c38_9 + t_r32_c38_10;
  assign t_r32_c38_12 = t_r32_c38_11 + p_33_39;
  assign out_32_38 = t_r32_c38_12 >> 4;

  assign t_r32_c39_0 = p_31_39 << 1;
  assign t_r32_c39_1 = p_32_38 << 1;
  assign t_r32_c39_2 = p_32_39 << 2;
  assign t_r32_c39_3 = p_32_40 << 1;
  assign t_r32_c39_4 = p_33_39 << 1;
  assign t_r32_c39_5 = t_r32_c39_0 + p_31_38;
  assign t_r32_c39_6 = t_r32_c39_1 + p_31_40;
  assign t_r32_c39_7 = t_r32_c39_2 + t_r32_c39_3;
  assign t_r32_c39_8 = t_r32_c39_4 + p_33_38;
  assign t_r32_c39_9 = t_r32_c39_5 + t_r32_c39_6;
  assign t_r32_c39_10 = t_r32_c39_7 + t_r32_c39_8;
  assign t_r32_c39_11 = t_r32_c39_9 + t_r32_c39_10;
  assign t_r32_c39_12 = t_r32_c39_11 + p_33_40;
  assign out_32_39 = t_r32_c39_12 >> 4;

  assign t_r32_c40_0 = p_31_40 << 1;
  assign t_r32_c40_1 = p_32_39 << 1;
  assign t_r32_c40_2 = p_32_40 << 2;
  assign t_r32_c40_3 = p_32_41 << 1;
  assign t_r32_c40_4 = p_33_40 << 1;
  assign t_r32_c40_5 = t_r32_c40_0 + p_31_39;
  assign t_r32_c40_6 = t_r32_c40_1 + p_31_41;
  assign t_r32_c40_7 = t_r32_c40_2 + t_r32_c40_3;
  assign t_r32_c40_8 = t_r32_c40_4 + p_33_39;
  assign t_r32_c40_9 = t_r32_c40_5 + t_r32_c40_6;
  assign t_r32_c40_10 = t_r32_c40_7 + t_r32_c40_8;
  assign t_r32_c40_11 = t_r32_c40_9 + t_r32_c40_10;
  assign t_r32_c40_12 = t_r32_c40_11 + p_33_41;
  assign out_32_40 = t_r32_c40_12 >> 4;

  assign t_r32_c41_0 = p_31_41 << 1;
  assign t_r32_c41_1 = p_32_40 << 1;
  assign t_r32_c41_2 = p_32_41 << 2;
  assign t_r32_c41_3 = p_32_42 << 1;
  assign t_r32_c41_4 = p_33_41 << 1;
  assign t_r32_c41_5 = t_r32_c41_0 + p_31_40;
  assign t_r32_c41_6 = t_r32_c41_1 + p_31_42;
  assign t_r32_c41_7 = t_r32_c41_2 + t_r32_c41_3;
  assign t_r32_c41_8 = t_r32_c41_4 + p_33_40;
  assign t_r32_c41_9 = t_r32_c41_5 + t_r32_c41_6;
  assign t_r32_c41_10 = t_r32_c41_7 + t_r32_c41_8;
  assign t_r32_c41_11 = t_r32_c41_9 + t_r32_c41_10;
  assign t_r32_c41_12 = t_r32_c41_11 + p_33_42;
  assign out_32_41 = t_r32_c41_12 >> 4;

  assign t_r32_c42_0 = p_31_42 << 1;
  assign t_r32_c42_1 = p_32_41 << 1;
  assign t_r32_c42_2 = p_32_42 << 2;
  assign t_r32_c42_3 = p_32_43 << 1;
  assign t_r32_c42_4 = p_33_42 << 1;
  assign t_r32_c42_5 = t_r32_c42_0 + p_31_41;
  assign t_r32_c42_6 = t_r32_c42_1 + p_31_43;
  assign t_r32_c42_7 = t_r32_c42_2 + t_r32_c42_3;
  assign t_r32_c42_8 = t_r32_c42_4 + p_33_41;
  assign t_r32_c42_9 = t_r32_c42_5 + t_r32_c42_6;
  assign t_r32_c42_10 = t_r32_c42_7 + t_r32_c42_8;
  assign t_r32_c42_11 = t_r32_c42_9 + t_r32_c42_10;
  assign t_r32_c42_12 = t_r32_c42_11 + p_33_43;
  assign out_32_42 = t_r32_c42_12 >> 4;

  assign t_r32_c43_0 = p_31_43 << 1;
  assign t_r32_c43_1 = p_32_42 << 1;
  assign t_r32_c43_2 = p_32_43 << 2;
  assign t_r32_c43_3 = p_32_44 << 1;
  assign t_r32_c43_4 = p_33_43 << 1;
  assign t_r32_c43_5 = t_r32_c43_0 + p_31_42;
  assign t_r32_c43_6 = t_r32_c43_1 + p_31_44;
  assign t_r32_c43_7 = t_r32_c43_2 + t_r32_c43_3;
  assign t_r32_c43_8 = t_r32_c43_4 + p_33_42;
  assign t_r32_c43_9 = t_r32_c43_5 + t_r32_c43_6;
  assign t_r32_c43_10 = t_r32_c43_7 + t_r32_c43_8;
  assign t_r32_c43_11 = t_r32_c43_9 + t_r32_c43_10;
  assign t_r32_c43_12 = t_r32_c43_11 + p_33_44;
  assign out_32_43 = t_r32_c43_12 >> 4;

  assign t_r32_c44_0 = p_31_44 << 1;
  assign t_r32_c44_1 = p_32_43 << 1;
  assign t_r32_c44_2 = p_32_44 << 2;
  assign t_r32_c44_3 = p_32_45 << 1;
  assign t_r32_c44_4 = p_33_44 << 1;
  assign t_r32_c44_5 = t_r32_c44_0 + p_31_43;
  assign t_r32_c44_6 = t_r32_c44_1 + p_31_45;
  assign t_r32_c44_7 = t_r32_c44_2 + t_r32_c44_3;
  assign t_r32_c44_8 = t_r32_c44_4 + p_33_43;
  assign t_r32_c44_9 = t_r32_c44_5 + t_r32_c44_6;
  assign t_r32_c44_10 = t_r32_c44_7 + t_r32_c44_8;
  assign t_r32_c44_11 = t_r32_c44_9 + t_r32_c44_10;
  assign t_r32_c44_12 = t_r32_c44_11 + p_33_45;
  assign out_32_44 = t_r32_c44_12 >> 4;

  assign t_r32_c45_0 = p_31_45 << 1;
  assign t_r32_c45_1 = p_32_44 << 1;
  assign t_r32_c45_2 = p_32_45 << 2;
  assign t_r32_c45_3 = p_32_46 << 1;
  assign t_r32_c45_4 = p_33_45 << 1;
  assign t_r32_c45_5 = t_r32_c45_0 + p_31_44;
  assign t_r32_c45_6 = t_r32_c45_1 + p_31_46;
  assign t_r32_c45_7 = t_r32_c45_2 + t_r32_c45_3;
  assign t_r32_c45_8 = t_r32_c45_4 + p_33_44;
  assign t_r32_c45_9 = t_r32_c45_5 + t_r32_c45_6;
  assign t_r32_c45_10 = t_r32_c45_7 + t_r32_c45_8;
  assign t_r32_c45_11 = t_r32_c45_9 + t_r32_c45_10;
  assign t_r32_c45_12 = t_r32_c45_11 + p_33_46;
  assign out_32_45 = t_r32_c45_12 >> 4;

  assign t_r32_c46_0 = p_31_46 << 1;
  assign t_r32_c46_1 = p_32_45 << 1;
  assign t_r32_c46_2 = p_32_46 << 2;
  assign t_r32_c46_3 = p_32_47 << 1;
  assign t_r32_c46_4 = p_33_46 << 1;
  assign t_r32_c46_5 = t_r32_c46_0 + p_31_45;
  assign t_r32_c46_6 = t_r32_c46_1 + p_31_47;
  assign t_r32_c46_7 = t_r32_c46_2 + t_r32_c46_3;
  assign t_r32_c46_8 = t_r32_c46_4 + p_33_45;
  assign t_r32_c46_9 = t_r32_c46_5 + t_r32_c46_6;
  assign t_r32_c46_10 = t_r32_c46_7 + t_r32_c46_8;
  assign t_r32_c46_11 = t_r32_c46_9 + t_r32_c46_10;
  assign t_r32_c46_12 = t_r32_c46_11 + p_33_47;
  assign out_32_46 = t_r32_c46_12 >> 4;

  assign t_r32_c47_0 = p_31_47 << 1;
  assign t_r32_c47_1 = p_32_46 << 1;
  assign t_r32_c47_2 = p_32_47 << 2;
  assign t_r32_c47_3 = p_32_48 << 1;
  assign t_r32_c47_4 = p_33_47 << 1;
  assign t_r32_c47_5 = t_r32_c47_0 + p_31_46;
  assign t_r32_c47_6 = t_r32_c47_1 + p_31_48;
  assign t_r32_c47_7 = t_r32_c47_2 + t_r32_c47_3;
  assign t_r32_c47_8 = t_r32_c47_4 + p_33_46;
  assign t_r32_c47_9 = t_r32_c47_5 + t_r32_c47_6;
  assign t_r32_c47_10 = t_r32_c47_7 + t_r32_c47_8;
  assign t_r32_c47_11 = t_r32_c47_9 + t_r32_c47_10;
  assign t_r32_c47_12 = t_r32_c47_11 + p_33_48;
  assign out_32_47 = t_r32_c47_12 >> 4;

  assign t_r32_c48_0 = p_31_48 << 1;
  assign t_r32_c48_1 = p_32_47 << 1;
  assign t_r32_c48_2 = p_32_48 << 2;
  assign t_r32_c48_3 = p_32_49 << 1;
  assign t_r32_c48_4 = p_33_48 << 1;
  assign t_r32_c48_5 = t_r32_c48_0 + p_31_47;
  assign t_r32_c48_6 = t_r32_c48_1 + p_31_49;
  assign t_r32_c48_7 = t_r32_c48_2 + t_r32_c48_3;
  assign t_r32_c48_8 = t_r32_c48_4 + p_33_47;
  assign t_r32_c48_9 = t_r32_c48_5 + t_r32_c48_6;
  assign t_r32_c48_10 = t_r32_c48_7 + t_r32_c48_8;
  assign t_r32_c48_11 = t_r32_c48_9 + t_r32_c48_10;
  assign t_r32_c48_12 = t_r32_c48_11 + p_33_49;
  assign out_32_48 = t_r32_c48_12 >> 4;

  assign t_r32_c49_0 = p_31_49 << 1;
  assign t_r32_c49_1 = p_32_48 << 1;
  assign t_r32_c49_2 = p_32_49 << 2;
  assign t_r32_c49_3 = p_32_50 << 1;
  assign t_r32_c49_4 = p_33_49 << 1;
  assign t_r32_c49_5 = t_r32_c49_0 + p_31_48;
  assign t_r32_c49_6 = t_r32_c49_1 + p_31_50;
  assign t_r32_c49_7 = t_r32_c49_2 + t_r32_c49_3;
  assign t_r32_c49_8 = t_r32_c49_4 + p_33_48;
  assign t_r32_c49_9 = t_r32_c49_5 + t_r32_c49_6;
  assign t_r32_c49_10 = t_r32_c49_7 + t_r32_c49_8;
  assign t_r32_c49_11 = t_r32_c49_9 + t_r32_c49_10;
  assign t_r32_c49_12 = t_r32_c49_11 + p_33_50;
  assign out_32_49 = t_r32_c49_12 >> 4;

  assign t_r32_c50_0 = p_31_50 << 1;
  assign t_r32_c50_1 = p_32_49 << 1;
  assign t_r32_c50_2 = p_32_50 << 2;
  assign t_r32_c50_3 = p_32_51 << 1;
  assign t_r32_c50_4 = p_33_50 << 1;
  assign t_r32_c50_5 = t_r32_c50_0 + p_31_49;
  assign t_r32_c50_6 = t_r32_c50_1 + p_31_51;
  assign t_r32_c50_7 = t_r32_c50_2 + t_r32_c50_3;
  assign t_r32_c50_8 = t_r32_c50_4 + p_33_49;
  assign t_r32_c50_9 = t_r32_c50_5 + t_r32_c50_6;
  assign t_r32_c50_10 = t_r32_c50_7 + t_r32_c50_8;
  assign t_r32_c50_11 = t_r32_c50_9 + t_r32_c50_10;
  assign t_r32_c50_12 = t_r32_c50_11 + p_33_51;
  assign out_32_50 = t_r32_c50_12 >> 4;

  assign t_r32_c51_0 = p_31_51 << 1;
  assign t_r32_c51_1 = p_32_50 << 1;
  assign t_r32_c51_2 = p_32_51 << 2;
  assign t_r32_c51_3 = p_32_52 << 1;
  assign t_r32_c51_4 = p_33_51 << 1;
  assign t_r32_c51_5 = t_r32_c51_0 + p_31_50;
  assign t_r32_c51_6 = t_r32_c51_1 + p_31_52;
  assign t_r32_c51_7 = t_r32_c51_2 + t_r32_c51_3;
  assign t_r32_c51_8 = t_r32_c51_4 + p_33_50;
  assign t_r32_c51_9 = t_r32_c51_5 + t_r32_c51_6;
  assign t_r32_c51_10 = t_r32_c51_7 + t_r32_c51_8;
  assign t_r32_c51_11 = t_r32_c51_9 + t_r32_c51_10;
  assign t_r32_c51_12 = t_r32_c51_11 + p_33_52;
  assign out_32_51 = t_r32_c51_12 >> 4;

  assign t_r32_c52_0 = p_31_52 << 1;
  assign t_r32_c52_1 = p_32_51 << 1;
  assign t_r32_c52_2 = p_32_52 << 2;
  assign t_r32_c52_3 = p_32_53 << 1;
  assign t_r32_c52_4 = p_33_52 << 1;
  assign t_r32_c52_5 = t_r32_c52_0 + p_31_51;
  assign t_r32_c52_6 = t_r32_c52_1 + p_31_53;
  assign t_r32_c52_7 = t_r32_c52_2 + t_r32_c52_3;
  assign t_r32_c52_8 = t_r32_c52_4 + p_33_51;
  assign t_r32_c52_9 = t_r32_c52_5 + t_r32_c52_6;
  assign t_r32_c52_10 = t_r32_c52_7 + t_r32_c52_8;
  assign t_r32_c52_11 = t_r32_c52_9 + t_r32_c52_10;
  assign t_r32_c52_12 = t_r32_c52_11 + p_33_53;
  assign out_32_52 = t_r32_c52_12 >> 4;

  assign t_r32_c53_0 = p_31_53 << 1;
  assign t_r32_c53_1 = p_32_52 << 1;
  assign t_r32_c53_2 = p_32_53 << 2;
  assign t_r32_c53_3 = p_32_54 << 1;
  assign t_r32_c53_4 = p_33_53 << 1;
  assign t_r32_c53_5 = t_r32_c53_0 + p_31_52;
  assign t_r32_c53_6 = t_r32_c53_1 + p_31_54;
  assign t_r32_c53_7 = t_r32_c53_2 + t_r32_c53_3;
  assign t_r32_c53_8 = t_r32_c53_4 + p_33_52;
  assign t_r32_c53_9 = t_r32_c53_5 + t_r32_c53_6;
  assign t_r32_c53_10 = t_r32_c53_7 + t_r32_c53_8;
  assign t_r32_c53_11 = t_r32_c53_9 + t_r32_c53_10;
  assign t_r32_c53_12 = t_r32_c53_11 + p_33_54;
  assign out_32_53 = t_r32_c53_12 >> 4;

  assign t_r32_c54_0 = p_31_54 << 1;
  assign t_r32_c54_1 = p_32_53 << 1;
  assign t_r32_c54_2 = p_32_54 << 2;
  assign t_r32_c54_3 = p_32_55 << 1;
  assign t_r32_c54_4 = p_33_54 << 1;
  assign t_r32_c54_5 = t_r32_c54_0 + p_31_53;
  assign t_r32_c54_6 = t_r32_c54_1 + p_31_55;
  assign t_r32_c54_7 = t_r32_c54_2 + t_r32_c54_3;
  assign t_r32_c54_8 = t_r32_c54_4 + p_33_53;
  assign t_r32_c54_9 = t_r32_c54_5 + t_r32_c54_6;
  assign t_r32_c54_10 = t_r32_c54_7 + t_r32_c54_8;
  assign t_r32_c54_11 = t_r32_c54_9 + t_r32_c54_10;
  assign t_r32_c54_12 = t_r32_c54_11 + p_33_55;
  assign out_32_54 = t_r32_c54_12 >> 4;

  assign t_r32_c55_0 = p_31_55 << 1;
  assign t_r32_c55_1 = p_32_54 << 1;
  assign t_r32_c55_2 = p_32_55 << 2;
  assign t_r32_c55_3 = p_32_56 << 1;
  assign t_r32_c55_4 = p_33_55 << 1;
  assign t_r32_c55_5 = t_r32_c55_0 + p_31_54;
  assign t_r32_c55_6 = t_r32_c55_1 + p_31_56;
  assign t_r32_c55_7 = t_r32_c55_2 + t_r32_c55_3;
  assign t_r32_c55_8 = t_r32_c55_4 + p_33_54;
  assign t_r32_c55_9 = t_r32_c55_5 + t_r32_c55_6;
  assign t_r32_c55_10 = t_r32_c55_7 + t_r32_c55_8;
  assign t_r32_c55_11 = t_r32_c55_9 + t_r32_c55_10;
  assign t_r32_c55_12 = t_r32_c55_11 + p_33_56;
  assign out_32_55 = t_r32_c55_12 >> 4;

  assign t_r32_c56_0 = p_31_56 << 1;
  assign t_r32_c56_1 = p_32_55 << 1;
  assign t_r32_c56_2 = p_32_56 << 2;
  assign t_r32_c56_3 = p_32_57 << 1;
  assign t_r32_c56_4 = p_33_56 << 1;
  assign t_r32_c56_5 = t_r32_c56_0 + p_31_55;
  assign t_r32_c56_6 = t_r32_c56_1 + p_31_57;
  assign t_r32_c56_7 = t_r32_c56_2 + t_r32_c56_3;
  assign t_r32_c56_8 = t_r32_c56_4 + p_33_55;
  assign t_r32_c56_9 = t_r32_c56_5 + t_r32_c56_6;
  assign t_r32_c56_10 = t_r32_c56_7 + t_r32_c56_8;
  assign t_r32_c56_11 = t_r32_c56_9 + t_r32_c56_10;
  assign t_r32_c56_12 = t_r32_c56_11 + p_33_57;
  assign out_32_56 = t_r32_c56_12 >> 4;

  assign t_r32_c57_0 = p_31_57 << 1;
  assign t_r32_c57_1 = p_32_56 << 1;
  assign t_r32_c57_2 = p_32_57 << 2;
  assign t_r32_c57_3 = p_32_58 << 1;
  assign t_r32_c57_4 = p_33_57 << 1;
  assign t_r32_c57_5 = t_r32_c57_0 + p_31_56;
  assign t_r32_c57_6 = t_r32_c57_1 + p_31_58;
  assign t_r32_c57_7 = t_r32_c57_2 + t_r32_c57_3;
  assign t_r32_c57_8 = t_r32_c57_4 + p_33_56;
  assign t_r32_c57_9 = t_r32_c57_5 + t_r32_c57_6;
  assign t_r32_c57_10 = t_r32_c57_7 + t_r32_c57_8;
  assign t_r32_c57_11 = t_r32_c57_9 + t_r32_c57_10;
  assign t_r32_c57_12 = t_r32_c57_11 + p_33_58;
  assign out_32_57 = t_r32_c57_12 >> 4;

  assign t_r32_c58_0 = p_31_58 << 1;
  assign t_r32_c58_1 = p_32_57 << 1;
  assign t_r32_c58_2 = p_32_58 << 2;
  assign t_r32_c58_3 = p_32_59 << 1;
  assign t_r32_c58_4 = p_33_58 << 1;
  assign t_r32_c58_5 = t_r32_c58_0 + p_31_57;
  assign t_r32_c58_6 = t_r32_c58_1 + p_31_59;
  assign t_r32_c58_7 = t_r32_c58_2 + t_r32_c58_3;
  assign t_r32_c58_8 = t_r32_c58_4 + p_33_57;
  assign t_r32_c58_9 = t_r32_c58_5 + t_r32_c58_6;
  assign t_r32_c58_10 = t_r32_c58_7 + t_r32_c58_8;
  assign t_r32_c58_11 = t_r32_c58_9 + t_r32_c58_10;
  assign t_r32_c58_12 = t_r32_c58_11 + p_33_59;
  assign out_32_58 = t_r32_c58_12 >> 4;

  assign t_r32_c59_0 = p_31_59 << 1;
  assign t_r32_c59_1 = p_32_58 << 1;
  assign t_r32_c59_2 = p_32_59 << 2;
  assign t_r32_c59_3 = p_32_60 << 1;
  assign t_r32_c59_4 = p_33_59 << 1;
  assign t_r32_c59_5 = t_r32_c59_0 + p_31_58;
  assign t_r32_c59_6 = t_r32_c59_1 + p_31_60;
  assign t_r32_c59_7 = t_r32_c59_2 + t_r32_c59_3;
  assign t_r32_c59_8 = t_r32_c59_4 + p_33_58;
  assign t_r32_c59_9 = t_r32_c59_5 + t_r32_c59_6;
  assign t_r32_c59_10 = t_r32_c59_7 + t_r32_c59_8;
  assign t_r32_c59_11 = t_r32_c59_9 + t_r32_c59_10;
  assign t_r32_c59_12 = t_r32_c59_11 + p_33_60;
  assign out_32_59 = t_r32_c59_12 >> 4;

  assign t_r32_c60_0 = p_31_60 << 1;
  assign t_r32_c60_1 = p_32_59 << 1;
  assign t_r32_c60_2 = p_32_60 << 2;
  assign t_r32_c60_3 = p_32_61 << 1;
  assign t_r32_c60_4 = p_33_60 << 1;
  assign t_r32_c60_5 = t_r32_c60_0 + p_31_59;
  assign t_r32_c60_6 = t_r32_c60_1 + p_31_61;
  assign t_r32_c60_7 = t_r32_c60_2 + t_r32_c60_3;
  assign t_r32_c60_8 = t_r32_c60_4 + p_33_59;
  assign t_r32_c60_9 = t_r32_c60_5 + t_r32_c60_6;
  assign t_r32_c60_10 = t_r32_c60_7 + t_r32_c60_8;
  assign t_r32_c60_11 = t_r32_c60_9 + t_r32_c60_10;
  assign t_r32_c60_12 = t_r32_c60_11 + p_33_61;
  assign out_32_60 = t_r32_c60_12 >> 4;

  assign t_r32_c61_0 = p_31_61 << 1;
  assign t_r32_c61_1 = p_32_60 << 1;
  assign t_r32_c61_2 = p_32_61 << 2;
  assign t_r32_c61_3 = p_32_62 << 1;
  assign t_r32_c61_4 = p_33_61 << 1;
  assign t_r32_c61_5 = t_r32_c61_0 + p_31_60;
  assign t_r32_c61_6 = t_r32_c61_1 + p_31_62;
  assign t_r32_c61_7 = t_r32_c61_2 + t_r32_c61_3;
  assign t_r32_c61_8 = t_r32_c61_4 + p_33_60;
  assign t_r32_c61_9 = t_r32_c61_5 + t_r32_c61_6;
  assign t_r32_c61_10 = t_r32_c61_7 + t_r32_c61_8;
  assign t_r32_c61_11 = t_r32_c61_9 + t_r32_c61_10;
  assign t_r32_c61_12 = t_r32_c61_11 + p_33_62;
  assign out_32_61 = t_r32_c61_12 >> 4;

  assign t_r32_c62_0 = p_31_62 << 1;
  assign t_r32_c62_1 = p_32_61 << 1;
  assign t_r32_c62_2 = p_32_62 << 2;
  assign t_r32_c62_3 = p_32_63 << 1;
  assign t_r32_c62_4 = p_33_62 << 1;
  assign t_r32_c62_5 = t_r32_c62_0 + p_31_61;
  assign t_r32_c62_6 = t_r32_c62_1 + p_31_63;
  assign t_r32_c62_7 = t_r32_c62_2 + t_r32_c62_3;
  assign t_r32_c62_8 = t_r32_c62_4 + p_33_61;
  assign t_r32_c62_9 = t_r32_c62_5 + t_r32_c62_6;
  assign t_r32_c62_10 = t_r32_c62_7 + t_r32_c62_8;
  assign t_r32_c62_11 = t_r32_c62_9 + t_r32_c62_10;
  assign t_r32_c62_12 = t_r32_c62_11 + p_33_63;
  assign out_32_62 = t_r32_c62_12 >> 4;

  assign t_r32_c63_0 = p_31_63 << 1;
  assign t_r32_c63_1 = p_32_62 << 1;
  assign t_r32_c63_2 = p_32_63 << 2;
  assign t_r32_c63_3 = p_32_64 << 1;
  assign t_r32_c63_4 = p_33_63 << 1;
  assign t_r32_c63_5 = t_r32_c63_0 + p_31_62;
  assign t_r32_c63_6 = t_r32_c63_1 + p_31_64;
  assign t_r32_c63_7 = t_r32_c63_2 + t_r32_c63_3;
  assign t_r32_c63_8 = t_r32_c63_4 + p_33_62;
  assign t_r32_c63_9 = t_r32_c63_5 + t_r32_c63_6;
  assign t_r32_c63_10 = t_r32_c63_7 + t_r32_c63_8;
  assign t_r32_c63_11 = t_r32_c63_9 + t_r32_c63_10;
  assign t_r32_c63_12 = t_r32_c63_11 + p_33_64;
  assign out_32_63 = t_r32_c63_12 >> 4;

  assign t_r32_c64_0 = p_31_64 << 1;
  assign t_r32_c64_1 = p_32_63 << 1;
  assign t_r32_c64_2 = p_32_64 << 2;
  assign t_r32_c64_3 = p_32_65 << 1;
  assign t_r32_c64_4 = p_33_64 << 1;
  assign t_r32_c64_5 = t_r32_c64_0 + p_31_63;
  assign t_r32_c64_6 = t_r32_c64_1 + p_31_65;
  assign t_r32_c64_7 = t_r32_c64_2 + t_r32_c64_3;
  assign t_r32_c64_8 = t_r32_c64_4 + p_33_63;
  assign t_r32_c64_9 = t_r32_c64_5 + t_r32_c64_6;
  assign t_r32_c64_10 = t_r32_c64_7 + t_r32_c64_8;
  assign t_r32_c64_11 = t_r32_c64_9 + t_r32_c64_10;
  assign t_r32_c64_12 = t_r32_c64_11 + p_33_65;
  assign out_32_64 = t_r32_c64_12 >> 4;

  assign t_r33_c1_0 = p_32_1 << 1;
  assign t_r33_c1_1 = p_33_0 << 1;
  assign t_r33_c1_2 = p_33_1 << 2;
  assign t_r33_c1_3 = p_33_2 << 1;
  assign t_r33_c1_4 = p_34_1 << 1;
  assign t_r33_c1_5 = t_r33_c1_0 + p_32_0;
  assign t_r33_c1_6 = t_r33_c1_1 + p_32_2;
  assign t_r33_c1_7 = t_r33_c1_2 + t_r33_c1_3;
  assign t_r33_c1_8 = t_r33_c1_4 + p_34_0;
  assign t_r33_c1_9 = t_r33_c1_5 + t_r33_c1_6;
  assign t_r33_c1_10 = t_r33_c1_7 + t_r33_c1_8;
  assign t_r33_c1_11 = t_r33_c1_9 + t_r33_c1_10;
  assign t_r33_c1_12 = t_r33_c1_11 + p_34_2;
  assign out_33_1 = t_r33_c1_12 >> 4;

  assign t_r33_c2_0 = p_32_2 << 1;
  assign t_r33_c2_1 = p_33_1 << 1;
  assign t_r33_c2_2 = p_33_2 << 2;
  assign t_r33_c2_3 = p_33_3 << 1;
  assign t_r33_c2_4 = p_34_2 << 1;
  assign t_r33_c2_5 = t_r33_c2_0 + p_32_1;
  assign t_r33_c2_6 = t_r33_c2_1 + p_32_3;
  assign t_r33_c2_7 = t_r33_c2_2 + t_r33_c2_3;
  assign t_r33_c2_8 = t_r33_c2_4 + p_34_1;
  assign t_r33_c2_9 = t_r33_c2_5 + t_r33_c2_6;
  assign t_r33_c2_10 = t_r33_c2_7 + t_r33_c2_8;
  assign t_r33_c2_11 = t_r33_c2_9 + t_r33_c2_10;
  assign t_r33_c2_12 = t_r33_c2_11 + p_34_3;
  assign out_33_2 = t_r33_c2_12 >> 4;

  assign t_r33_c3_0 = p_32_3 << 1;
  assign t_r33_c3_1 = p_33_2 << 1;
  assign t_r33_c3_2 = p_33_3 << 2;
  assign t_r33_c3_3 = p_33_4 << 1;
  assign t_r33_c3_4 = p_34_3 << 1;
  assign t_r33_c3_5 = t_r33_c3_0 + p_32_2;
  assign t_r33_c3_6 = t_r33_c3_1 + p_32_4;
  assign t_r33_c3_7 = t_r33_c3_2 + t_r33_c3_3;
  assign t_r33_c3_8 = t_r33_c3_4 + p_34_2;
  assign t_r33_c3_9 = t_r33_c3_5 + t_r33_c3_6;
  assign t_r33_c3_10 = t_r33_c3_7 + t_r33_c3_8;
  assign t_r33_c3_11 = t_r33_c3_9 + t_r33_c3_10;
  assign t_r33_c3_12 = t_r33_c3_11 + p_34_4;
  assign out_33_3 = t_r33_c3_12 >> 4;

  assign t_r33_c4_0 = p_32_4 << 1;
  assign t_r33_c4_1 = p_33_3 << 1;
  assign t_r33_c4_2 = p_33_4 << 2;
  assign t_r33_c4_3 = p_33_5 << 1;
  assign t_r33_c4_4 = p_34_4 << 1;
  assign t_r33_c4_5 = t_r33_c4_0 + p_32_3;
  assign t_r33_c4_6 = t_r33_c4_1 + p_32_5;
  assign t_r33_c4_7 = t_r33_c4_2 + t_r33_c4_3;
  assign t_r33_c4_8 = t_r33_c4_4 + p_34_3;
  assign t_r33_c4_9 = t_r33_c4_5 + t_r33_c4_6;
  assign t_r33_c4_10 = t_r33_c4_7 + t_r33_c4_8;
  assign t_r33_c4_11 = t_r33_c4_9 + t_r33_c4_10;
  assign t_r33_c4_12 = t_r33_c4_11 + p_34_5;
  assign out_33_4 = t_r33_c4_12 >> 4;

  assign t_r33_c5_0 = p_32_5 << 1;
  assign t_r33_c5_1 = p_33_4 << 1;
  assign t_r33_c5_2 = p_33_5 << 2;
  assign t_r33_c5_3 = p_33_6 << 1;
  assign t_r33_c5_4 = p_34_5 << 1;
  assign t_r33_c5_5 = t_r33_c5_0 + p_32_4;
  assign t_r33_c5_6 = t_r33_c5_1 + p_32_6;
  assign t_r33_c5_7 = t_r33_c5_2 + t_r33_c5_3;
  assign t_r33_c5_8 = t_r33_c5_4 + p_34_4;
  assign t_r33_c5_9 = t_r33_c5_5 + t_r33_c5_6;
  assign t_r33_c5_10 = t_r33_c5_7 + t_r33_c5_8;
  assign t_r33_c5_11 = t_r33_c5_9 + t_r33_c5_10;
  assign t_r33_c5_12 = t_r33_c5_11 + p_34_6;
  assign out_33_5 = t_r33_c5_12 >> 4;

  assign t_r33_c6_0 = p_32_6 << 1;
  assign t_r33_c6_1 = p_33_5 << 1;
  assign t_r33_c6_2 = p_33_6 << 2;
  assign t_r33_c6_3 = p_33_7 << 1;
  assign t_r33_c6_4 = p_34_6 << 1;
  assign t_r33_c6_5 = t_r33_c6_0 + p_32_5;
  assign t_r33_c6_6 = t_r33_c6_1 + p_32_7;
  assign t_r33_c6_7 = t_r33_c6_2 + t_r33_c6_3;
  assign t_r33_c6_8 = t_r33_c6_4 + p_34_5;
  assign t_r33_c6_9 = t_r33_c6_5 + t_r33_c6_6;
  assign t_r33_c6_10 = t_r33_c6_7 + t_r33_c6_8;
  assign t_r33_c6_11 = t_r33_c6_9 + t_r33_c6_10;
  assign t_r33_c6_12 = t_r33_c6_11 + p_34_7;
  assign out_33_6 = t_r33_c6_12 >> 4;

  assign t_r33_c7_0 = p_32_7 << 1;
  assign t_r33_c7_1 = p_33_6 << 1;
  assign t_r33_c7_2 = p_33_7 << 2;
  assign t_r33_c7_3 = p_33_8 << 1;
  assign t_r33_c7_4 = p_34_7 << 1;
  assign t_r33_c7_5 = t_r33_c7_0 + p_32_6;
  assign t_r33_c7_6 = t_r33_c7_1 + p_32_8;
  assign t_r33_c7_7 = t_r33_c7_2 + t_r33_c7_3;
  assign t_r33_c7_8 = t_r33_c7_4 + p_34_6;
  assign t_r33_c7_9 = t_r33_c7_5 + t_r33_c7_6;
  assign t_r33_c7_10 = t_r33_c7_7 + t_r33_c7_8;
  assign t_r33_c7_11 = t_r33_c7_9 + t_r33_c7_10;
  assign t_r33_c7_12 = t_r33_c7_11 + p_34_8;
  assign out_33_7 = t_r33_c7_12 >> 4;

  assign t_r33_c8_0 = p_32_8 << 1;
  assign t_r33_c8_1 = p_33_7 << 1;
  assign t_r33_c8_2 = p_33_8 << 2;
  assign t_r33_c8_3 = p_33_9 << 1;
  assign t_r33_c8_4 = p_34_8 << 1;
  assign t_r33_c8_5 = t_r33_c8_0 + p_32_7;
  assign t_r33_c8_6 = t_r33_c8_1 + p_32_9;
  assign t_r33_c8_7 = t_r33_c8_2 + t_r33_c8_3;
  assign t_r33_c8_8 = t_r33_c8_4 + p_34_7;
  assign t_r33_c8_9 = t_r33_c8_5 + t_r33_c8_6;
  assign t_r33_c8_10 = t_r33_c8_7 + t_r33_c8_8;
  assign t_r33_c8_11 = t_r33_c8_9 + t_r33_c8_10;
  assign t_r33_c8_12 = t_r33_c8_11 + p_34_9;
  assign out_33_8 = t_r33_c8_12 >> 4;

  assign t_r33_c9_0 = p_32_9 << 1;
  assign t_r33_c9_1 = p_33_8 << 1;
  assign t_r33_c9_2 = p_33_9 << 2;
  assign t_r33_c9_3 = p_33_10 << 1;
  assign t_r33_c9_4 = p_34_9 << 1;
  assign t_r33_c9_5 = t_r33_c9_0 + p_32_8;
  assign t_r33_c9_6 = t_r33_c9_1 + p_32_10;
  assign t_r33_c9_7 = t_r33_c9_2 + t_r33_c9_3;
  assign t_r33_c9_8 = t_r33_c9_4 + p_34_8;
  assign t_r33_c9_9 = t_r33_c9_5 + t_r33_c9_6;
  assign t_r33_c9_10 = t_r33_c9_7 + t_r33_c9_8;
  assign t_r33_c9_11 = t_r33_c9_9 + t_r33_c9_10;
  assign t_r33_c9_12 = t_r33_c9_11 + p_34_10;
  assign out_33_9 = t_r33_c9_12 >> 4;

  assign t_r33_c10_0 = p_32_10 << 1;
  assign t_r33_c10_1 = p_33_9 << 1;
  assign t_r33_c10_2 = p_33_10 << 2;
  assign t_r33_c10_3 = p_33_11 << 1;
  assign t_r33_c10_4 = p_34_10 << 1;
  assign t_r33_c10_5 = t_r33_c10_0 + p_32_9;
  assign t_r33_c10_6 = t_r33_c10_1 + p_32_11;
  assign t_r33_c10_7 = t_r33_c10_2 + t_r33_c10_3;
  assign t_r33_c10_8 = t_r33_c10_4 + p_34_9;
  assign t_r33_c10_9 = t_r33_c10_5 + t_r33_c10_6;
  assign t_r33_c10_10 = t_r33_c10_7 + t_r33_c10_8;
  assign t_r33_c10_11 = t_r33_c10_9 + t_r33_c10_10;
  assign t_r33_c10_12 = t_r33_c10_11 + p_34_11;
  assign out_33_10 = t_r33_c10_12 >> 4;

  assign t_r33_c11_0 = p_32_11 << 1;
  assign t_r33_c11_1 = p_33_10 << 1;
  assign t_r33_c11_2 = p_33_11 << 2;
  assign t_r33_c11_3 = p_33_12 << 1;
  assign t_r33_c11_4 = p_34_11 << 1;
  assign t_r33_c11_5 = t_r33_c11_0 + p_32_10;
  assign t_r33_c11_6 = t_r33_c11_1 + p_32_12;
  assign t_r33_c11_7 = t_r33_c11_2 + t_r33_c11_3;
  assign t_r33_c11_8 = t_r33_c11_4 + p_34_10;
  assign t_r33_c11_9 = t_r33_c11_5 + t_r33_c11_6;
  assign t_r33_c11_10 = t_r33_c11_7 + t_r33_c11_8;
  assign t_r33_c11_11 = t_r33_c11_9 + t_r33_c11_10;
  assign t_r33_c11_12 = t_r33_c11_11 + p_34_12;
  assign out_33_11 = t_r33_c11_12 >> 4;

  assign t_r33_c12_0 = p_32_12 << 1;
  assign t_r33_c12_1 = p_33_11 << 1;
  assign t_r33_c12_2 = p_33_12 << 2;
  assign t_r33_c12_3 = p_33_13 << 1;
  assign t_r33_c12_4 = p_34_12 << 1;
  assign t_r33_c12_5 = t_r33_c12_0 + p_32_11;
  assign t_r33_c12_6 = t_r33_c12_1 + p_32_13;
  assign t_r33_c12_7 = t_r33_c12_2 + t_r33_c12_3;
  assign t_r33_c12_8 = t_r33_c12_4 + p_34_11;
  assign t_r33_c12_9 = t_r33_c12_5 + t_r33_c12_6;
  assign t_r33_c12_10 = t_r33_c12_7 + t_r33_c12_8;
  assign t_r33_c12_11 = t_r33_c12_9 + t_r33_c12_10;
  assign t_r33_c12_12 = t_r33_c12_11 + p_34_13;
  assign out_33_12 = t_r33_c12_12 >> 4;

  assign t_r33_c13_0 = p_32_13 << 1;
  assign t_r33_c13_1 = p_33_12 << 1;
  assign t_r33_c13_2 = p_33_13 << 2;
  assign t_r33_c13_3 = p_33_14 << 1;
  assign t_r33_c13_4 = p_34_13 << 1;
  assign t_r33_c13_5 = t_r33_c13_0 + p_32_12;
  assign t_r33_c13_6 = t_r33_c13_1 + p_32_14;
  assign t_r33_c13_7 = t_r33_c13_2 + t_r33_c13_3;
  assign t_r33_c13_8 = t_r33_c13_4 + p_34_12;
  assign t_r33_c13_9 = t_r33_c13_5 + t_r33_c13_6;
  assign t_r33_c13_10 = t_r33_c13_7 + t_r33_c13_8;
  assign t_r33_c13_11 = t_r33_c13_9 + t_r33_c13_10;
  assign t_r33_c13_12 = t_r33_c13_11 + p_34_14;
  assign out_33_13 = t_r33_c13_12 >> 4;

  assign t_r33_c14_0 = p_32_14 << 1;
  assign t_r33_c14_1 = p_33_13 << 1;
  assign t_r33_c14_2 = p_33_14 << 2;
  assign t_r33_c14_3 = p_33_15 << 1;
  assign t_r33_c14_4 = p_34_14 << 1;
  assign t_r33_c14_5 = t_r33_c14_0 + p_32_13;
  assign t_r33_c14_6 = t_r33_c14_1 + p_32_15;
  assign t_r33_c14_7 = t_r33_c14_2 + t_r33_c14_3;
  assign t_r33_c14_8 = t_r33_c14_4 + p_34_13;
  assign t_r33_c14_9 = t_r33_c14_5 + t_r33_c14_6;
  assign t_r33_c14_10 = t_r33_c14_7 + t_r33_c14_8;
  assign t_r33_c14_11 = t_r33_c14_9 + t_r33_c14_10;
  assign t_r33_c14_12 = t_r33_c14_11 + p_34_15;
  assign out_33_14 = t_r33_c14_12 >> 4;

  assign t_r33_c15_0 = p_32_15 << 1;
  assign t_r33_c15_1 = p_33_14 << 1;
  assign t_r33_c15_2 = p_33_15 << 2;
  assign t_r33_c15_3 = p_33_16 << 1;
  assign t_r33_c15_4 = p_34_15 << 1;
  assign t_r33_c15_5 = t_r33_c15_0 + p_32_14;
  assign t_r33_c15_6 = t_r33_c15_1 + p_32_16;
  assign t_r33_c15_7 = t_r33_c15_2 + t_r33_c15_3;
  assign t_r33_c15_8 = t_r33_c15_4 + p_34_14;
  assign t_r33_c15_9 = t_r33_c15_5 + t_r33_c15_6;
  assign t_r33_c15_10 = t_r33_c15_7 + t_r33_c15_8;
  assign t_r33_c15_11 = t_r33_c15_9 + t_r33_c15_10;
  assign t_r33_c15_12 = t_r33_c15_11 + p_34_16;
  assign out_33_15 = t_r33_c15_12 >> 4;

  assign t_r33_c16_0 = p_32_16 << 1;
  assign t_r33_c16_1 = p_33_15 << 1;
  assign t_r33_c16_2 = p_33_16 << 2;
  assign t_r33_c16_3 = p_33_17 << 1;
  assign t_r33_c16_4 = p_34_16 << 1;
  assign t_r33_c16_5 = t_r33_c16_0 + p_32_15;
  assign t_r33_c16_6 = t_r33_c16_1 + p_32_17;
  assign t_r33_c16_7 = t_r33_c16_2 + t_r33_c16_3;
  assign t_r33_c16_8 = t_r33_c16_4 + p_34_15;
  assign t_r33_c16_9 = t_r33_c16_5 + t_r33_c16_6;
  assign t_r33_c16_10 = t_r33_c16_7 + t_r33_c16_8;
  assign t_r33_c16_11 = t_r33_c16_9 + t_r33_c16_10;
  assign t_r33_c16_12 = t_r33_c16_11 + p_34_17;
  assign out_33_16 = t_r33_c16_12 >> 4;

  assign t_r33_c17_0 = p_32_17 << 1;
  assign t_r33_c17_1 = p_33_16 << 1;
  assign t_r33_c17_2 = p_33_17 << 2;
  assign t_r33_c17_3 = p_33_18 << 1;
  assign t_r33_c17_4 = p_34_17 << 1;
  assign t_r33_c17_5 = t_r33_c17_0 + p_32_16;
  assign t_r33_c17_6 = t_r33_c17_1 + p_32_18;
  assign t_r33_c17_7 = t_r33_c17_2 + t_r33_c17_3;
  assign t_r33_c17_8 = t_r33_c17_4 + p_34_16;
  assign t_r33_c17_9 = t_r33_c17_5 + t_r33_c17_6;
  assign t_r33_c17_10 = t_r33_c17_7 + t_r33_c17_8;
  assign t_r33_c17_11 = t_r33_c17_9 + t_r33_c17_10;
  assign t_r33_c17_12 = t_r33_c17_11 + p_34_18;
  assign out_33_17 = t_r33_c17_12 >> 4;

  assign t_r33_c18_0 = p_32_18 << 1;
  assign t_r33_c18_1 = p_33_17 << 1;
  assign t_r33_c18_2 = p_33_18 << 2;
  assign t_r33_c18_3 = p_33_19 << 1;
  assign t_r33_c18_4 = p_34_18 << 1;
  assign t_r33_c18_5 = t_r33_c18_0 + p_32_17;
  assign t_r33_c18_6 = t_r33_c18_1 + p_32_19;
  assign t_r33_c18_7 = t_r33_c18_2 + t_r33_c18_3;
  assign t_r33_c18_8 = t_r33_c18_4 + p_34_17;
  assign t_r33_c18_9 = t_r33_c18_5 + t_r33_c18_6;
  assign t_r33_c18_10 = t_r33_c18_7 + t_r33_c18_8;
  assign t_r33_c18_11 = t_r33_c18_9 + t_r33_c18_10;
  assign t_r33_c18_12 = t_r33_c18_11 + p_34_19;
  assign out_33_18 = t_r33_c18_12 >> 4;

  assign t_r33_c19_0 = p_32_19 << 1;
  assign t_r33_c19_1 = p_33_18 << 1;
  assign t_r33_c19_2 = p_33_19 << 2;
  assign t_r33_c19_3 = p_33_20 << 1;
  assign t_r33_c19_4 = p_34_19 << 1;
  assign t_r33_c19_5 = t_r33_c19_0 + p_32_18;
  assign t_r33_c19_6 = t_r33_c19_1 + p_32_20;
  assign t_r33_c19_7 = t_r33_c19_2 + t_r33_c19_3;
  assign t_r33_c19_8 = t_r33_c19_4 + p_34_18;
  assign t_r33_c19_9 = t_r33_c19_5 + t_r33_c19_6;
  assign t_r33_c19_10 = t_r33_c19_7 + t_r33_c19_8;
  assign t_r33_c19_11 = t_r33_c19_9 + t_r33_c19_10;
  assign t_r33_c19_12 = t_r33_c19_11 + p_34_20;
  assign out_33_19 = t_r33_c19_12 >> 4;

  assign t_r33_c20_0 = p_32_20 << 1;
  assign t_r33_c20_1 = p_33_19 << 1;
  assign t_r33_c20_2 = p_33_20 << 2;
  assign t_r33_c20_3 = p_33_21 << 1;
  assign t_r33_c20_4 = p_34_20 << 1;
  assign t_r33_c20_5 = t_r33_c20_0 + p_32_19;
  assign t_r33_c20_6 = t_r33_c20_1 + p_32_21;
  assign t_r33_c20_7 = t_r33_c20_2 + t_r33_c20_3;
  assign t_r33_c20_8 = t_r33_c20_4 + p_34_19;
  assign t_r33_c20_9 = t_r33_c20_5 + t_r33_c20_6;
  assign t_r33_c20_10 = t_r33_c20_7 + t_r33_c20_8;
  assign t_r33_c20_11 = t_r33_c20_9 + t_r33_c20_10;
  assign t_r33_c20_12 = t_r33_c20_11 + p_34_21;
  assign out_33_20 = t_r33_c20_12 >> 4;

  assign t_r33_c21_0 = p_32_21 << 1;
  assign t_r33_c21_1 = p_33_20 << 1;
  assign t_r33_c21_2 = p_33_21 << 2;
  assign t_r33_c21_3 = p_33_22 << 1;
  assign t_r33_c21_4 = p_34_21 << 1;
  assign t_r33_c21_5 = t_r33_c21_0 + p_32_20;
  assign t_r33_c21_6 = t_r33_c21_1 + p_32_22;
  assign t_r33_c21_7 = t_r33_c21_2 + t_r33_c21_3;
  assign t_r33_c21_8 = t_r33_c21_4 + p_34_20;
  assign t_r33_c21_9 = t_r33_c21_5 + t_r33_c21_6;
  assign t_r33_c21_10 = t_r33_c21_7 + t_r33_c21_8;
  assign t_r33_c21_11 = t_r33_c21_9 + t_r33_c21_10;
  assign t_r33_c21_12 = t_r33_c21_11 + p_34_22;
  assign out_33_21 = t_r33_c21_12 >> 4;

  assign t_r33_c22_0 = p_32_22 << 1;
  assign t_r33_c22_1 = p_33_21 << 1;
  assign t_r33_c22_2 = p_33_22 << 2;
  assign t_r33_c22_3 = p_33_23 << 1;
  assign t_r33_c22_4 = p_34_22 << 1;
  assign t_r33_c22_5 = t_r33_c22_0 + p_32_21;
  assign t_r33_c22_6 = t_r33_c22_1 + p_32_23;
  assign t_r33_c22_7 = t_r33_c22_2 + t_r33_c22_3;
  assign t_r33_c22_8 = t_r33_c22_4 + p_34_21;
  assign t_r33_c22_9 = t_r33_c22_5 + t_r33_c22_6;
  assign t_r33_c22_10 = t_r33_c22_7 + t_r33_c22_8;
  assign t_r33_c22_11 = t_r33_c22_9 + t_r33_c22_10;
  assign t_r33_c22_12 = t_r33_c22_11 + p_34_23;
  assign out_33_22 = t_r33_c22_12 >> 4;

  assign t_r33_c23_0 = p_32_23 << 1;
  assign t_r33_c23_1 = p_33_22 << 1;
  assign t_r33_c23_2 = p_33_23 << 2;
  assign t_r33_c23_3 = p_33_24 << 1;
  assign t_r33_c23_4 = p_34_23 << 1;
  assign t_r33_c23_5 = t_r33_c23_0 + p_32_22;
  assign t_r33_c23_6 = t_r33_c23_1 + p_32_24;
  assign t_r33_c23_7 = t_r33_c23_2 + t_r33_c23_3;
  assign t_r33_c23_8 = t_r33_c23_4 + p_34_22;
  assign t_r33_c23_9 = t_r33_c23_5 + t_r33_c23_6;
  assign t_r33_c23_10 = t_r33_c23_7 + t_r33_c23_8;
  assign t_r33_c23_11 = t_r33_c23_9 + t_r33_c23_10;
  assign t_r33_c23_12 = t_r33_c23_11 + p_34_24;
  assign out_33_23 = t_r33_c23_12 >> 4;

  assign t_r33_c24_0 = p_32_24 << 1;
  assign t_r33_c24_1 = p_33_23 << 1;
  assign t_r33_c24_2 = p_33_24 << 2;
  assign t_r33_c24_3 = p_33_25 << 1;
  assign t_r33_c24_4 = p_34_24 << 1;
  assign t_r33_c24_5 = t_r33_c24_0 + p_32_23;
  assign t_r33_c24_6 = t_r33_c24_1 + p_32_25;
  assign t_r33_c24_7 = t_r33_c24_2 + t_r33_c24_3;
  assign t_r33_c24_8 = t_r33_c24_4 + p_34_23;
  assign t_r33_c24_9 = t_r33_c24_5 + t_r33_c24_6;
  assign t_r33_c24_10 = t_r33_c24_7 + t_r33_c24_8;
  assign t_r33_c24_11 = t_r33_c24_9 + t_r33_c24_10;
  assign t_r33_c24_12 = t_r33_c24_11 + p_34_25;
  assign out_33_24 = t_r33_c24_12 >> 4;

  assign t_r33_c25_0 = p_32_25 << 1;
  assign t_r33_c25_1 = p_33_24 << 1;
  assign t_r33_c25_2 = p_33_25 << 2;
  assign t_r33_c25_3 = p_33_26 << 1;
  assign t_r33_c25_4 = p_34_25 << 1;
  assign t_r33_c25_5 = t_r33_c25_0 + p_32_24;
  assign t_r33_c25_6 = t_r33_c25_1 + p_32_26;
  assign t_r33_c25_7 = t_r33_c25_2 + t_r33_c25_3;
  assign t_r33_c25_8 = t_r33_c25_4 + p_34_24;
  assign t_r33_c25_9 = t_r33_c25_5 + t_r33_c25_6;
  assign t_r33_c25_10 = t_r33_c25_7 + t_r33_c25_8;
  assign t_r33_c25_11 = t_r33_c25_9 + t_r33_c25_10;
  assign t_r33_c25_12 = t_r33_c25_11 + p_34_26;
  assign out_33_25 = t_r33_c25_12 >> 4;

  assign t_r33_c26_0 = p_32_26 << 1;
  assign t_r33_c26_1 = p_33_25 << 1;
  assign t_r33_c26_2 = p_33_26 << 2;
  assign t_r33_c26_3 = p_33_27 << 1;
  assign t_r33_c26_4 = p_34_26 << 1;
  assign t_r33_c26_5 = t_r33_c26_0 + p_32_25;
  assign t_r33_c26_6 = t_r33_c26_1 + p_32_27;
  assign t_r33_c26_7 = t_r33_c26_2 + t_r33_c26_3;
  assign t_r33_c26_8 = t_r33_c26_4 + p_34_25;
  assign t_r33_c26_9 = t_r33_c26_5 + t_r33_c26_6;
  assign t_r33_c26_10 = t_r33_c26_7 + t_r33_c26_8;
  assign t_r33_c26_11 = t_r33_c26_9 + t_r33_c26_10;
  assign t_r33_c26_12 = t_r33_c26_11 + p_34_27;
  assign out_33_26 = t_r33_c26_12 >> 4;

  assign t_r33_c27_0 = p_32_27 << 1;
  assign t_r33_c27_1 = p_33_26 << 1;
  assign t_r33_c27_2 = p_33_27 << 2;
  assign t_r33_c27_3 = p_33_28 << 1;
  assign t_r33_c27_4 = p_34_27 << 1;
  assign t_r33_c27_5 = t_r33_c27_0 + p_32_26;
  assign t_r33_c27_6 = t_r33_c27_1 + p_32_28;
  assign t_r33_c27_7 = t_r33_c27_2 + t_r33_c27_3;
  assign t_r33_c27_8 = t_r33_c27_4 + p_34_26;
  assign t_r33_c27_9 = t_r33_c27_5 + t_r33_c27_6;
  assign t_r33_c27_10 = t_r33_c27_7 + t_r33_c27_8;
  assign t_r33_c27_11 = t_r33_c27_9 + t_r33_c27_10;
  assign t_r33_c27_12 = t_r33_c27_11 + p_34_28;
  assign out_33_27 = t_r33_c27_12 >> 4;

  assign t_r33_c28_0 = p_32_28 << 1;
  assign t_r33_c28_1 = p_33_27 << 1;
  assign t_r33_c28_2 = p_33_28 << 2;
  assign t_r33_c28_3 = p_33_29 << 1;
  assign t_r33_c28_4 = p_34_28 << 1;
  assign t_r33_c28_5 = t_r33_c28_0 + p_32_27;
  assign t_r33_c28_6 = t_r33_c28_1 + p_32_29;
  assign t_r33_c28_7 = t_r33_c28_2 + t_r33_c28_3;
  assign t_r33_c28_8 = t_r33_c28_4 + p_34_27;
  assign t_r33_c28_9 = t_r33_c28_5 + t_r33_c28_6;
  assign t_r33_c28_10 = t_r33_c28_7 + t_r33_c28_8;
  assign t_r33_c28_11 = t_r33_c28_9 + t_r33_c28_10;
  assign t_r33_c28_12 = t_r33_c28_11 + p_34_29;
  assign out_33_28 = t_r33_c28_12 >> 4;

  assign t_r33_c29_0 = p_32_29 << 1;
  assign t_r33_c29_1 = p_33_28 << 1;
  assign t_r33_c29_2 = p_33_29 << 2;
  assign t_r33_c29_3 = p_33_30 << 1;
  assign t_r33_c29_4 = p_34_29 << 1;
  assign t_r33_c29_5 = t_r33_c29_0 + p_32_28;
  assign t_r33_c29_6 = t_r33_c29_1 + p_32_30;
  assign t_r33_c29_7 = t_r33_c29_2 + t_r33_c29_3;
  assign t_r33_c29_8 = t_r33_c29_4 + p_34_28;
  assign t_r33_c29_9 = t_r33_c29_5 + t_r33_c29_6;
  assign t_r33_c29_10 = t_r33_c29_7 + t_r33_c29_8;
  assign t_r33_c29_11 = t_r33_c29_9 + t_r33_c29_10;
  assign t_r33_c29_12 = t_r33_c29_11 + p_34_30;
  assign out_33_29 = t_r33_c29_12 >> 4;

  assign t_r33_c30_0 = p_32_30 << 1;
  assign t_r33_c30_1 = p_33_29 << 1;
  assign t_r33_c30_2 = p_33_30 << 2;
  assign t_r33_c30_3 = p_33_31 << 1;
  assign t_r33_c30_4 = p_34_30 << 1;
  assign t_r33_c30_5 = t_r33_c30_0 + p_32_29;
  assign t_r33_c30_6 = t_r33_c30_1 + p_32_31;
  assign t_r33_c30_7 = t_r33_c30_2 + t_r33_c30_3;
  assign t_r33_c30_8 = t_r33_c30_4 + p_34_29;
  assign t_r33_c30_9 = t_r33_c30_5 + t_r33_c30_6;
  assign t_r33_c30_10 = t_r33_c30_7 + t_r33_c30_8;
  assign t_r33_c30_11 = t_r33_c30_9 + t_r33_c30_10;
  assign t_r33_c30_12 = t_r33_c30_11 + p_34_31;
  assign out_33_30 = t_r33_c30_12 >> 4;

  assign t_r33_c31_0 = p_32_31 << 1;
  assign t_r33_c31_1 = p_33_30 << 1;
  assign t_r33_c31_2 = p_33_31 << 2;
  assign t_r33_c31_3 = p_33_32 << 1;
  assign t_r33_c31_4 = p_34_31 << 1;
  assign t_r33_c31_5 = t_r33_c31_0 + p_32_30;
  assign t_r33_c31_6 = t_r33_c31_1 + p_32_32;
  assign t_r33_c31_7 = t_r33_c31_2 + t_r33_c31_3;
  assign t_r33_c31_8 = t_r33_c31_4 + p_34_30;
  assign t_r33_c31_9 = t_r33_c31_5 + t_r33_c31_6;
  assign t_r33_c31_10 = t_r33_c31_7 + t_r33_c31_8;
  assign t_r33_c31_11 = t_r33_c31_9 + t_r33_c31_10;
  assign t_r33_c31_12 = t_r33_c31_11 + p_34_32;
  assign out_33_31 = t_r33_c31_12 >> 4;

  assign t_r33_c32_0 = p_32_32 << 1;
  assign t_r33_c32_1 = p_33_31 << 1;
  assign t_r33_c32_2 = p_33_32 << 2;
  assign t_r33_c32_3 = p_33_33 << 1;
  assign t_r33_c32_4 = p_34_32 << 1;
  assign t_r33_c32_5 = t_r33_c32_0 + p_32_31;
  assign t_r33_c32_6 = t_r33_c32_1 + p_32_33;
  assign t_r33_c32_7 = t_r33_c32_2 + t_r33_c32_3;
  assign t_r33_c32_8 = t_r33_c32_4 + p_34_31;
  assign t_r33_c32_9 = t_r33_c32_5 + t_r33_c32_6;
  assign t_r33_c32_10 = t_r33_c32_7 + t_r33_c32_8;
  assign t_r33_c32_11 = t_r33_c32_9 + t_r33_c32_10;
  assign t_r33_c32_12 = t_r33_c32_11 + p_34_33;
  assign out_33_32 = t_r33_c32_12 >> 4;

  assign t_r33_c33_0 = p_32_33 << 1;
  assign t_r33_c33_1 = p_33_32 << 1;
  assign t_r33_c33_2 = p_33_33 << 2;
  assign t_r33_c33_3 = p_33_34 << 1;
  assign t_r33_c33_4 = p_34_33 << 1;
  assign t_r33_c33_5 = t_r33_c33_0 + p_32_32;
  assign t_r33_c33_6 = t_r33_c33_1 + p_32_34;
  assign t_r33_c33_7 = t_r33_c33_2 + t_r33_c33_3;
  assign t_r33_c33_8 = t_r33_c33_4 + p_34_32;
  assign t_r33_c33_9 = t_r33_c33_5 + t_r33_c33_6;
  assign t_r33_c33_10 = t_r33_c33_7 + t_r33_c33_8;
  assign t_r33_c33_11 = t_r33_c33_9 + t_r33_c33_10;
  assign t_r33_c33_12 = t_r33_c33_11 + p_34_34;
  assign out_33_33 = t_r33_c33_12 >> 4;

  assign t_r33_c34_0 = p_32_34 << 1;
  assign t_r33_c34_1 = p_33_33 << 1;
  assign t_r33_c34_2 = p_33_34 << 2;
  assign t_r33_c34_3 = p_33_35 << 1;
  assign t_r33_c34_4 = p_34_34 << 1;
  assign t_r33_c34_5 = t_r33_c34_0 + p_32_33;
  assign t_r33_c34_6 = t_r33_c34_1 + p_32_35;
  assign t_r33_c34_7 = t_r33_c34_2 + t_r33_c34_3;
  assign t_r33_c34_8 = t_r33_c34_4 + p_34_33;
  assign t_r33_c34_9 = t_r33_c34_5 + t_r33_c34_6;
  assign t_r33_c34_10 = t_r33_c34_7 + t_r33_c34_8;
  assign t_r33_c34_11 = t_r33_c34_9 + t_r33_c34_10;
  assign t_r33_c34_12 = t_r33_c34_11 + p_34_35;
  assign out_33_34 = t_r33_c34_12 >> 4;

  assign t_r33_c35_0 = p_32_35 << 1;
  assign t_r33_c35_1 = p_33_34 << 1;
  assign t_r33_c35_2 = p_33_35 << 2;
  assign t_r33_c35_3 = p_33_36 << 1;
  assign t_r33_c35_4 = p_34_35 << 1;
  assign t_r33_c35_5 = t_r33_c35_0 + p_32_34;
  assign t_r33_c35_6 = t_r33_c35_1 + p_32_36;
  assign t_r33_c35_7 = t_r33_c35_2 + t_r33_c35_3;
  assign t_r33_c35_8 = t_r33_c35_4 + p_34_34;
  assign t_r33_c35_9 = t_r33_c35_5 + t_r33_c35_6;
  assign t_r33_c35_10 = t_r33_c35_7 + t_r33_c35_8;
  assign t_r33_c35_11 = t_r33_c35_9 + t_r33_c35_10;
  assign t_r33_c35_12 = t_r33_c35_11 + p_34_36;
  assign out_33_35 = t_r33_c35_12 >> 4;

  assign t_r33_c36_0 = p_32_36 << 1;
  assign t_r33_c36_1 = p_33_35 << 1;
  assign t_r33_c36_2 = p_33_36 << 2;
  assign t_r33_c36_3 = p_33_37 << 1;
  assign t_r33_c36_4 = p_34_36 << 1;
  assign t_r33_c36_5 = t_r33_c36_0 + p_32_35;
  assign t_r33_c36_6 = t_r33_c36_1 + p_32_37;
  assign t_r33_c36_7 = t_r33_c36_2 + t_r33_c36_3;
  assign t_r33_c36_8 = t_r33_c36_4 + p_34_35;
  assign t_r33_c36_9 = t_r33_c36_5 + t_r33_c36_6;
  assign t_r33_c36_10 = t_r33_c36_7 + t_r33_c36_8;
  assign t_r33_c36_11 = t_r33_c36_9 + t_r33_c36_10;
  assign t_r33_c36_12 = t_r33_c36_11 + p_34_37;
  assign out_33_36 = t_r33_c36_12 >> 4;

  assign t_r33_c37_0 = p_32_37 << 1;
  assign t_r33_c37_1 = p_33_36 << 1;
  assign t_r33_c37_2 = p_33_37 << 2;
  assign t_r33_c37_3 = p_33_38 << 1;
  assign t_r33_c37_4 = p_34_37 << 1;
  assign t_r33_c37_5 = t_r33_c37_0 + p_32_36;
  assign t_r33_c37_6 = t_r33_c37_1 + p_32_38;
  assign t_r33_c37_7 = t_r33_c37_2 + t_r33_c37_3;
  assign t_r33_c37_8 = t_r33_c37_4 + p_34_36;
  assign t_r33_c37_9 = t_r33_c37_5 + t_r33_c37_6;
  assign t_r33_c37_10 = t_r33_c37_7 + t_r33_c37_8;
  assign t_r33_c37_11 = t_r33_c37_9 + t_r33_c37_10;
  assign t_r33_c37_12 = t_r33_c37_11 + p_34_38;
  assign out_33_37 = t_r33_c37_12 >> 4;

  assign t_r33_c38_0 = p_32_38 << 1;
  assign t_r33_c38_1 = p_33_37 << 1;
  assign t_r33_c38_2 = p_33_38 << 2;
  assign t_r33_c38_3 = p_33_39 << 1;
  assign t_r33_c38_4 = p_34_38 << 1;
  assign t_r33_c38_5 = t_r33_c38_0 + p_32_37;
  assign t_r33_c38_6 = t_r33_c38_1 + p_32_39;
  assign t_r33_c38_7 = t_r33_c38_2 + t_r33_c38_3;
  assign t_r33_c38_8 = t_r33_c38_4 + p_34_37;
  assign t_r33_c38_9 = t_r33_c38_5 + t_r33_c38_6;
  assign t_r33_c38_10 = t_r33_c38_7 + t_r33_c38_8;
  assign t_r33_c38_11 = t_r33_c38_9 + t_r33_c38_10;
  assign t_r33_c38_12 = t_r33_c38_11 + p_34_39;
  assign out_33_38 = t_r33_c38_12 >> 4;

  assign t_r33_c39_0 = p_32_39 << 1;
  assign t_r33_c39_1 = p_33_38 << 1;
  assign t_r33_c39_2 = p_33_39 << 2;
  assign t_r33_c39_3 = p_33_40 << 1;
  assign t_r33_c39_4 = p_34_39 << 1;
  assign t_r33_c39_5 = t_r33_c39_0 + p_32_38;
  assign t_r33_c39_6 = t_r33_c39_1 + p_32_40;
  assign t_r33_c39_7 = t_r33_c39_2 + t_r33_c39_3;
  assign t_r33_c39_8 = t_r33_c39_4 + p_34_38;
  assign t_r33_c39_9 = t_r33_c39_5 + t_r33_c39_6;
  assign t_r33_c39_10 = t_r33_c39_7 + t_r33_c39_8;
  assign t_r33_c39_11 = t_r33_c39_9 + t_r33_c39_10;
  assign t_r33_c39_12 = t_r33_c39_11 + p_34_40;
  assign out_33_39 = t_r33_c39_12 >> 4;

  assign t_r33_c40_0 = p_32_40 << 1;
  assign t_r33_c40_1 = p_33_39 << 1;
  assign t_r33_c40_2 = p_33_40 << 2;
  assign t_r33_c40_3 = p_33_41 << 1;
  assign t_r33_c40_4 = p_34_40 << 1;
  assign t_r33_c40_5 = t_r33_c40_0 + p_32_39;
  assign t_r33_c40_6 = t_r33_c40_1 + p_32_41;
  assign t_r33_c40_7 = t_r33_c40_2 + t_r33_c40_3;
  assign t_r33_c40_8 = t_r33_c40_4 + p_34_39;
  assign t_r33_c40_9 = t_r33_c40_5 + t_r33_c40_6;
  assign t_r33_c40_10 = t_r33_c40_7 + t_r33_c40_8;
  assign t_r33_c40_11 = t_r33_c40_9 + t_r33_c40_10;
  assign t_r33_c40_12 = t_r33_c40_11 + p_34_41;
  assign out_33_40 = t_r33_c40_12 >> 4;

  assign t_r33_c41_0 = p_32_41 << 1;
  assign t_r33_c41_1 = p_33_40 << 1;
  assign t_r33_c41_2 = p_33_41 << 2;
  assign t_r33_c41_3 = p_33_42 << 1;
  assign t_r33_c41_4 = p_34_41 << 1;
  assign t_r33_c41_5 = t_r33_c41_0 + p_32_40;
  assign t_r33_c41_6 = t_r33_c41_1 + p_32_42;
  assign t_r33_c41_7 = t_r33_c41_2 + t_r33_c41_3;
  assign t_r33_c41_8 = t_r33_c41_4 + p_34_40;
  assign t_r33_c41_9 = t_r33_c41_5 + t_r33_c41_6;
  assign t_r33_c41_10 = t_r33_c41_7 + t_r33_c41_8;
  assign t_r33_c41_11 = t_r33_c41_9 + t_r33_c41_10;
  assign t_r33_c41_12 = t_r33_c41_11 + p_34_42;
  assign out_33_41 = t_r33_c41_12 >> 4;

  assign t_r33_c42_0 = p_32_42 << 1;
  assign t_r33_c42_1 = p_33_41 << 1;
  assign t_r33_c42_2 = p_33_42 << 2;
  assign t_r33_c42_3 = p_33_43 << 1;
  assign t_r33_c42_4 = p_34_42 << 1;
  assign t_r33_c42_5 = t_r33_c42_0 + p_32_41;
  assign t_r33_c42_6 = t_r33_c42_1 + p_32_43;
  assign t_r33_c42_7 = t_r33_c42_2 + t_r33_c42_3;
  assign t_r33_c42_8 = t_r33_c42_4 + p_34_41;
  assign t_r33_c42_9 = t_r33_c42_5 + t_r33_c42_6;
  assign t_r33_c42_10 = t_r33_c42_7 + t_r33_c42_8;
  assign t_r33_c42_11 = t_r33_c42_9 + t_r33_c42_10;
  assign t_r33_c42_12 = t_r33_c42_11 + p_34_43;
  assign out_33_42 = t_r33_c42_12 >> 4;

  assign t_r33_c43_0 = p_32_43 << 1;
  assign t_r33_c43_1 = p_33_42 << 1;
  assign t_r33_c43_2 = p_33_43 << 2;
  assign t_r33_c43_3 = p_33_44 << 1;
  assign t_r33_c43_4 = p_34_43 << 1;
  assign t_r33_c43_5 = t_r33_c43_0 + p_32_42;
  assign t_r33_c43_6 = t_r33_c43_1 + p_32_44;
  assign t_r33_c43_7 = t_r33_c43_2 + t_r33_c43_3;
  assign t_r33_c43_8 = t_r33_c43_4 + p_34_42;
  assign t_r33_c43_9 = t_r33_c43_5 + t_r33_c43_6;
  assign t_r33_c43_10 = t_r33_c43_7 + t_r33_c43_8;
  assign t_r33_c43_11 = t_r33_c43_9 + t_r33_c43_10;
  assign t_r33_c43_12 = t_r33_c43_11 + p_34_44;
  assign out_33_43 = t_r33_c43_12 >> 4;

  assign t_r33_c44_0 = p_32_44 << 1;
  assign t_r33_c44_1 = p_33_43 << 1;
  assign t_r33_c44_2 = p_33_44 << 2;
  assign t_r33_c44_3 = p_33_45 << 1;
  assign t_r33_c44_4 = p_34_44 << 1;
  assign t_r33_c44_5 = t_r33_c44_0 + p_32_43;
  assign t_r33_c44_6 = t_r33_c44_1 + p_32_45;
  assign t_r33_c44_7 = t_r33_c44_2 + t_r33_c44_3;
  assign t_r33_c44_8 = t_r33_c44_4 + p_34_43;
  assign t_r33_c44_9 = t_r33_c44_5 + t_r33_c44_6;
  assign t_r33_c44_10 = t_r33_c44_7 + t_r33_c44_8;
  assign t_r33_c44_11 = t_r33_c44_9 + t_r33_c44_10;
  assign t_r33_c44_12 = t_r33_c44_11 + p_34_45;
  assign out_33_44 = t_r33_c44_12 >> 4;

  assign t_r33_c45_0 = p_32_45 << 1;
  assign t_r33_c45_1 = p_33_44 << 1;
  assign t_r33_c45_2 = p_33_45 << 2;
  assign t_r33_c45_3 = p_33_46 << 1;
  assign t_r33_c45_4 = p_34_45 << 1;
  assign t_r33_c45_5 = t_r33_c45_0 + p_32_44;
  assign t_r33_c45_6 = t_r33_c45_1 + p_32_46;
  assign t_r33_c45_7 = t_r33_c45_2 + t_r33_c45_3;
  assign t_r33_c45_8 = t_r33_c45_4 + p_34_44;
  assign t_r33_c45_9 = t_r33_c45_5 + t_r33_c45_6;
  assign t_r33_c45_10 = t_r33_c45_7 + t_r33_c45_8;
  assign t_r33_c45_11 = t_r33_c45_9 + t_r33_c45_10;
  assign t_r33_c45_12 = t_r33_c45_11 + p_34_46;
  assign out_33_45 = t_r33_c45_12 >> 4;

  assign t_r33_c46_0 = p_32_46 << 1;
  assign t_r33_c46_1 = p_33_45 << 1;
  assign t_r33_c46_2 = p_33_46 << 2;
  assign t_r33_c46_3 = p_33_47 << 1;
  assign t_r33_c46_4 = p_34_46 << 1;
  assign t_r33_c46_5 = t_r33_c46_0 + p_32_45;
  assign t_r33_c46_6 = t_r33_c46_1 + p_32_47;
  assign t_r33_c46_7 = t_r33_c46_2 + t_r33_c46_3;
  assign t_r33_c46_8 = t_r33_c46_4 + p_34_45;
  assign t_r33_c46_9 = t_r33_c46_5 + t_r33_c46_6;
  assign t_r33_c46_10 = t_r33_c46_7 + t_r33_c46_8;
  assign t_r33_c46_11 = t_r33_c46_9 + t_r33_c46_10;
  assign t_r33_c46_12 = t_r33_c46_11 + p_34_47;
  assign out_33_46 = t_r33_c46_12 >> 4;

  assign t_r33_c47_0 = p_32_47 << 1;
  assign t_r33_c47_1 = p_33_46 << 1;
  assign t_r33_c47_2 = p_33_47 << 2;
  assign t_r33_c47_3 = p_33_48 << 1;
  assign t_r33_c47_4 = p_34_47 << 1;
  assign t_r33_c47_5 = t_r33_c47_0 + p_32_46;
  assign t_r33_c47_6 = t_r33_c47_1 + p_32_48;
  assign t_r33_c47_7 = t_r33_c47_2 + t_r33_c47_3;
  assign t_r33_c47_8 = t_r33_c47_4 + p_34_46;
  assign t_r33_c47_9 = t_r33_c47_5 + t_r33_c47_6;
  assign t_r33_c47_10 = t_r33_c47_7 + t_r33_c47_8;
  assign t_r33_c47_11 = t_r33_c47_9 + t_r33_c47_10;
  assign t_r33_c47_12 = t_r33_c47_11 + p_34_48;
  assign out_33_47 = t_r33_c47_12 >> 4;

  assign t_r33_c48_0 = p_32_48 << 1;
  assign t_r33_c48_1 = p_33_47 << 1;
  assign t_r33_c48_2 = p_33_48 << 2;
  assign t_r33_c48_3 = p_33_49 << 1;
  assign t_r33_c48_4 = p_34_48 << 1;
  assign t_r33_c48_5 = t_r33_c48_0 + p_32_47;
  assign t_r33_c48_6 = t_r33_c48_1 + p_32_49;
  assign t_r33_c48_7 = t_r33_c48_2 + t_r33_c48_3;
  assign t_r33_c48_8 = t_r33_c48_4 + p_34_47;
  assign t_r33_c48_9 = t_r33_c48_5 + t_r33_c48_6;
  assign t_r33_c48_10 = t_r33_c48_7 + t_r33_c48_8;
  assign t_r33_c48_11 = t_r33_c48_9 + t_r33_c48_10;
  assign t_r33_c48_12 = t_r33_c48_11 + p_34_49;
  assign out_33_48 = t_r33_c48_12 >> 4;

  assign t_r33_c49_0 = p_32_49 << 1;
  assign t_r33_c49_1 = p_33_48 << 1;
  assign t_r33_c49_2 = p_33_49 << 2;
  assign t_r33_c49_3 = p_33_50 << 1;
  assign t_r33_c49_4 = p_34_49 << 1;
  assign t_r33_c49_5 = t_r33_c49_0 + p_32_48;
  assign t_r33_c49_6 = t_r33_c49_1 + p_32_50;
  assign t_r33_c49_7 = t_r33_c49_2 + t_r33_c49_3;
  assign t_r33_c49_8 = t_r33_c49_4 + p_34_48;
  assign t_r33_c49_9 = t_r33_c49_5 + t_r33_c49_6;
  assign t_r33_c49_10 = t_r33_c49_7 + t_r33_c49_8;
  assign t_r33_c49_11 = t_r33_c49_9 + t_r33_c49_10;
  assign t_r33_c49_12 = t_r33_c49_11 + p_34_50;
  assign out_33_49 = t_r33_c49_12 >> 4;

  assign t_r33_c50_0 = p_32_50 << 1;
  assign t_r33_c50_1 = p_33_49 << 1;
  assign t_r33_c50_2 = p_33_50 << 2;
  assign t_r33_c50_3 = p_33_51 << 1;
  assign t_r33_c50_4 = p_34_50 << 1;
  assign t_r33_c50_5 = t_r33_c50_0 + p_32_49;
  assign t_r33_c50_6 = t_r33_c50_1 + p_32_51;
  assign t_r33_c50_7 = t_r33_c50_2 + t_r33_c50_3;
  assign t_r33_c50_8 = t_r33_c50_4 + p_34_49;
  assign t_r33_c50_9 = t_r33_c50_5 + t_r33_c50_6;
  assign t_r33_c50_10 = t_r33_c50_7 + t_r33_c50_8;
  assign t_r33_c50_11 = t_r33_c50_9 + t_r33_c50_10;
  assign t_r33_c50_12 = t_r33_c50_11 + p_34_51;
  assign out_33_50 = t_r33_c50_12 >> 4;

  assign t_r33_c51_0 = p_32_51 << 1;
  assign t_r33_c51_1 = p_33_50 << 1;
  assign t_r33_c51_2 = p_33_51 << 2;
  assign t_r33_c51_3 = p_33_52 << 1;
  assign t_r33_c51_4 = p_34_51 << 1;
  assign t_r33_c51_5 = t_r33_c51_0 + p_32_50;
  assign t_r33_c51_6 = t_r33_c51_1 + p_32_52;
  assign t_r33_c51_7 = t_r33_c51_2 + t_r33_c51_3;
  assign t_r33_c51_8 = t_r33_c51_4 + p_34_50;
  assign t_r33_c51_9 = t_r33_c51_5 + t_r33_c51_6;
  assign t_r33_c51_10 = t_r33_c51_7 + t_r33_c51_8;
  assign t_r33_c51_11 = t_r33_c51_9 + t_r33_c51_10;
  assign t_r33_c51_12 = t_r33_c51_11 + p_34_52;
  assign out_33_51 = t_r33_c51_12 >> 4;

  assign t_r33_c52_0 = p_32_52 << 1;
  assign t_r33_c52_1 = p_33_51 << 1;
  assign t_r33_c52_2 = p_33_52 << 2;
  assign t_r33_c52_3 = p_33_53 << 1;
  assign t_r33_c52_4 = p_34_52 << 1;
  assign t_r33_c52_5 = t_r33_c52_0 + p_32_51;
  assign t_r33_c52_6 = t_r33_c52_1 + p_32_53;
  assign t_r33_c52_7 = t_r33_c52_2 + t_r33_c52_3;
  assign t_r33_c52_8 = t_r33_c52_4 + p_34_51;
  assign t_r33_c52_9 = t_r33_c52_5 + t_r33_c52_6;
  assign t_r33_c52_10 = t_r33_c52_7 + t_r33_c52_8;
  assign t_r33_c52_11 = t_r33_c52_9 + t_r33_c52_10;
  assign t_r33_c52_12 = t_r33_c52_11 + p_34_53;
  assign out_33_52 = t_r33_c52_12 >> 4;

  assign t_r33_c53_0 = p_32_53 << 1;
  assign t_r33_c53_1 = p_33_52 << 1;
  assign t_r33_c53_2 = p_33_53 << 2;
  assign t_r33_c53_3 = p_33_54 << 1;
  assign t_r33_c53_4 = p_34_53 << 1;
  assign t_r33_c53_5 = t_r33_c53_0 + p_32_52;
  assign t_r33_c53_6 = t_r33_c53_1 + p_32_54;
  assign t_r33_c53_7 = t_r33_c53_2 + t_r33_c53_3;
  assign t_r33_c53_8 = t_r33_c53_4 + p_34_52;
  assign t_r33_c53_9 = t_r33_c53_5 + t_r33_c53_6;
  assign t_r33_c53_10 = t_r33_c53_7 + t_r33_c53_8;
  assign t_r33_c53_11 = t_r33_c53_9 + t_r33_c53_10;
  assign t_r33_c53_12 = t_r33_c53_11 + p_34_54;
  assign out_33_53 = t_r33_c53_12 >> 4;

  assign t_r33_c54_0 = p_32_54 << 1;
  assign t_r33_c54_1 = p_33_53 << 1;
  assign t_r33_c54_2 = p_33_54 << 2;
  assign t_r33_c54_3 = p_33_55 << 1;
  assign t_r33_c54_4 = p_34_54 << 1;
  assign t_r33_c54_5 = t_r33_c54_0 + p_32_53;
  assign t_r33_c54_6 = t_r33_c54_1 + p_32_55;
  assign t_r33_c54_7 = t_r33_c54_2 + t_r33_c54_3;
  assign t_r33_c54_8 = t_r33_c54_4 + p_34_53;
  assign t_r33_c54_9 = t_r33_c54_5 + t_r33_c54_6;
  assign t_r33_c54_10 = t_r33_c54_7 + t_r33_c54_8;
  assign t_r33_c54_11 = t_r33_c54_9 + t_r33_c54_10;
  assign t_r33_c54_12 = t_r33_c54_11 + p_34_55;
  assign out_33_54 = t_r33_c54_12 >> 4;

  assign t_r33_c55_0 = p_32_55 << 1;
  assign t_r33_c55_1 = p_33_54 << 1;
  assign t_r33_c55_2 = p_33_55 << 2;
  assign t_r33_c55_3 = p_33_56 << 1;
  assign t_r33_c55_4 = p_34_55 << 1;
  assign t_r33_c55_5 = t_r33_c55_0 + p_32_54;
  assign t_r33_c55_6 = t_r33_c55_1 + p_32_56;
  assign t_r33_c55_7 = t_r33_c55_2 + t_r33_c55_3;
  assign t_r33_c55_8 = t_r33_c55_4 + p_34_54;
  assign t_r33_c55_9 = t_r33_c55_5 + t_r33_c55_6;
  assign t_r33_c55_10 = t_r33_c55_7 + t_r33_c55_8;
  assign t_r33_c55_11 = t_r33_c55_9 + t_r33_c55_10;
  assign t_r33_c55_12 = t_r33_c55_11 + p_34_56;
  assign out_33_55 = t_r33_c55_12 >> 4;

  assign t_r33_c56_0 = p_32_56 << 1;
  assign t_r33_c56_1 = p_33_55 << 1;
  assign t_r33_c56_2 = p_33_56 << 2;
  assign t_r33_c56_3 = p_33_57 << 1;
  assign t_r33_c56_4 = p_34_56 << 1;
  assign t_r33_c56_5 = t_r33_c56_0 + p_32_55;
  assign t_r33_c56_6 = t_r33_c56_1 + p_32_57;
  assign t_r33_c56_7 = t_r33_c56_2 + t_r33_c56_3;
  assign t_r33_c56_8 = t_r33_c56_4 + p_34_55;
  assign t_r33_c56_9 = t_r33_c56_5 + t_r33_c56_6;
  assign t_r33_c56_10 = t_r33_c56_7 + t_r33_c56_8;
  assign t_r33_c56_11 = t_r33_c56_9 + t_r33_c56_10;
  assign t_r33_c56_12 = t_r33_c56_11 + p_34_57;
  assign out_33_56 = t_r33_c56_12 >> 4;

  assign t_r33_c57_0 = p_32_57 << 1;
  assign t_r33_c57_1 = p_33_56 << 1;
  assign t_r33_c57_2 = p_33_57 << 2;
  assign t_r33_c57_3 = p_33_58 << 1;
  assign t_r33_c57_4 = p_34_57 << 1;
  assign t_r33_c57_5 = t_r33_c57_0 + p_32_56;
  assign t_r33_c57_6 = t_r33_c57_1 + p_32_58;
  assign t_r33_c57_7 = t_r33_c57_2 + t_r33_c57_3;
  assign t_r33_c57_8 = t_r33_c57_4 + p_34_56;
  assign t_r33_c57_9 = t_r33_c57_5 + t_r33_c57_6;
  assign t_r33_c57_10 = t_r33_c57_7 + t_r33_c57_8;
  assign t_r33_c57_11 = t_r33_c57_9 + t_r33_c57_10;
  assign t_r33_c57_12 = t_r33_c57_11 + p_34_58;
  assign out_33_57 = t_r33_c57_12 >> 4;

  assign t_r33_c58_0 = p_32_58 << 1;
  assign t_r33_c58_1 = p_33_57 << 1;
  assign t_r33_c58_2 = p_33_58 << 2;
  assign t_r33_c58_3 = p_33_59 << 1;
  assign t_r33_c58_4 = p_34_58 << 1;
  assign t_r33_c58_5 = t_r33_c58_0 + p_32_57;
  assign t_r33_c58_6 = t_r33_c58_1 + p_32_59;
  assign t_r33_c58_7 = t_r33_c58_2 + t_r33_c58_3;
  assign t_r33_c58_8 = t_r33_c58_4 + p_34_57;
  assign t_r33_c58_9 = t_r33_c58_5 + t_r33_c58_6;
  assign t_r33_c58_10 = t_r33_c58_7 + t_r33_c58_8;
  assign t_r33_c58_11 = t_r33_c58_9 + t_r33_c58_10;
  assign t_r33_c58_12 = t_r33_c58_11 + p_34_59;
  assign out_33_58 = t_r33_c58_12 >> 4;

  assign t_r33_c59_0 = p_32_59 << 1;
  assign t_r33_c59_1 = p_33_58 << 1;
  assign t_r33_c59_2 = p_33_59 << 2;
  assign t_r33_c59_3 = p_33_60 << 1;
  assign t_r33_c59_4 = p_34_59 << 1;
  assign t_r33_c59_5 = t_r33_c59_0 + p_32_58;
  assign t_r33_c59_6 = t_r33_c59_1 + p_32_60;
  assign t_r33_c59_7 = t_r33_c59_2 + t_r33_c59_3;
  assign t_r33_c59_8 = t_r33_c59_4 + p_34_58;
  assign t_r33_c59_9 = t_r33_c59_5 + t_r33_c59_6;
  assign t_r33_c59_10 = t_r33_c59_7 + t_r33_c59_8;
  assign t_r33_c59_11 = t_r33_c59_9 + t_r33_c59_10;
  assign t_r33_c59_12 = t_r33_c59_11 + p_34_60;
  assign out_33_59 = t_r33_c59_12 >> 4;

  assign t_r33_c60_0 = p_32_60 << 1;
  assign t_r33_c60_1 = p_33_59 << 1;
  assign t_r33_c60_2 = p_33_60 << 2;
  assign t_r33_c60_3 = p_33_61 << 1;
  assign t_r33_c60_4 = p_34_60 << 1;
  assign t_r33_c60_5 = t_r33_c60_0 + p_32_59;
  assign t_r33_c60_6 = t_r33_c60_1 + p_32_61;
  assign t_r33_c60_7 = t_r33_c60_2 + t_r33_c60_3;
  assign t_r33_c60_8 = t_r33_c60_4 + p_34_59;
  assign t_r33_c60_9 = t_r33_c60_5 + t_r33_c60_6;
  assign t_r33_c60_10 = t_r33_c60_7 + t_r33_c60_8;
  assign t_r33_c60_11 = t_r33_c60_9 + t_r33_c60_10;
  assign t_r33_c60_12 = t_r33_c60_11 + p_34_61;
  assign out_33_60 = t_r33_c60_12 >> 4;

  assign t_r33_c61_0 = p_32_61 << 1;
  assign t_r33_c61_1 = p_33_60 << 1;
  assign t_r33_c61_2 = p_33_61 << 2;
  assign t_r33_c61_3 = p_33_62 << 1;
  assign t_r33_c61_4 = p_34_61 << 1;
  assign t_r33_c61_5 = t_r33_c61_0 + p_32_60;
  assign t_r33_c61_6 = t_r33_c61_1 + p_32_62;
  assign t_r33_c61_7 = t_r33_c61_2 + t_r33_c61_3;
  assign t_r33_c61_8 = t_r33_c61_4 + p_34_60;
  assign t_r33_c61_9 = t_r33_c61_5 + t_r33_c61_6;
  assign t_r33_c61_10 = t_r33_c61_7 + t_r33_c61_8;
  assign t_r33_c61_11 = t_r33_c61_9 + t_r33_c61_10;
  assign t_r33_c61_12 = t_r33_c61_11 + p_34_62;
  assign out_33_61 = t_r33_c61_12 >> 4;

  assign t_r33_c62_0 = p_32_62 << 1;
  assign t_r33_c62_1 = p_33_61 << 1;
  assign t_r33_c62_2 = p_33_62 << 2;
  assign t_r33_c62_3 = p_33_63 << 1;
  assign t_r33_c62_4 = p_34_62 << 1;
  assign t_r33_c62_5 = t_r33_c62_0 + p_32_61;
  assign t_r33_c62_6 = t_r33_c62_1 + p_32_63;
  assign t_r33_c62_7 = t_r33_c62_2 + t_r33_c62_3;
  assign t_r33_c62_8 = t_r33_c62_4 + p_34_61;
  assign t_r33_c62_9 = t_r33_c62_5 + t_r33_c62_6;
  assign t_r33_c62_10 = t_r33_c62_7 + t_r33_c62_8;
  assign t_r33_c62_11 = t_r33_c62_9 + t_r33_c62_10;
  assign t_r33_c62_12 = t_r33_c62_11 + p_34_63;
  assign out_33_62 = t_r33_c62_12 >> 4;

  assign t_r33_c63_0 = p_32_63 << 1;
  assign t_r33_c63_1 = p_33_62 << 1;
  assign t_r33_c63_2 = p_33_63 << 2;
  assign t_r33_c63_3 = p_33_64 << 1;
  assign t_r33_c63_4 = p_34_63 << 1;
  assign t_r33_c63_5 = t_r33_c63_0 + p_32_62;
  assign t_r33_c63_6 = t_r33_c63_1 + p_32_64;
  assign t_r33_c63_7 = t_r33_c63_2 + t_r33_c63_3;
  assign t_r33_c63_8 = t_r33_c63_4 + p_34_62;
  assign t_r33_c63_9 = t_r33_c63_5 + t_r33_c63_6;
  assign t_r33_c63_10 = t_r33_c63_7 + t_r33_c63_8;
  assign t_r33_c63_11 = t_r33_c63_9 + t_r33_c63_10;
  assign t_r33_c63_12 = t_r33_c63_11 + p_34_64;
  assign out_33_63 = t_r33_c63_12 >> 4;

  assign t_r33_c64_0 = p_32_64 << 1;
  assign t_r33_c64_1 = p_33_63 << 1;
  assign t_r33_c64_2 = p_33_64 << 2;
  assign t_r33_c64_3 = p_33_65 << 1;
  assign t_r33_c64_4 = p_34_64 << 1;
  assign t_r33_c64_5 = t_r33_c64_0 + p_32_63;
  assign t_r33_c64_6 = t_r33_c64_1 + p_32_65;
  assign t_r33_c64_7 = t_r33_c64_2 + t_r33_c64_3;
  assign t_r33_c64_8 = t_r33_c64_4 + p_34_63;
  assign t_r33_c64_9 = t_r33_c64_5 + t_r33_c64_6;
  assign t_r33_c64_10 = t_r33_c64_7 + t_r33_c64_8;
  assign t_r33_c64_11 = t_r33_c64_9 + t_r33_c64_10;
  assign t_r33_c64_12 = t_r33_c64_11 + p_34_65;
  assign out_33_64 = t_r33_c64_12 >> 4;

  assign t_r34_c1_0 = p_33_1 << 1;
  assign t_r34_c1_1 = p_34_0 << 1;
  assign t_r34_c1_2 = p_34_1 << 2;
  assign t_r34_c1_3 = p_34_2 << 1;
  assign t_r34_c1_4 = p_35_1 << 1;
  assign t_r34_c1_5 = t_r34_c1_0 + p_33_0;
  assign t_r34_c1_6 = t_r34_c1_1 + p_33_2;
  assign t_r34_c1_7 = t_r34_c1_2 + t_r34_c1_3;
  assign t_r34_c1_8 = t_r34_c1_4 + p_35_0;
  assign t_r34_c1_9 = t_r34_c1_5 + t_r34_c1_6;
  assign t_r34_c1_10 = t_r34_c1_7 + t_r34_c1_8;
  assign t_r34_c1_11 = t_r34_c1_9 + t_r34_c1_10;
  assign t_r34_c1_12 = t_r34_c1_11 + p_35_2;
  assign out_34_1 = t_r34_c1_12 >> 4;

  assign t_r34_c2_0 = p_33_2 << 1;
  assign t_r34_c2_1 = p_34_1 << 1;
  assign t_r34_c2_2 = p_34_2 << 2;
  assign t_r34_c2_3 = p_34_3 << 1;
  assign t_r34_c2_4 = p_35_2 << 1;
  assign t_r34_c2_5 = t_r34_c2_0 + p_33_1;
  assign t_r34_c2_6 = t_r34_c2_1 + p_33_3;
  assign t_r34_c2_7 = t_r34_c2_2 + t_r34_c2_3;
  assign t_r34_c2_8 = t_r34_c2_4 + p_35_1;
  assign t_r34_c2_9 = t_r34_c2_5 + t_r34_c2_6;
  assign t_r34_c2_10 = t_r34_c2_7 + t_r34_c2_8;
  assign t_r34_c2_11 = t_r34_c2_9 + t_r34_c2_10;
  assign t_r34_c2_12 = t_r34_c2_11 + p_35_3;
  assign out_34_2 = t_r34_c2_12 >> 4;

  assign t_r34_c3_0 = p_33_3 << 1;
  assign t_r34_c3_1 = p_34_2 << 1;
  assign t_r34_c3_2 = p_34_3 << 2;
  assign t_r34_c3_3 = p_34_4 << 1;
  assign t_r34_c3_4 = p_35_3 << 1;
  assign t_r34_c3_5 = t_r34_c3_0 + p_33_2;
  assign t_r34_c3_6 = t_r34_c3_1 + p_33_4;
  assign t_r34_c3_7 = t_r34_c3_2 + t_r34_c3_3;
  assign t_r34_c3_8 = t_r34_c3_4 + p_35_2;
  assign t_r34_c3_9 = t_r34_c3_5 + t_r34_c3_6;
  assign t_r34_c3_10 = t_r34_c3_7 + t_r34_c3_8;
  assign t_r34_c3_11 = t_r34_c3_9 + t_r34_c3_10;
  assign t_r34_c3_12 = t_r34_c3_11 + p_35_4;
  assign out_34_3 = t_r34_c3_12 >> 4;

  assign t_r34_c4_0 = p_33_4 << 1;
  assign t_r34_c4_1 = p_34_3 << 1;
  assign t_r34_c4_2 = p_34_4 << 2;
  assign t_r34_c4_3 = p_34_5 << 1;
  assign t_r34_c4_4 = p_35_4 << 1;
  assign t_r34_c4_5 = t_r34_c4_0 + p_33_3;
  assign t_r34_c4_6 = t_r34_c4_1 + p_33_5;
  assign t_r34_c4_7 = t_r34_c4_2 + t_r34_c4_3;
  assign t_r34_c4_8 = t_r34_c4_4 + p_35_3;
  assign t_r34_c4_9 = t_r34_c4_5 + t_r34_c4_6;
  assign t_r34_c4_10 = t_r34_c4_7 + t_r34_c4_8;
  assign t_r34_c4_11 = t_r34_c4_9 + t_r34_c4_10;
  assign t_r34_c4_12 = t_r34_c4_11 + p_35_5;
  assign out_34_4 = t_r34_c4_12 >> 4;

  assign t_r34_c5_0 = p_33_5 << 1;
  assign t_r34_c5_1 = p_34_4 << 1;
  assign t_r34_c5_2 = p_34_5 << 2;
  assign t_r34_c5_3 = p_34_6 << 1;
  assign t_r34_c5_4 = p_35_5 << 1;
  assign t_r34_c5_5 = t_r34_c5_0 + p_33_4;
  assign t_r34_c5_6 = t_r34_c5_1 + p_33_6;
  assign t_r34_c5_7 = t_r34_c5_2 + t_r34_c5_3;
  assign t_r34_c5_8 = t_r34_c5_4 + p_35_4;
  assign t_r34_c5_9 = t_r34_c5_5 + t_r34_c5_6;
  assign t_r34_c5_10 = t_r34_c5_7 + t_r34_c5_8;
  assign t_r34_c5_11 = t_r34_c5_9 + t_r34_c5_10;
  assign t_r34_c5_12 = t_r34_c5_11 + p_35_6;
  assign out_34_5 = t_r34_c5_12 >> 4;

  assign t_r34_c6_0 = p_33_6 << 1;
  assign t_r34_c6_1 = p_34_5 << 1;
  assign t_r34_c6_2 = p_34_6 << 2;
  assign t_r34_c6_3 = p_34_7 << 1;
  assign t_r34_c6_4 = p_35_6 << 1;
  assign t_r34_c6_5 = t_r34_c6_0 + p_33_5;
  assign t_r34_c6_6 = t_r34_c6_1 + p_33_7;
  assign t_r34_c6_7 = t_r34_c6_2 + t_r34_c6_3;
  assign t_r34_c6_8 = t_r34_c6_4 + p_35_5;
  assign t_r34_c6_9 = t_r34_c6_5 + t_r34_c6_6;
  assign t_r34_c6_10 = t_r34_c6_7 + t_r34_c6_8;
  assign t_r34_c6_11 = t_r34_c6_9 + t_r34_c6_10;
  assign t_r34_c6_12 = t_r34_c6_11 + p_35_7;
  assign out_34_6 = t_r34_c6_12 >> 4;

  assign t_r34_c7_0 = p_33_7 << 1;
  assign t_r34_c7_1 = p_34_6 << 1;
  assign t_r34_c7_2 = p_34_7 << 2;
  assign t_r34_c7_3 = p_34_8 << 1;
  assign t_r34_c7_4 = p_35_7 << 1;
  assign t_r34_c7_5 = t_r34_c7_0 + p_33_6;
  assign t_r34_c7_6 = t_r34_c7_1 + p_33_8;
  assign t_r34_c7_7 = t_r34_c7_2 + t_r34_c7_3;
  assign t_r34_c7_8 = t_r34_c7_4 + p_35_6;
  assign t_r34_c7_9 = t_r34_c7_5 + t_r34_c7_6;
  assign t_r34_c7_10 = t_r34_c7_7 + t_r34_c7_8;
  assign t_r34_c7_11 = t_r34_c7_9 + t_r34_c7_10;
  assign t_r34_c7_12 = t_r34_c7_11 + p_35_8;
  assign out_34_7 = t_r34_c7_12 >> 4;

  assign t_r34_c8_0 = p_33_8 << 1;
  assign t_r34_c8_1 = p_34_7 << 1;
  assign t_r34_c8_2 = p_34_8 << 2;
  assign t_r34_c8_3 = p_34_9 << 1;
  assign t_r34_c8_4 = p_35_8 << 1;
  assign t_r34_c8_5 = t_r34_c8_0 + p_33_7;
  assign t_r34_c8_6 = t_r34_c8_1 + p_33_9;
  assign t_r34_c8_7 = t_r34_c8_2 + t_r34_c8_3;
  assign t_r34_c8_8 = t_r34_c8_4 + p_35_7;
  assign t_r34_c8_9 = t_r34_c8_5 + t_r34_c8_6;
  assign t_r34_c8_10 = t_r34_c8_7 + t_r34_c8_8;
  assign t_r34_c8_11 = t_r34_c8_9 + t_r34_c8_10;
  assign t_r34_c8_12 = t_r34_c8_11 + p_35_9;
  assign out_34_8 = t_r34_c8_12 >> 4;

  assign t_r34_c9_0 = p_33_9 << 1;
  assign t_r34_c9_1 = p_34_8 << 1;
  assign t_r34_c9_2 = p_34_9 << 2;
  assign t_r34_c9_3 = p_34_10 << 1;
  assign t_r34_c9_4 = p_35_9 << 1;
  assign t_r34_c9_5 = t_r34_c9_0 + p_33_8;
  assign t_r34_c9_6 = t_r34_c9_1 + p_33_10;
  assign t_r34_c9_7 = t_r34_c9_2 + t_r34_c9_3;
  assign t_r34_c9_8 = t_r34_c9_4 + p_35_8;
  assign t_r34_c9_9 = t_r34_c9_5 + t_r34_c9_6;
  assign t_r34_c9_10 = t_r34_c9_7 + t_r34_c9_8;
  assign t_r34_c9_11 = t_r34_c9_9 + t_r34_c9_10;
  assign t_r34_c9_12 = t_r34_c9_11 + p_35_10;
  assign out_34_9 = t_r34_c9_12 >> 4;

  assign t_r34_c10_0 = p_33_10 << 1;
  assign t_r34_c10_1 = p_34_9 << 1;
  assign t_r34_c10_2 = p_34_10 << 2;
  assign t_r34_c10_3 = p_34_11 << 1;
  assign t_r34_c10_4 = p_35_10 << 1;
  assign t_r34_c10_5 = t_r34_c10_0 + p_33_9;
  assign t_r34_c10_6 = t_r34_c10_1 + p_33_11;
  assign t_r34_c10_7 = t_r34_c10_2 + t_r34_c10_3;
  assign t_r34_c10_8 = t_r34_c10_4 + p_35_9;
  assign t_r34_c10_9 = t_r34_c10_5 + t_r34_c10_6;
  assign t_r34_c10_10 = t_r34_c10_7 + t_r34_c10_8;
  assign t_r34_c10_11 = t_r34_c10_9 + t_r34_c10_10;
  assign t_r34_c10_12 = t_r34_c10_11 + p_35_11;
  assign out_34_10 = t_r34_c10_12 >> 4;

  assign t_r34_c11_0 = p_33_11 << 1;
  assign t_r34_c11_1 = p_34_10 << 1;
  assign t_r34_c11_2 = p_34_11 << 2;
  assign t_r34_c11_3 = p_34_12 << 1;
  assign t_r34_c11_4 = p_35_11 << 1;
  assign t_r34_c11_5 = t_r34_c11_0 + p_33_10;
  assign t_r34_c11_6 = t_r34_c11_1 + p_33_12;
  assign t_r34_c11_7 = t_r34_c11_2 + t_r34_c11_3;
  assign t_r34_c11_8 = t_r34_c11_4 + p_35_10;
  assign t_r34_c11_9 = t_r34_c11_5 + t_r34_c11_6;
  assign t_r34_c11_10 = t_r34_c11_7 + t_r34_c11_8;
  assign t_r34_c11_11 = t_r34_c11_9 + t_r34_c11_10;
  assign t_r34_c11_12 = t_r34_c11_11 + p_35_12;
  assign out_34_11 = t_r34_c11_12 >> 4;

  assign t_r34_c12_0 = p_33_12 << 1;
  assign t_r34_c12_1 = p_34_11 << 1;
  assign t_r34_c12_2 = p_34_12 << 2;
  assign t_r34_c12_3 = p_34_13 << 1;
  assign t_r34_c12_4 = p_35_12 << 1;
  assign t_r34_c12_5 = t_r34_c12_0 + p_33_11;
  assign t_r34_c12_6 = t_r34_c12_1 + p_33_13;
  assign t_r34_c12_7 = t_r34_c12_2 + t_r34_c12_3;
  assign t_r34_c12_8 = t_r34_c12_4 + p_35_11;
  assign t_r34_c12_9 = t_r34_c12_5 + t_r34_c12_6;
  assign t_r34_c12_10 = t_r34_c12_7 + t_r34_c12_8;
  assign t_r34_c12_11 = t_r34_c12_9 + t_r34_c12_10;
  assign t_r34_c12_12 = t_r34_c12_11 + p_35_13;
  assign out_34_12 = t_r34_c12_12 >> 4;

  assign t_r34_c13_0 = p_33_13 << 1;
  assign t_r34_c13_1 = p_34_12 << 1;
  assign t_r34_c13_2 = p_34_13 << 2;
  assign t_r34_c13_3 = p_34_14 << 1;
  assign t_r34_c13_4 = p_35_13 << 1;
  assign t_r34_c13_5 = t_r34_c13_0 + p_33_12;
  assign t_r34_c13_6 = t_r34_c13_1 + p_33_14;
  assign t_r34_c13_7 = t_r34_c13_2 + t_r34_c13_3;
  assign t_r34_c13_8 = t_r34_c13_4 + p_35_12;
  assign t_r34_c13_9 = t_r34_c13_5 + t_r34_c13_6;
  assign t_r34_c13_10 = t_r34_c13_7 + t_r34_c13_8;
  assign t_r34_c13_11 = t_r34_c13_9 + t_r34_c13_10;
  assign t_r34_c13_12 = t_r34_c13_11 + p_35_14;
  assign out_34_13 = t_r34_c13_12 >> 4;

  assign t_r34_c14_0 = p_33_14 << 1;
  assign t_r34_c14_1 = p_34_13 << 1;
  assign t_r34_c14_2 = p_34_14 << 2;
  assign t_r34_c14_3 = p_34_15 << 1;
  assign t_r34_c14_4 = p_35_14 << 1;
  assign t_r34_c14_5 = t_r34_c14_0 + p_33_13;
  assign t_r34_c14_6 = t_r34_c14_1 + p_33_15;
  assign t_r34_c14_7 = t_r34_c14_2 + t_r34_c14_3;
  assign t_r34_c14_8 = t_r34_c14_4 + p_35_13;
  assign t_r34_c14_9 = t_r34_c14_5 + t_r34_c14_6;
  assign t_r34_c14_10 = t_r34_c14_7 + t_r34_c14_8;
  assign t_r34_c14_11 = t_r34_c14_9 + t_r34_c14_10;
  assign t_r34_c14_12 = t_r34_c14_11 + p_35_15;
  assign out_34_14 = t_r34_c14_12 >> 4;

  assign t_r34_c15_0 = p_33_15 << 1;
  assign t_r34_c15_1 = p_34_14 << 1;
  assign t_r34_c15_2 = p_34_15 << 2;
  assign t_r34_c15_3 = p_34_16 << 1;
  assign t_r34_c15_4 = p_35_15 << 1;
  assign t_r34_c15_5 = t_r34_c15_0 + p_33_14;
  assign t_r34_c15_6 = t_r34_c15_1 + p_33_16;
  assign t_r34_c15_7 = t_r34_c15_2 + t_r34_c15_3;
  assign t_r34_c15_8 = t_r34_c15_4 + p_35_14;
  assign t_r34_c15_9 = t_r34_c15_5 + t_r34_c15_6;
  assign t_r34_c15_10 = t_r34_c15_7 + t_r34_c15_8;
  assign t_r34_c15_11 = t_r34_c15_9 + t_r34_c15_10;
  assign t_r34_c15_12 = t_r34_c15_11 + p_35_16;
  assign out_34_15 = t_r34_c15_12 >> 4;

  assign t_r34_c16_0 = p_33_16 << 1;
  assign t_r34_c16_1 = p_34_15 << 1;
  assign t_r34_c16_2 = p_34_16 << 2;
  assign t_r34_c16_3 = p_34_17 << 1;
  assign t_r34_c16_4 = p_35_16 << 1;
  assign t_r34_c16_5 = t_r34_c16_0 + p_33_15;
  assign t_r34_c16_6 = t_r34_c16_1 + p_33_17;
  assign t_r34_c16_7 = t_r34_c16_2 + t_r34_c16_3;
  assign t_r34_c16_8 = t_r34_c16_4 + p_35_15;
  assign t_r34_c16_9 = t_r34_c16_5 + t_r34_c16_6;
  assign t_r34_c16_10 = t_r34_c16_7 + t_r34_c16_8;
  assign t_r34_c16_11 = t_r34_c16_9 + t_r34_c16_10;
  assign t_r34_c16_12 = t_r34_c16_11 + p_35_17;
  assign out_34_16 = t_r34_c16_12 >> 4;

  assign t_r34_c17_0 = p_33_17 << 1;
  assign t_r34_c17_1 = p_34_16 << 1;
  assign t_r34_c17_2 = p_34_17 << 2;
  assign t_r34_c17_3 = p_34_18 << 1;
  assign t_r34_c17_4 = p_35_17 << 1;
  assign t_r34_c17_5 = t_r34_c17_0 + p_33_16;
  assign t_r34_c17_6 = t_r34_c17_1 + p_33_18;
  assign t_r34_c17_7 = t_r34_c17_2 + t_r34_c17_3;
  assign t_r34_c17_8 = t_r34_c17_4 + p_35_16;
  assign t_r34_c17_9 = t_r34_c17_5 + t_r34_c17_6;
  assign t_r34_c17_10 = t_r34_c17_7 + t_r34_c17_8;
  assign t_r34_c17_11 = t_r34_c17_9 + t_r34_c17_10;
  assign t_r34_c17_12 = t_r34_c17_11 + p_35_18;
  assign out_34_17 = t_r34_c17_12 >> 4;

  assign t_r34_c18_0 = p_33_18 << 1;
  assign t_r34_c18_1 = p_34_17 << 1;
  assign t_r34_c18_2 = p_34_18 << 2;
  assign t_r34_c18_3 = p_34_19 << 1;
  assign t_r34_c18_4 = p_35_18 << 1;
  assign t_r34_c18_5 = t_r34_c18_0 + p_33_17;
  assign t_r34_c18_6 = t_r34_c18_1 + p_33_19;
  assign t_r34_c18_7 = t_r34_c18_2 + t_r34_c18_3;
  assign t_r34_c18_8 = t_r34_c18_4 + p_35_17;
  assign t_r34_c18_9 = t_r34_c18_5 + t_r34_c18_6;
  assign t_r34_c18_10 = t_r34_c18_7 + t_r34_c18_8;
  assign t_r34_c18_11 = t_r34_c18_9 + t_r34_c18_10;
  assign t_r34_c18_12 = t_r34_c18_11 + p_35_19;
  assign out_34_18 = t_r34_c18_12 >> 4;

  assign t_r34_c19_0 = p_33_19 << 1;
  assign t_r34_c19_1 = p_34_18 << 1;
  assign t_r34_c19_2 = p_34_19 << 2;
  assign t_r34_c19_3 = p_34_20 << 1;
  assign t_r34_c19_4 = p_35_19 << 1;
  assign t_r34_c19_5 = t_r34_c19_0 + p_33_18;
  assign t_r34_c19_6 = t_r34_c19_1 + p_33_20;
  assign t_r34_c19_7 = t_r34_c19_2 + t_r34_c19_3;
  assign t_r34_c19_8 = t_r34_c19_4 + p_35_18;
  assign t_r34_c19_9 = t_r34_c19_5 + t_r34_c19_6;
  assign t_r34_c19_10 = t_r34_c19_7 + t_r34_c19_8;
  assign t_r34_c19_11 = t_r34_c19_9 + t_r34_c19_10;
  assign t_r34_c19_12 = t_r34_c19_11 + p_35_20;
  assign out_34_19 = t_r34_c19_12 >> 4;

  assign t_r34_c20_0 = p_33_20 << 1;
  assign t_r34_c20_1 = p_34_19 << 1;
  assign t_r34_c20_2 = p_34_20 << 2;
  assign t_r34_c20_3 = p_34_21 << 1;
  assign t_r34_c20_4 = p_35_20 << 1;
  assign t_r34_c20_5 = t_r34_c20_0 + p_33_19;
  assign t_r34_c20_6 = t_r34_c20_1 + p_33_21;
  assign t_r34_c20_7 = t_r34_c20_2 + t_r34_c20_3;
  assign t_r34_c20_8 = t_r34_c20_4 + p_35_19;
  assign t_r34_c20_9 = t_r34_c20_5 + t_r34_c20_6;
  assign t_r34_c20_10 = t_r34_c20_7 + t_r34_c20_8;
  assign t_r34_c20_11 = t_r34_c20_9 + t_r34_c20_10;
  assign t_r34_c20_12 = t_r34_c20_11 + p_35_21;
  assign out_34_20 = t_r34_c20_12 >> 4;

  assign t_r34_c21_0 = p_33_21 << 1;
  assign t_r34_c21_1 = p_34_20 << 1;
  assign t_r34_c21_2 = p_34_21 << 2;
  assign t_r34_c21_3 = p_34_22 << 1;
  assign t_r34_c21_4 = p_35_21 << 1;
  assign t_r34_c21_5 = t_r34_c21_0 + p_33_20;
  assign t_r34_c21_6 = t_r34_c21_1 + p_33_22;
  assign t_r34_c21_7 = t_r34_c21_2 + t_r34_c21_3;
  assign t_r34_c21_8 = t_r34_c21_4 + p_35_20;
  assign t_r34_c21_9 = t_r34_c21_5 + t_r34_c21_6;
  assign t_r34_c21_10 = t_r34_c21_7 + t_r34_c21_8;
  assign t_r34_c21_11 = t_r34_c21_9 + t_r34_c21_10;
  assign t_r34_c21_12 = t_r34_c21_11 + p_35_22;
  assign out_34_21 = t_r34_c21_12 >> 4;

  assign t_r34_c22_0 = p_33_22 << 1;
  assign t_r34_c22_1 = p_34_21 << 1;
  assign t_r34_c22_2 = p_34_22 << 2;
  assign t_r34_c22_3 = p_34_23 << 1;
  assign t_r34_c22_4 = p_35_22 << 1;
  assign t_r34_c22_5 = t_r34_c22_0 + p_33_21;
  assign t_r34_c22_6 = t_r34_c22_1 + p_33_23;
  assign t_r34_c22_7 = t_r34_c22_2 + t_r34_c22_3;
  assign t_r34_c22_8 = t_r34_c22_4 + p_35_21;
  assign t_r34_c22_9 = t_r34_c22_5 + t_r34_c22_6;
  assign t_r34_c22_10 = t_r34_c22_7 + t_r34_c22_8;
  assign t_r34_c22_11 = t_r34_c22_9 + t_r34_c22_10;
  assign t_r34_c22_12 = t_r34_c22_11 + p_35_23;
  assign out_34_22 = t_r34_c22_12 >> 4;

  assign t_r34_c23_0 = p_33_23 << 1;
  assign t_r34_c23_1 = p_34_22 << 1;
  assign t_r34_c23_2 = p_34_23 << 2;
  assign t_r34_c23_3 = p_34_24 << 1;
  assign t_r34_c23_4 = p_35_23 << 1;
  assign t_r34_c23_5 = t_r34_c23_0 + p_33_22;
  assign t_r34_c23_6 = t_r34_c23_1 + p_33_24;
  assign t_r34_c23_7 = t_r34_c23_2 + t_r34_c23_3;
  assign t_r34_c23_8 = t_r34_c23_4 + p_35_22;
  assign t_r34_c23_9 = t_r34_c23_5 + t_r34_c23_6;
  assign t_r34_c23_10 = t_r34_c23_7 + t_r34_c23_8;
  assign t_r34_c23_11 = t_r34_c23_9 + t_r34_c23_10;
  assign t_r34_c23_12 = t_r34_c23_11 + p_35_24;
  assign out_34_23 = t_r34_c23_12 >> 4;

  assign t_r34_c24_0 = p_33_24 << 1;
  assign t_r34_c24_1 = p_34_23 << 1;
  assign t_r34_c24_2 = p_34_24 << 2;
  assign t_r34_c24_3 = p_34_25 << 1;
  assign t_r34_c24_4 = p_35_24 << 1;
  assign t_r34_c24_5 = t_r34_c24_0 + p_33_23;
  assign t_r34_c24_6 = t_r34_c24_1 + p_33_25;
  assign t_r34_c24_7 = t_r34_c24_2 + t_r34_c24_3;
  assign t_r34_c24_8 = t_r34_c24_4 + p_35_23;
  assign t_r34_c24_9 = t_r34_c24_5 + t_r34_c24_6;
  assign t_r34_c24_10 = t_r34_c24_7 + t_r34_c24_8;
  assign t_r34_c24_11 = t_r34_c24_9 + t_r34_c24_10;
  assign t_r34_c24_12 = t_r34_c24_11 + p_35_25;
  assign out_34_24 = t_r34_c24_12 >> 4;

  assign t_r34_c25_0 = p_33_25 << 1;
  assign t_r34_c25_1 = p_34_24 << 1;
  assign t_r34_c25_2 = p_34_25 << 2;
  assign t_r34_c25_3 = p_34_26 << 1;
  assign t_r34_c25_4 = p_35_25 << 1;
  assign t_r34_c25_5 = t_r34_c25_0 + p_33_24;
  assign t_r34_c25_6 = t_r34_c25_1 + p_33_26;
  assign t_r34_c25_7 = t_r34_c25_2 + t_r34_c25_3;
  assign t_r34_c25_8 = t_r34_c25_4 + p_35_24;
  assign t_r34_c25_9 = t_r34_c25_5 + t_r34_c25_6;
  assign t_r34_c25_10 = t_r34_c25_7 + t_r34_c25_8;
  assign t_r34_c25_11 = t_r34_c25_9 + t_r34_c25_10;
  assign t_r34_c25_12 = t_r34_c25_11 + p_35_26;
  assign out_34_25 = t_r34_c25_12 >> 4;

  assign t_r34_c26_0 = p_33_26 << 1;
  assign t_r34_c26_1 = p_34_25 << 1;
  assign t_r34_c26_2 = p_34_26 << 2;
  assign t_r34_c26_3 = p_34_27 << 1;
  assign t_r34_c26_4 = p_35_26 << 1;
  assign t_r34_c26_5 = t_r34_c26_0 + p_33_25;
  assign t_r34_c26_6 = t_r34_c26_1 + p_33_27;
  assign t_r34_c26_7 = t_r34_c26_2 + t_r34_c26_3;
  assign t_r34_c26_8 = t_r34_c26_4 + p_35_25;
  assign t_r34_c26_9 = t_r34_c26_5 + t_r34_c26_6;
  assign t_r34_c26_10 = t_r34_c26_7 + t_r34_c26_8;
  assign t_r34_c26_11 = t_r34_c26_9 + t_r34_c26_10;
  assign t_r34_c26_12 = t_r34_c26_11 + p_35_27;
  assign out_34_26 = t_r34_c26_12 >> 4;

  assign t_r34_c27_0 = p_33_27 << 1;
  assign t_r34_c27_1 = p_34_26 << 1;
  assign t_r34_c27_2 = p_34_27 << 2;
  assign t_r34_c27_3 = p_34_28 << 1;
  assign t_r34_c27_4 = p_35_27 << 1;
  assign t_r34_c27_5 = t_r34_c27_0 + p_33_26;
  assign t_r34_c27_6 = t_r34_c27_1 + p_33_28;
  assign t_r34_c27_7 = t_r34_c27_2 + t_r34_c27_3;
  assign t_r34_c27_8 = t_r34_c27_4 + p_35_26;
  assign t_r34_c27_9 = t_r34_c27_5 + t_r34_c27_6;
  assign t_r34_c27_10 = t_r34_c27_7 + t_r34_c27_8;
  assign t_r34_c27_11 = t_r34_c27_9 + t_r34_c27_10;
  assign t_r34_c27_12 = t_r34_c27_11 + p_35_28;
  assign out_34_27 = t_r34_c27_12 >> 4;

  assign t_r34_c28_0 = p_33_28 << 1;
  assign t_r34_c28_1 = p_34_27 << 1;
  assign t_r34_c28_2 = p_34_28 << 2;
  assign t_r34_c28_3 = p_34_29 << 1;
  assign t_r34_c28_4 = p_35_28 << 1;
  assign t_r34_c28_5 = t_r34_c28_0 + p_33_27;
  assign t_r34_c28_6 = t_r34_c28_1 + p_33_29;
  assign t_r34_c28_7 = t_r34_c28_2 + t_r34_c28_3;
  assign t_r34_c28_8 = t_r34_c28_4 + p_35_27;
  assign t_r34_c28_9 = t_r34_c28_5 + t_r34_c28_6;
  assign t_r34_c28_10 = t_r34_c28_7 + t_r34_c28_8;
  assign t_r34_c28_11 = t_r34_c28_9 + t_r34_c28_10;
  assign t_r34_c28_12 = t_r34_c28_11 + p_35_29;
  assign out_34_28 = t_r34_c28_12 >> 4;

  assign t_r34_c29_0 = p_33_29 << 1;
  assign t_r34_c29_1 = p_34_28 << 1;
  assign t_r34_c29_2 = p_34_29 << 2;
  assign t_r34_c29_3 = p_34_30 << 1;
  assign t_r34_c29_4 = p_35_29 << 1;
  assign t_r34_c29_5 = t_r34_c29_0 + p_33_28;
  assign t_r34_c29_6 = t_r34_c29_1 + p_33_30;
  assign t_r34_c29_7 = t_r34_c29_2 + t_r34_c29_3;
  assign t_r34_c29_8 = t_r34_c29_4 + p_35_28;
  assign t_r34_c29_9 = t_r34_c29_5 + t_r34_c29_6;
  assign t_r34_c29_10 = t_r34_c29_7 + t_r34_c29_8;
  assign t_r34_c29_11 = t_r34_c29_9 + t_r34_c29_10;
  assign t_r34_c29_12 = t_r34_c29_11 + p_35_30;
  assign out_34_29 = t_r34_c29_12 >> 4;

  assign t_r34_c30_0 = p_33_30 << 1;
  assign t_r34_c30_1 = p_34_29 << 1;
  assign t_r34_c30_2 = p_34_30 << 2;
  assign t_r34_c30_3 = p_34_31 << 1;
  assign t_r34_c30_4 = p_35_30 << 1;
  assign t_r34_c30_5 = t_r34_c30_0 + p_33_29;
  assign t_r34_c30_6 = t_r34_c30_1 + p_33_31;
  assign t_r34_c30_7 = t_r34_c30_2 + t_r34_c30_3;
  assign t_r34_c30_8 = t_r34_c30_4 + p_35_29;
  assign t_r34_c30_9 = t_r34_c30_5 + t_r34_c30_6;
  assign t_r34_c30_10 = t_r34_c30_7 + t_r34_c30_8;
  assign t_r34_c30_11 = t_r34_c30_9 + t_r34_c30_10;
  assign t_r34_c30_12 = t_r34_c30_11 + p_35_31;
  assign out_34_30 = t_r34_c30_12 >> 4;

  assign t_r34_c31_0 = p_33_31 << 1;
  assign t_r34_c31_1 = p_34_30 << 1;
  assign t_r34_c31_2 = p_34_31 << 2;
  assign t_r34_c31_3 = p_34_32 << 1;
  assign t_r34_c31_4 = p_35_31 << 1;
  assign t_r34_c31_5 = t_r34_c31_0 + p_33_30;
  assign t_r34_c31_6 = t_r34_c31_1 + p_33_32;
  assign t_r34_c31_7 = t_r34_c31_2 + t_r34_c31_3;
  assign t_r34_c31_8 = t_r34_c31_4 + p_35_30;
  assign t_r34_c31_9 = t_r34_c31_5 + t_r34_c31_6;
  assign t_r34_c31_10 = t_r34_c31_7 + t_r34_c31_8;
  assign t_r34_c31_11 = t_r34_c31_9 + t_r34_c31_10;
  assign t_r34_c31_12 = t_r34_c31_11 + p_35_32;
  assign out_34_31 = t_r34_c31_12 >> 4;

  assign t_r34_c32_0 = p_33_32 << 1;
  assign t_r34_c32_1 = p_34_31 << 1;
  assign t_r34_c32_2 = p_34_32 << 2;
  assign t_r34_c32_3 = p_34_33 << 1;
  assign t_r34_c32_4 = p_35_32 << 1;
  assign t_r34_c32_5 = t_r34_c32_0 + p_33_31;
  assign t_r34_c32_6 = t_r34_c32_1 + p_33_33;
  assign t_r34_c32_7 = t_r34_c32_2 + t_r34_c32_3;
  assign t_r34_c32_8 = t_r34_c32_4 + p_35_31;
  assign t_r34_c32_9 = t_r34_c32_5 + t_r34_c32_6;
  assign t_r34_c32_10 = t_r34_c32_7 + t_r34_c32_8;
  assign t_r34_c32_11 = t_r34_c32_9 + t_r34_c32_10;
  assign t_r34_c32_12 = t_r34_c32_11 + p_35_33;
  assign out_34_32 = t_r34_c32_12 >> 4;

  assign t_r34_c33_0 = p_33_33 << 1;
  assign t_r34_c33_1 = p_34_32 << 1;
  assign t_r34_c33_2 = p_34_33 << 2;
  assign t_r34_c33_3 = p_34_34 << 1;
  assign t_r34_c33_4 = p_35_33 << 1;
  assign t_r34_c33_5 = t_r34_c33_0 + p_33_32;
  assign t_r34_c33_6 = t_r34_c33_1 + p_33_34;
  assign t_r34_c33_7 = t_r34_c33_2 + t_r34_c33_3;
  assign t_r34_c33_8 = t_r34_c33_4 + p_35_32;
  assign t_r34_c33_9 = t_r34_c33_5 + t_r34_c33_6;
  assign t_r34_c33_10 = t_r34_c33_7 + t_r34_c33_8;
  assign t_r34_c33_11 = t_r34_c33_9 + t_r34_c33_10;
  assign t_r34_c33_12 = t_r34_c33_11 + p_35_34;
  assign out_34_33 = t_r34_c33_12 >> 4;

  assign t_r34_c34_0 = p_33_34 << 1;
  assign t_r34_c34_1 = p_34_33 << 1;
  assign t_r34_c34_2 = p_34_34 << 2;
  assign t_r34_c34_3 = p_34_35 << 1;
  assign t_r34_c34_4 = p_35_34 << 1;
  assign t_r34_c34_5 = t_r34_c34_0 + p_33_33;
  assign t_r34_c34_6 = t_r34_c34_1 + p_33_35;
  assign t_r34_c34_7 = t_r34_c34_2 + t_r34_c34_3;
  assign t_r34_c34_8 = t_r34_c34_4 + p_35_33;
  assign t_r34_c34_9 = t_r34_c34_5 + t_r34_c34_6;
  assign t_r34_c34_10 = t_r34_c34_7 + t_r34_c34_8;
  assign t_r34_c34_11 = t_r34_c34_9 + t_r34_c34_10;
  assign t_r34_c34_12 = t_r34_c34_11 + p_35_35;
  assign out_34_34 = t_r34_c34_12 >> 4;

  assign t_r34_c35_0 = p_33_35 << 1;
  assign t_r34_c35_1 = p_34_34 << 1;
  assign t_r34_c35_2 = p_34_35 << 2;
  assign t_r34_c35_3 = p_34_36 << 1;
  assign t_r34_c35_4 = p_35_35 << 1;
  assign t_r34_c35_5 = t_r34_c35_0 + p_33_34;
  assign t_r34_c35_6 = t_r34_c35_1 + p_33_36;
  assign t_r34_c35_7 = t_r34_c35_2 + t_r34_c35_3;
  assign t_r34_c35_8 = t_r34_c35_4 + p_35_34;
  assign t_r34_c35_9 = t_r34_c35_5 + t_r34_c35_6;
  assign t_r34_c35_10 = t_r34_c35_7 + t_r34_c35_8;
  assign t_r34_c35_11 = t_r34_c35_9 + t_r34_c35_10;
  assign t_r34_c35_12 = t_r34_c35_11 + p_35_36;
  assign out_34_35 = t_r34_c35_12 >> 4;

  assign t_r34_c36_0 = p_33_36 << 1;
  assign t_r34_c36_1 = p_34_35 << 1;
  assign t_r34_c36_2 = p_34_36 << 2;
  assign t_r34_c36_3 = p_34_37 << 1;
  assign t_r34_c36_4 = p_35_36 << 1;
  assign t_r34_c36_5 = t_r34_c36_0 + p_33_35;
  assign t_r34_c36_6 = t_r34_c36_1 + p_33_37;
  assign t_r34_c36_7 = t_r34_c36_2 + t_r34_c36_3;
  assign t_r34_c36_8 = t_r34_c36_4 + p_35_35;
  assign t_r34_c36_9 = t_r34_c36_5 + t_r34_c36_6;
  assign t_r34_c36_10 = t_r34_c36_7 + t_r34_c36_8;
  assign t_r34_c36_11 = t_r34_c36_9 + t_r34_c36_10;
  assign t_r34_c36_12 = t_r34_c36_11 + p_35_37;
  assign out_34_36 = t_r34_c36_12 >> 4;

  assign t_r34_c37_0 = p_33_37 << 1;
  assign t_r34_c37_1 = p_34_36 << 1;
  assign t_r34_c37_2 = p_34_37 << 2;
  assign t_r34_c37_3 = p_34_38 << 1;
  assign t_r34_c37_4 = p_35_37 << 1;
  assign t_r34_c37_5 = t_r34_c37_0 + p_33_36;
  assign t_r34_c37_6 = t_r34_c37_1 + p_33_38;
  assign t_r34_c37_7 = t_r34_c37_2 + t_r34_c37_3;
  assign t_r34_c37_8 = t_r34_c37_4 + p_35_36;
  assign t_r34_c37_9 = t_r34_c37_5 + t_r34_c37_6;
  assign t_r34_c37_10 = t_r34_c37_7 + t_r34_c37_8;
  assign t_r34_c37_11 = t_r34_c37_9 + t_r34_c37_10;
  assign t_r34_c37_12 = t_r34_c37_11 + p_35_38;
  assign out_34_37 = t_r34_c37_12 >> 4;

  assign t_r34_c38_0 = p_33_38 << 1;
  assign t_r34_c38_1 = p_34_37 << 1;
  assign t_r34_c38_2 = p_34_38 << 2;
  assign t_r34_c38_3 = p_34_39 << 1;
  assign t_r34_c38_4 = p_35_38 << 1;
  assign t_r34_c38_5 = t_r34_c38_0 + p_33_37;
  assign t_r34_c38_6 = t_r34_c38_1 + p_33_39;
  assign t_r34_c38_7 = t_r34_c38_2 + t_r34_c38_3;
  assign t_r34_c38_8 = t_r34_c38_4 + p_35_37;
  assign t_r34_c38_9 = t_r34_c38_5 + t_r34_c38_6;
  assign t_r34_c38_10 = t_r34_c38_7 + t_r34_c38_8;
  assign t_r34_c38_11 = t_r34_c38_9 + t_r34_c38_10;
  assign t_r34_c38_12 = t_r34_c38_11 + p_35_39;
  assign out_34_38 = t_r34_c38_12 >> 4;

  assign t_r34_c39_0 = p_33_39 << 1;
  assign t_r34_c39_1 = p_34_38 << 1;
  assign t_r34_c39_2 = p_34_39 << 2;
  assign t_r34_c39_3 = p_34_40 << 1;
  assign t_r34_c39_4 = p_35_39 << 1;
  assign t_r34_c39_5 = t_r34_c39_0 + p_33_38;
  assign t_r34_c39_6 = t_r34_c39_1 + p_33_40;
  assign t_r34_c39_7 = t_r34_c39_2 + t_r34_c39_3;
  assign t_r34_c39_8 = t_r34_c39_4 + p_35_38;
  assign t_r34_c39_9 = t_r34_c39_5 + t_r34_c39_6;
  assign t_r34_c39_10 = t_r34_c39_7 + t_r34_c39_8;
  assign t_r34_c39_11 = t_r34_c39_9 + t_r34_c39_10;
  assign t_r34_c39_12 = t_r34_c39_11 + p_35_40;
  assign out_34_39 = t_r34_c39_12 >> 4;

  assign t_r34_c40_0 = p_33_40 << 1;
  assign t_r34_c40_1 = p_34_39 << 1;
  assign t_r34_c40_2 = p_34_40 << 2;
  assign t_r34_c40_3 = p_34_41 << 1;
  assign t_r34_c40_4 = p_35_40 << 1;
  assign t_r34_c40_5 = t_r34_c40_0 + p_33_39;
  assign t_r34_c40_6 = t_r34_c40_1 + p_33_41;
  assign t_r34_c40_7 = t_r34_c40_2 + t_r34_c40_3;
  assign t_r34_c40_8 = t_r34_c40_4 + p_35_39;
  assign t_r34_c40_9 = t_r34_c40_5 + t_r34_c40_6;
  assign t_r34_c40_10 = t_r34_c40_7 + t_r34_c40_8;
  assign t_r34_c40_11 = t_r34_c40_9 + t_r34_c40_10;
  assign t_r34_c40_12 = t_r34_c40_11 + p_35_41;
  assign out_34_40 = t_r34_c40_12 >> 4;

  assign t_r34_c41_0 = p_33_41 << 1;
  assign t_r34_c41_1 = p_34_40 << 1;
  assign t_r34_c41_2 = p_34_41 << 2;
  assign t_r34_c41_3 = p_34_42 << 1;
  assign t_r34_c41_4 = p_35_41 << 1;
  assign t_r34_c41_5 = t_r34_c41_0 + p_33_40;
  assign t_r34_c41_6 = t_r34_c41_1 + p_33_42;
  assign t_r34_c41_7 = t_r34_c41_2 + t_r34_c41_3;
  assign t_r34_c41_8 = t_r34_c41_4 + p_35_40;
  assign t_r34_c41_9 = t_r34_c41_5 + t_r34_c41_6;
  assign t_r34_c41_10 = t_r34_c41_7 + t_r34_c41_8;
  assign t_r34_c41_11 = t_r34_c41_9 + t_r34_c41_10;
  assign t_r34_c41_12 = t_r34_c41_11 + p_35_42;
  assign out_34_41 = t_r34_c41_12 >> 4;

  assign t_r34_c42_0 = p_33_42 << 1;
  assign t_r34_c42_1 = p_34_41 << 1;
  assign t_r34_c42_2 = p_34_42 << 2;
  assign t_r34_c42_3 = p_34_43 << 1;
  assign t_r34_c42_4 = p_35_42 << 1;
  assign t_r34_c42_5 = t_r34_c42_0 + p_33_41;
  assign t_r34_c42_6 = t_r34_c42_1 + p_33_43;
  assign t_r34_c42_7 = t_r34_c42_2 + t_r34_c42_3;
  assign t_r34_c42_8 = t_r34_c42_4 + p_35_41;
  assign t_r34_c42_9 = t_r34_c42_5 + t_r34_c42_6;
  assign t_r34_c42_10 = t_r34_c42_7 + t_r34_c42_8;
  assign t_r34_c42_11 = t_r34_c42_9 + t_r34_c42_10;
  assign t_r34_c42_12 = t_r34_c42_11 + p_35_43;
  assign out_34_42 = t_r34_c42_12 >> 4;

  assign t_r34_c43_0 = p_33_43 << 1;
  assign t_r34_c43_1 = p_34_42 << 1;
  assign t_r34_c43_2 = p_34_43 << 2;
  assign t_r34_c43_3 = p_34_44 << 1;
  assign t_r34_c43_4 = p_35_43 << 1;
  assign t_r34_c43_5 = t_r34_c43_0 + p_33_42;
  assign t_r34_c43_6 = t_r34_c43_1 + p_33_44;
  assign t_r34_c43_7 = t_r34_c43_2 + t_r34_c43_3;
  assign t_r34_c43_8 = t_r34_c43_4 + p_35_42;
  assign t_r34_c43_9 = t_r34_c43_5 + t_r34_c43_6;
  assign t_r34_c43_10 = t_r34_c43_7 + t_r34_c43_8;
  assign t_r34_c43_11 = t_r34_c43_9 + t_r34_c43_10;
  assign t_r34_c43_12 = t_r34_c43_11 + p_35_44;
  assign out_34_43 = t_r34_c43_12 >> 4;

  assign t_r34_c44_0 = p_33_44 << 1;
  assign t_r34_c44_1 = p_34_43 << 1;
  assign t_r34_c44_2 = p_34_44 << 2;
  assign t_r34_c44_3 = p_34_45 << 1;
  assign t_r34_c44_4 = p_35_44 << 1;
  assign t_r34_c44_5 = t_r34_c44_0 + p_33_43;
  assign t_r34_c44_6 = t_r34_c44_1 + p_33_45;
  assign t_r34_c44_7 = t_r34_c44_2 + t_r34_c44_3;
  assign t_r34_c44_8 = t_r34_c44_4 + p_35_43;
  assign t_r34_c44_9 = t_r34_c44_5 + t_r34_c44_6;
  assign t_r34_c44_10 = t_r34_c44_7 + t_r34_c44_8;
  assign t_r34_c44_11 = t_r34_c44_9 + t_r34_c44_10;
  assign t_r34_c44_12 = t_r34_c44_11 + p_35_45;
  assign out_34_44 = t_r34_c44_12 >> 4;

  assign t_r34_c45_0 = p_33_45 << 1;
  assign t_r34_c45_1 = p_34_44 << 1;
  assign t_r34_c45_2 = p_34_45 << 2;
  assign t_r34_c45_3 = p_34_46 << 1;
  assign t_r34_c45_4 = p_35_45 << 1;
  assign t_r34_c45_5 = t_r34_c45_0 + p_33_44;
  assign t_r34_c45_6 = t_r34_c45_1 + p_33_46;
  assign t_r34_c45_7 = t_r34_c45_2 + t_r34_c45_3;
  assign t_r34_c45_8 = t_r34_c45_4 + p_35_44;
  assign t_r34_c45_9 = t_r34_c45_5 + t_r34_c45_6;
  assign t_r34_c45_10 = t_r34_c45_7 + t_r34_c45_8;
  assign t_r34_c45_11 = t_r34_c45_9 + t_r34_c45_10;
  assign t_r34_c45_12 = t_r34_c45_11 + p_35_46;
  assign out_34_45 = t_r34_c45_12 >> 4;

  assign t_r34_c46_0 = p_33_46 << 1;
  assign t_r34_c46_1 = p_34_45 << 1;
  assign t_r34_c46_2 = p_34_46 << 2;
  assign t_r34_c46_3 = p_34_47 << 1;
  assign t_r34_c46_4 = p_35_46 << 1;
  assign t_r34_c46_5 = t_r34_c46_0 + p_33_45;
  assign t_r34_c46_6 = t_r34_c46_1 + p_33_47;
  assign t_r34_c46_7 = t_r34_c46_2 + t_r34_c46_3;
  assign t_r34_c46_8 = t_r34_c46_4 + p_35_45;
  assign t_r34_c46_9 = t_r34_c46_5 + t_r34_c46_6;
  assign t_r34_c46_10 = t_r34_c46_7 + t_r34_c46_8;
  assign t_r34_c46_11 = t_r34_c46_9 + t_r34_c46_10;
  assign t_r34_c46_12 = t_r34_c46_11 + p_35_47;
  assign out_34_46 = t_r34_c46_12 >> 4;

  assign t_r34_c47_0 = p_33_47 << 1;
  assign t_r34_c47_1 = p_34_46 << 1;
  assign t_r34_c47_2 = p_34_47 << 2;
  assign t_r34_c47_3 = p_34_48 << 1;
  assign t_r34_c47_4 = p_35_47 << 1;
  assign t_r34_c47_5 = t_r34_c47_0 + p_33_46;
  assign t_r34_c47_6 = t_r34_c47_1 + p_33_48;
  assign t_r34_c47_7 = t_r34_c47_2 + t_r34_c47_3;
  assign t_r34_c47_8 = t_r34_c47_4 + p_35_46;
  assign t_r34_c47_9 = t_r34_c47_5 + t_r34_c47_6;
  assign t_r34_c47_10 = t_r34_c47_7 + t_r34_c47_8;
  assign t_r34_c47_11 = t_r34_c47_9 + t_r34_c47_10;
  assign t_r34_c47_12 = t_r34_c47_11 + p_35_48;
  assign out_34_47 = t_r34_c47_12 >> 4;

  assign t_r34_c48_0 = p_33_48 << 1;
  assign t_r34_c48_1 = p_34_47 << 1;
  assign t_r34_c48_2 = p_34_48 << 2;
  assign t_r34_c48_3 = p_34_49 << 1;
  assign t_r34_c48_4 = p_35_48 << 1;
  assign t_r34_c48_5 = t_r34_c48_0 + p_33_47;
  assign t_r34_c48_6 = t_r34_c48_1 + p_33_49;
  assign t_r34_c48_7 = t_r34_c48_2 + t_r34_c48_3;
  assign t_r34_c48_8 = t_r34_c48_4 + p_35_47;
  assign t_r34_c48_9 = t_r34_c48_5 + t_r34_c48_6;
  assign t_r34_c48_10 = t_r34_c48_7 + t_r34_c48_8;
  assign t_r34_c48_11 = t_r34_c48_9 + t_r34_c48_10;
  assign t_r34_c48_12 = t_r34_c48_11 + p_35_49;
  assign out_34_48 = t_r34_c48_12 >> 4;

  assign t_r34_c49_0 = p_33_49 << 1;
  assign t_r34_c49_1 = p_34_48 << 1;
  assign t_r34_c49_2 = p_34_49 << 2;
  assign t_r34_c49_3 = p_34_50 << 1;
  assign t_r34_c49_4 = p_35_49 << 1;
  assign t_r34_c49_5 = t_r34_c49_0 + p_33_48;
  assign t_r34_c49_6 = t_r34_c49_1 + p_33_50;
  assign t_r34_c49_7 = t_r34_c49_2 + t_r34_c49_3;
  assign t_r34_c49_8 = t_r34_c49_4 + p_35_48;
  assign t_r34_c49_9 = t_r34_c49_5 + t_r34_c49_6;
  assign t_r34_c49_10 = t_r34_c49_7 + t_r34_c49_8;
  assign t_r34_c49_11 = t_r34_c49_9 + t_r34_c49_10;
  assign t_r34_c49_12 = t_r34_c49_11 + p_35_50;
  assign out_34_49 = t_r34_c49_12 >> 4;

  assign t_r34_c50_0 = p_33_50 << 1;
  assign t_r34_c50_1 = p_34_49 << 1;
  assign t_r34_c50_2 = p_34_50 << 2;
  assign t_r34_c50_3 = p_34_51 << 1;
  assign t_r34_c50_4 = p_35_50 << 1;
  assign t_r34_c50_5 = t_r34_c50_0 + p_33_49;
  assign t_r34_c50_6 = t_r34_c50_1 + p_33_51;
  assign t_r34_c50_7 = t_r34_c50_2 + t_r34_c50_3;
  assign t_r34_c50_8 = t_r34_c50_4 + p_35_49;
  assign t_r34_c50_9 = t_r34_c50_5 + t_r34_c50_6;
  assign t_r34_c50_10 = t_r34_c50_7 + t_r34_c50_8;
  assign t_r34_c50_11 = t_r34_c50_9 + t_r34_c50_10;
  assign t_r34_c50_12 = t_r34_c50_11 + p_35_51;
  assign out_34_50 = t_r34_c50_12 >> 4;

  assign t_r34_c51_0 = p_33_51 << 1;
  assign t_r34_c51_1 = p_34_50 << 1;
  assign t_r34_c51_2 = p_34_51 << 2;
  assign t_r34_c51_3 = p_34_52 << 1;
  assign t_r34_c51_4 = p_35_51 << 1;
  assign t_r34_c51_5 = t_r34_c51_0 + p_33_50;
  assign t_r34_c51_6 = t_r34_c51_1 + p_33_52;
  assign t_r34_c51_7 = t_r34_c51_2 + t_r34_c51_3;
  assign t_r34_c51_8 = t_r34_c51_4 + p_35_50;
  assign t_r34_c51_9 = t_r34_c51_5 + t_r34_c51_6;
  assign t_r34_c51_10 = t_r34_c51_7 + t_r34_c51_8;
  assign t_r34_c51_11 = t_r34_c51_9 + t_r34_c51_10;
  assign t_r34_c51_12 = t_r34_c51_11 + p_35_52;
  assign out_34_51 = t_r34_c51_12 >> 4;

  assign t_r34_c52_0 = p_33_52 << 1;
  assign t_r34_c52_1 = p_34_51 << 1;
  assign t_r34_c52_2 = p_34_52 << 2;
  assign t_r34_c52_3 = p_34_53 << 1;
  assign t_r34_c52_4 = p_35_52 << 1;
  assign t_r34_c52_5 = t_r34_c52_0 + p_33_51;
  assign t_r34_c52_6 = t_r34_c52_1 + p_33_53;
  assign t_r34_c52_7 = t_r34_c52_2 + t_r34_c52_3;
  assign t_r34_c52_8 = t_r34_c52_4 + p_35_51;
  assign t_r34_c52_9 = t_r34_c52_5 + t_r34_c52_6;
  assign t_r34_c52_10 = t_r34_c52_7 + t_r34_c52_8;
  assign t_r34_c52_11 = t_r34_c52_9 + t_r34_c52_10;
  assign t_r34_c52_12 = t_r34_c52_11 + p_35_53;
  assign out_34_52 = t_r34_c52_12 >> 4;

  assign t_r34_c53_0 = p_33_53 << 1;
  assign t_r34_c53_1 = p_34_52 << 1;
  assign t_r34_c53_2 = p_34_53 << 2;
  assign t_r34_c53_3 = p_34_54 << 1;
  assign t_r34_c53_4 = p_35_53 << 1;
  assign t_r34_c53_5 = t_r34_c53_0 + p_33_52;
  assign t_r34_c53_6 = t_r34_c53_1 + p_33_54;
  assign t_r34_c53_7 = t_r34_c53_2 + t_r34_c53_3;
  assign t_r34_c53_8 = t_r34_c53_4 + p_35_52;
  assign t_r34_c53_9 = t_r34_c53_5 + t_r34_c53_6;
  assign t_r34_c53_10 = t_r34_c53_7 + t_r34_c53_8;
  assign t_r34_c53_11 = t_r34_c53_9 + t_r34_c53_10;
  assign t_r34_c53_12 = t_r34_c53_11 + p_35_54;
  assign out_34_53 = t_r34_c53_12 >> 4;

  assign t_r34_c54_0 = p_33_54 << 1;
  assign t_r34_c54_1 = p_34_53 << 1;
  assign t_r34_c54_2 = p_34_54 << 2;
  assign t_r34_c54_3 = p_34_55 << 1;
  assign t_r34_c54_4 = p_35_54 << 1;
  assign t_r34_c54_5 = t_r34_c54_0 + p_33_53;
  assign t_r34_c54_6 = t_r34_c54_1 + p_33_55;
  assign t_r34_c54_7 = t_r34_c54_2 + t_r34_c54_3;
  assign t_r34_c54_8 = t_r34_c54_4 + p_35_53;
  assign t_r34_c54_9 = t_r34_c54_5 + t_r34_c54_6;
  assign t_r34_c54_10 = t_r34_c54_7 + t_r34_c54_8;
  assign t_r34_c54_11 = t_r34_c54_9 + t_r34_c54_10;
  assign t_r34_c54_12 = t_r34_c54_11 + p_35_55;
  assign out_34_54 = t_r34_c54_12 >> 4;

  assign t_r34_c55_0 = p_33_55 << 1;
  assign t_r34_c55_1 = p_34_54 << 1;
  assign t_r34_c55_2 = p_34_55 << 2;
  assign t_r34_c55_3 = p_34_56 << 1;
  assign t_r34_c55_4 = p_35_55 << 1;
  assign t_r34_c55_5 = t_r34_c55_0 + p_33_54;
  assign t_r34_c55_6 = t_r34_c55_1 + p_33_56;
  assign t_r34_c55_7 = t_r34_c55_2 + t_r34_c55_3;
  assign t_r34_c55_8 = t_r34_c55_4 + p_35_54;
  assign t_r34_c55_9 = t_r34_c55_5 + t_r34_c55_6;
  assign t_r34_c55_10 = t_r34_c55_7 + t_r34_c55_8;
  assign t_r34_c55_11 = t_r34_c55_9 + t_r34_c55_10;
  assign t_r34_c55_12 = t_r34_c55_11 + p_35_56;
  assign out_34_55 = t_r34_c55_12 >> 4;

  assign t_r34_c56_0 = p_33_56 << 1;
  assign t_r34_c56_1 = p_34_55 << 1;
  assign t_r34_c56_2 = p_34_56 << 2;
  assign t_r34_c56_3 = p_34_57 << 1;
  assign t_r34_c56_4 = p_35_56 << 1;
  assign t_r34_c56_5 = t_r34_c56_0 + p_33_55;
  assign t_r34_c56_6 = t_r34_c56_1 + p_33_57;
  assign t_r34_c56_7 = t_r34_c56_2 + t_r34_c56_3;
  assign t_r34_c56_8 = t_r34_c56_4 + p_35_55;
  assign t_r34_c56_9 = t_r34_c56_5 + t_r34_c56_6;
  assign t_r34_c56_10 = t_r34_c56_7 + t_r34_c56_8;
  assign t_r34_c56_11 = t_r34_c56_9 + t_r34_c56_10;
  assign t_r34_c56_12 = t_r34_c56_11 + p_35_57;
  assign out_34_56 = t_r34_c56_12 >> 4;

  assign t_r34_c57_0 = p_33_57 << 1;
  assign t_r34_c57_1 = p_34_56 << 1;
  assign t_r34_c57_2 = p_34_57 << 2;
  assign t_r34_c57_3 = p_34_58 << 1;
  assign t_r34_c57_4 = p_35_57 << 1;
  assign t_r34_c57_5 = t_r34_c57_0 + p_33_56;
  assign t_r34_c57_6 = t_r34_c57_1 + p_33_58;
  assign t_r34_c57_7 = t_r34_c57_2 + t_r34_c57_3;
  assign t_r34_c57_8 = t_r34_c57_4 + p_35_56;
  assign t_r34_c57_9 = t_r34_c57_5 + t_r34_c57_6;
  assign t_r34_c57_10 = t_r34_c57_7 + t_r34_c57_8;
  assign t_r34_c57_11 = t_r34_c57_9 + t_r34_c57_10;
  assign t_r34_c57_12 = t_r34_c57_11 + p_35_58;
  assign out_34_57 = t_r34_c57_12 >> 4;

  assign t_r34_c58_0 = p_33_58 << 1;
  assign t_r34_c58_1 = p_34_57 << 1;
  assign t_r34_c58_2 = p_34_58 << 2;
  assign t_r34_c58_3 = p_34_59 << 1;
  assign t_r34_c58_4 = p_35_58 << 1;
  assign t_r34_c58_5 = t_r34_c58_0 + p_33_57;
  assign t_r34_c58_6 = t_r34_c58_1 + p_33_59;
  assign t_r34_c58_7 = t_r34_c58_2 + t_r34_c58_3;
  assign t_r34_c58_8 = t_r34_c58_4 + p_35_57;
  assign t_r34_c58_9 = t_r34_c58_5 + t_r34_c58_6;
  assign t_r34_c58_10 = t_r34_c58_7 + t_r34_c58_8;
  assign t_r34_c58_11 = t_r34_c58_9 + t_r34_c58_10;
  assign t_r34_c58_12 = t_r34_c58_11 + p_35_59;
  assign out_34_58 = t_r34_c58_12 >> 4;

  assign t_r34_c59_0 = p_33_59 << 1;
  assign t_r34_c59_1 = p_34_58 << 1;
  assign t_r34_c59_2 = p_34_59 << 2;
  assign t_r34_c59_3 = p_34_60 << 1;
  assign t_r34_c59_4 = p_35_59 << 1;
  assign t_r34_c59_5 = t_r34_c59_0 + p_33_58;
  assign t_r34_c59_6 = t_r34_c59_1 + p_33_60;
  assign t_r34_c59_7 = t_r34_c59_2 + t_r34_c59_3;
  assign t_r34_c59_8 = t_r34_c59_4 + p_35_58;
  assign t_r34_c59_9 = t_r34_c59_5 + t_r34_c59_6;
  assign t_r34_c59_10 = t_r34_c59_7 + t_r34_c59_8;
  assign t_r34_c59_11 = t_r34_c59_9 + t_r34_c59_10;
  assign t_r34_c59_12 = t_r34_c59_11 + p_35_60;
  assign out_34_59 = t_r34_c59_12 >> 4;

  assign t_r34_c60_0 = p_33_60 << 1;
  assign t_r34_c60_1 = p_34_59 << 1;
  assign t_r34_c60_2 = p_34_60 << 2;
  assign t_r34_c60_3 = p_34_61 << 1;
  assign t_r34_c60_4 = p_35_60 << 1;
  assign t_r34_c60_5 = t_r34_c60_0 + p_33_59;
  assign t_r34_c60_6 = t_r34_c60_1 + p_33_61;
  assign t_r34_c60_7 = t_r34_c60_2 + t_r34_c60_3;
  assign t_r34_c60_8 = t_r34_c60_4 + p_35_59;
  assign t_r34_c60_9 = t_r34_c60_5 + t_r34_c60_6;
  assign t_r34_c60_10 = t_r34_c60_7 + t_r34_c60_8;
  assign t_r34_c60_11 = t_r34_c60_9 + t_r34_c60_10;
  assign t_r34_c60_12 = t_r34_c60_11 + p_35_61;
  assign out_34_60 = t_r34_c60_12 >> 4;

  assign t_r34_c61_0 = p_33_61 << 1;
  assign t_r34_c61_1 = p_34_60 << 1;
  assign t_r34_c61_2 = p_34_61 << 2;
  assign t_r34_c61_3 = p_34_62 << 1;
  assign t_r34_c61_4 = p_35_61 << 1;
  assign t_r34_c61_5 = t_r34_c61_0 + p_33_60;
  assign t_r34_c61_6 = t_r34_c61_1 + p_33_62;
  assign t_r34_c61_7 = t_r34_c61_2 + t_r34_c61_3;
  assign t_r34_c61_8 = t_r34_c61_4 + p_35_60;
  assign t_r34_c61_9 = t_r34_c61_5 + t_r34_c61_6;
  assign t_r34_c61_10 = t_r34_c61_7 + t_r34_c61_8;
  assign t_r34_c61_11 = t_r34_c61_9 + t_r34_c61_10;
  assign t_r34_c61_12 = t_r34_c61_11 + p_35_62;
  assign out_34_61 = t_r34_c61_12 >> 4;

  assign t_r34_c62_0 = p_33_62 << 1;
  assign t_r34_c62_1 = p_34_61 << 1;
  assign t_r34_c62_2 = p_34_62 << 2;
  assign t_r34_c62_3 = p_34_63 << 1;
  assign t_r34_c62_4 = p_35_62 << 1;
  assign t_r34_c62_5 = t_r34_c62_0 + p_33_61;
  assign t_r34_c62_6 = t_r34_c62_1 + p_33_63;
  assign t_r34_c62_7 = t_r34_c62_2 + t_r34_c62_3;
  assign t_r34_c62_8 = t_r34_c62_4 + p_35_61;
  assign t_r34_c62_9 = t_r34_c62_5 + t_r34_c62_6;
  assign t_r34_c62_10 = t_r34_c62_7 + t_r34_c62_8;
  assign t_r34_c62_11 = t_r34_c62_9 + t_r34_c62_10;
  assign t_r34_c62_12 = t_r34_c62_11 + p_35_63;
  assign out_34_62 = t_r34_c62_12 >> 4;

  assign t_r34_c63_0 = p_33_63 << 1;
  assign t_r34_c63_1 = p_34_62 << 1;
  assign t_r34_c63_2 = p_34_63 << 2;
  assign t_r34_c63_3 = p_34_64 << 1;
  assign t_r34_c63_4 = p_35_63 << 1;
  assign t_r34_c63_5 = t_r34_c63_0 + p_33_62;
  assign t_r34_c63_6 = t_r34_c63_1 + p_33_64;
  assign t_r34_c63_7 = t_r34_c63_2 + t_r34_c63_3;
  assign t_r34_c63_8 = t_r34_c63_4 + p_35_62;
  assign t_r34_c63_9 = t_r34_c63_5 + t_r34_c63_6;
  assign t_r34_c63_10 = t_r34_c63_7 + t_r34_c63_8;
  assign t_r34_c63_11 = t_r34_c63_9 + t_r34_c63_10;
  assign t_r34_c63_12 = t_r34_c63_11 + p_35_64;
  assign out_34_63 = t_r34_c63_12 >> 4;

  assign t_r34_c64_0 = p_33_64 << 1;
  assign t_r34_c64_1 = p_34_63 << 1;
  assign t_r34_c64_2 = p_34_64 << 2;
  assign t_r34_c64_3 = p_34_65 << 1;
  assign t_r34_c64_4 = p_35_64 << 1;
  assign t_r34_c64_5 = t_r34_c64_0 + p_33_63;
  assign t_r34_c64_6 = t_r34_c64_1 + p_33_65;
  assign t_r34_c64_7 = t_r34_c64_2 + t_r34_c64_3;
  assign t_r34_c64_8 = t_r34_c64_4 + p_35_63;
  assign t_r34_c64_9 = t_r34_c64_5 + t_r34_c64_6;
  assign t_r34_c64_10 = t_r34_c64_7 + t_r34_c64_8;
  assign t_r34_c64_11 = t_r34_c64_9 + t_r34_c64_10;
  assign t_r34_c64_12 = t_r34_c64_11 + p_35_65;
  assign out_34_64 = t_r34_c64_12 >> 4;

  assign t_r35_c1_0 = p_34_1 << 1;
  assign t_r35_c1_1 = p_35_0 << 1;
  assign t_r35_c1_2 = p_35_1 << 2;
  assign t_r35_c1_3 = p_35_2 << 1;
  assign t_r35_c1_4 = p_36_1 << 1;
  assign t_r35_c1_5 = t_r35_c1_0 + p_34_0;
  assign t_r35_c1_6 = t_r35_c1_1 + p_34_2;
  assign t_r35_c1_7 = t_r35_c1_2 + t_r35_c1_3;
  assign t_r35_c1_8 = t_r35_c1_4 + p_36_0;
  assign t_r35_c1_9 = t_r35_c1_5 + t_r35_c1_6;
  assign t_r35_c1_10 = t_r35_c1_7 + t_r35_c1_8;
  assign t_r35_c1_11 = t_r35_c1_9 + t_r35_c1_10;
  assign t_r35_c1_12 = t_r35_c1_11 + p_36_2;
  assign out_35_1 = t_r35_c1_12 >> 4;

  assign t_r35_c2_0 = p_34_2 << 1;
  assign t_r35_c2_1 = p_35_1 << 1;
  assign t_r35_c2_2 = p_35_2 << 2;
  assign t_r35_c2_3 = p_35_3 << 1;
  assign t_r35_c2_4 = p_36_2 << 1;
  assign t_r35_c2_5 = t_r35_c2_0 + p_34_1;
  assign t_r35_c2_6 = t_r35_c2_1 + p_34_3;
  assign t_r35_c2_7 = t_r35_c2_2 + t_r35_c2_3;
  assign t_r35_c2_8 = t_r35_c2_4 + p_36_1;
  assign t_r35_c2_9 = t_r35_c2_5 + t_r35_c2_6;
  assign t_r35_c2_10 = t_r35_c2_7 + t_r35_c2_8;
  assign t_r35_c2_11 = t_r35_c2_9 + t_r35_c2_10;
  assign t_r35_c2_12 = t_r35_c2_11 + p_36_3;
  assign out_35_2 = t_r35_c2_12 >> 4;

  assign t_r35_c3_0 = p_34_3 << 1;
  assign t_r35_c3_1 = p_35_2 << 1;
  assign t_r35_c3_2 = p_35_3 << 2;
  assign t_r35_c3_3 = p_35_4 << 1;
  assign t_r35_c3_4 = p_36_3 << 1;
  assign t_r35_c3_5 = t_r35_c3_0 + p_34_2;
  assign t_r35_c3_6 = t_r35_c3_1 + p_34_4;
  assign t_r35_c3_7 = t_r35_c3_2 + t_r35_c3_3;
  assign t_r35_c3_8 = t_r35_c3_4 + p_36_2;
  assign t_r35_c3_9 = t_r35_c3_5 + t_r35_c3_6;
  assign t_r35_c3_10 = t_r35_c3_7 + t_r35_c3_8;
  assign t_r35_c3_11 = t_r35_c3_9 + t_r35_c3_10;
  assign t_r35_c3_12 = t_r35_c3_11 + p_36_4;
  assign out_35_3 = t_r35_c3_12 >> 4;

  assign t_r35_c4_0 = p_34_4 << 1;
  assign t_r35_c4_1 = p_35_3 << 1;
  assign t_r35_c4_2 = p_35_4 << 2;
  assign t_r35_c4_3 = p_35_5 << 1;
  assign t_r35_c4_4 = p_36_4 << 1;
  assign t_r35_c4_5 = t_r35_c4_0 + p_34_3;
  assign t_r35_c4_6 = t_r35_c4_1 + p_34_5;
  assign t_r35_c4_7 = t_r35_c4_2 + t_r35_c4_3;
  assign t_r35_c4_8 = t_r35_c4_4 + p_36_3;
  assign t_r35_c4_9 = t_r35_c4_5 + t_r35_c4_6;
  assign t_r35_c4_10 = t_r35_c4_7 + t_r35_c4_8;
  assign t_r35_c4_11 = t_r35_c4_9 + t_r35_c4_10;
  assign t_r35_c4_12 = t_r35_c4_11 + p_36_5;
  assign out_35_4 = t_r35_c4_12 >> 4;

  assign t_r35_c5_0 = p_34_5 << 1;
  assign t_r35_c5_1 = p_35_4 << 1;
  assign t_r35_c5_2 = p_35_5 << 2;
  assign t_r35_c5_3 = p_35_6 << 1;
  assign t_r35_c5_4 = p_36_5 << 1;
  assign t_r35_c5_5 = t_r35_c5_0 + p_34_4;
  assign t_r35_c5_6 = t_r35_c5_1 + p_34_6;
  assign t_r35_c5_7 = t_r35_c5_2 + t_r35_c5_3;
  assign t_r35_c5_8 = t_r35_c5_4 + p_36_4;
  assign t_r35_c5_9 = t_r35_c5_5 + t_r35_c5_6;
  assign t_r35_c5_10 = t_r35_c5_7 + t_r35_c5_8;
  assign t_r35_c5_11 = t_r35_c5_9 + t_r35_c5_10;
  assign t_r35_c5_12 = t_r35_c5_11 + p_36_6;
  assign out_35_5 = t_r35_c5_12 >> 4;

  assign t_r35_c6_0 = p_34_6 << 1;
  assign t_r35_c6_1 = p_35_5 << 1;
  assign t_r35_c6_2 = p_35_6 << 2;
  assign t_r35_c6_3 = p_35_7 << 1;
  assign t_r35_c6_4 = p_36_6 << 1;
  assign t_r35_c6_5 = t_r35_c6_0 + p_34_5;
  assign t_r35_c6_6 = t_r35_c6_1 + p_34_7;
  assign t_r35_c6_7 = t_r35_c6_2 + t_r35_c6_3;
  assign t_r35_c6_8 = t_r35_c6_4 + p_36_5;
  assign t_r35_c6_9 = t_r35_c6_5 + t_r35_c6_6;
  assign t_r35_c6_10 = t_r35_c6_7 + t_r35_c6_8;
  assign t_r35_c6_11 = t_r35_c6_9 + t_r35_c6_10;
  assign t_r35_c6_12 = t_r35_c6_11 + p_36_7;
  assign out_35_6 = t_r35_c6_12 >> 4;

  assign t_r35_c7_0 = p_34_7 << 1;
  assign t_r35_c7_1 = p_35_6 << 1;
  assign t_r35_c7_2 = p_35_7 << 2;
  assign t_r35_c7_3 = p_35_8 << 1;
  assign t_r35_c7_4 = p_36_7 << 1;
  assign t_r35_c7_5 = t_r35_c7_0 + p_34_6;
  assign t_r35_c7_6 = t_r35_c7_1 + p_34_8;
  assign t_r35_c7_7 = t_r35_c7_2 + t_r35_c7_3;
  assign t_r35_c7_8 = t_r35_c7_4 + p_36_6;
  assign t_r35_c7_9 = t_r35_c7_5 + t_r35_c7_6;
  assign t_r35_c7_10 = t_r35_c7_7 + t_r35_c7_8;
  assign t_r35_c7_11 = t_r35_c7_9 + t_r35_c7_10;
  assign t_r35_c7_12 = t_r35_c7_11 + p_36_8;
  assign out_35_7 = t_r35_c7_12 >> 4;

  assign t_r35_c8_0 = p_34_8 << 1;
  assign t_r35_c8_1 = p_35_7 << 1;
  assign t_r35_c8_2 = p_35_8 << 2;
  assign t_r35_c8_3 = p_35_9 << 1;
  assign t_r35_c8_4 = p_36_8 << 1;
  assign t_r35_c8_5 = t_r35_c8_0 + p_34_7;
  assign t_r35_c8_6 = t_r35_c8_1 + p_34_9;
  assign t_r35_c8_7 = t_r35_c8_2 + t_r35_c8_3;
  assign t_r35_c8_8 = t_r35_c8_4 + p_36_7;
  assign t_r35_c8_9 = t_r35_c8_5 + t_r35_c8_6;
  assign t_r35_c8_10 = t_r35_c8_7 + t_r35_c8_8;
  assign t_r35_c8_11 = t_r35_c8_9 + t_r35_c8_10;
  assign t_r35_c8_12 = t_r35_c8_11 + p_36_9;
  assign out_35_8 = t_r35_c8_12 >> 4;

  assign t_r35_c9_0 = p_34_9 << 1;
  assign t_r35_c9_1 = p_35_8 << 1;
  assign t_r35_c9_2 = p_35_9 << 2;
  assign t_r35_c9_3 = p_35_10 << 1;
  assign t_r35_c9_4 = p_36_9 << 1;
  assign t_r35_c9_5 = t_r35_c9_0 + p_34_8;
  assign t_r35_c9_6 = t_r35_c9_1 + p_34_10;
  assign t_r35_c9_7 = t_r35_c9_2 + t_r35_c9_3;
  assign t_r35_c9_8 = t_r35_c9_4 + p_36_8;
  assign t_r35_c9_9 = t_r35_c9_5 + t_r35_c9_6;
  assign t_r35_c9_10 = t_r35_c9_7 + t_r35_c9_8;
  assign t_r35_c9_11 = t_r35_c9_9 + t_r35_c9_10;
  assign t_r35_c9_12 = t_r35_c9_11 + p_36_10;
  assign out_35_9 = t_r35_c9_12 >> 4;

  assign t_r35_c10_0 = p_34_10 << 1;
  assign t_r35_c10_1 = p_35_9 << 1;
  assign t_r35_c10_2 = p_35_10 << 2;
  assign t_r35_c10_3 = p_35_11 << 1;
  assign t_r35_c10_4 = p_36_10 << 1;
  assign t_r35_c10_5 = t_r35_c10_0 + p_34_9;
  assign t_r35_c10_6 = t_r35_c10_1 + p_34_11;
  assign t_r35_c10_7 = t_r35_c10_2 + t_r35_c10_3;
  assign t_r35_c10_8 = t_r35_c10_4 + p_36_9;
  assign t_r35_c10_9 = t_r35_c10_5 + t_r35_c10_6;
  assign t_r35_c10_10 = t_r35_c10_7 + t_r35_c10_8;
  assign t_r35_c10_11 = t_r35_c10_9 + t_r35_c10_10;
  assign t_r35_c10_12 = t_r35_c10_11 + p_36_11;
  assign out_35_10 = t_r35_c10_12 >> 4;

  assign t_r35_c11_0 = p_34_11 << 1;
  assign t_r35_c11_1 = p_35_10 << 1;
  assign t_r35_c11_2 = p_35_11 << 2;
  assign t_r35_c11_3 = p_35_12 << 1;
  assign t_r35_c11_4 = p_36_11 << 1;
  assign t_r35_c11_5 = t_r35_c11_0 + p_34_10;
  assign t_r35_c11_6 = t_r35_c11_1 + p_34_12;
  assign t_r35_c11_7 = t_r35_c11_2 + t_r35_c11_3;
  assign t_r35_c11_8 = t_r35_c11_4 + p_36_10;
  assign t_r35_c11_9 = t_r35_c11_5 + t_r35_c11_6;
  assign t_r35_c11_10 = t_r35_c11_7 + t_r35_c11_8;
  assign t_r35_c11_11 = t_r35_c11_9 + t_r35_c11_10;
  assign t_r35_c11_12 = t_r35_c11_11 + p_36_12;
  assign out_35_11 = t_r35_c11_12 >> 4;

  assign t_r35_c12_0 = p_34_12 << 1;
  assign t_r35_c12_1 = p_35_11 << 1;
  assign t_r35_c12_2 = p_35_12 << 2;
  assign t_r35_c12_3 = p_35_13 << 1;
  assign t_r35_c12_4 = p_36_12 << 1;
  assign t_r35_c12_5 = t_r35_c12_0 + p_34_11;
  assign t_r35_c12_6 = t_r35_c12_1 + p_34_13;
  assign t_r35_c12_7 = t_r35_c12_2 + t_r35_c12_3;
  assign t_r35_c12_8 = t_r35_c12_4 + p_36_11;
  assign t_r35_c12_9 = t_r35_c12_5 + t_r35_c12_6;
  assign t_r35_c12_10 = t_r35_c12_7 + t_r35_c12_8;
  assign t_r35_c12_11 = t_r35_c12_9 + t_r35_c12_10;
  assign t_r35_c12_12 = t_r35_c12_11 + p_36_13;
  assign out_35_12 = t_r35_c12_12 >> 4;

  assign t_r35_c13_0 = p_34_13 << 1;
  assign t_r35_c13_1 = p_35_12 << 1;
  assign t_r35_c13_2 = p_35_13 << 2;
  assign t_r35_c13_3 = p_35_14 << 1;
  assign t_r35_c13_4 = p_36_13 << 1;
  assign t_r35_c13_5 = t_r35_c13_0 + p_34_12;
  assign t_r35_c13_6 = t_r35_c13_1 + p_34_14;
  assign t_r35_c13_7 = t_r35_c13_2 + t_r35_c13_3;
  assign t_r35_c13_8 = t_r35_c13_4 + p_36_12;
  assign t_r35_c13_9 = t_r35_c13_5 + t_r35_c13_6;
  assign t_r35_c13_10 = t_r35_c13_7 + t_r35_c13_8;
  assign t_r35_c13_11 = t_r35_c13_9 + t_r35_c13_10;
  assign t_r35_c13_12 = t_r35_c13_11 + p_36_14;
  assign out_35_13 = t_r35_c13_12 >> 4;

  assign t_r35_c14_0 = p_34_14 << 1;
  assign t_r35_c14_1 = p_35_13 << 1;
  assign t_r35_c14_2 = p_35_14 << 2;
  assign t_r35_c14_3 = p_35_15 << 1;
  assign t_r35_c14_4 = p_36_14 << 1;
  assign t_r35_c14_5 = t_r35_c14_0 + p_34_13;
  assign t_r35_c14_6 = t_r35_c14_1 + p_34_15;
  assign t_r35_c14_7 = t_r35_c14_2 + t_r35_c14_3;
  assign t_r35_c14_8 = t_r35_c14_4 + p_36_13;
  assign t_r35_c14_9 = t_r35_c14_5 + t_r35_c14_6;
  assign t_r35_c14_10 = t_r35_c14_7 + t_r35_c14_8;
  assign t_r35_c14_11 = t_r35_c14_9 + t_r35_c14_10;
  assign t_r35_c14_12 = t_r35_c14_11 + p_36_15;
  assign out_35_14 = t_r35_c14_12 >> 4;

  assign t_r35_c15_0 = p_34_15 << 1;
  assign t_r35_c15_1 = p_35_14 << 1;
  assign t_r35_c15_2 = p_35_15 << 2;
  assign t_r35_c15_3 = p_35_16 << 1;
  assign t_r35_c15_4 = p_36_15 << 1;
  assign t_r35_c15_5 = t_r35_c15_0 + p_34_14;
  assign t_r35_c15_6 = t_r35_c15_1 + p_34_16;
  assign t_r35_c15_7 = t_r35_c15_2 + t_r35_c15_3;
  assign t_r35_c15_8 = t_r35_c15_4 + p_36_14;
  assign t_r35_c15_9 = t_r35_c15_5 + t_r35_c15_6;
  assign t_r35_c15_10 = t_r35_c15_7 + t_r35_c15_8;
  assign t_r35_c15_11 = t_r35_c15_9 + t_r35_c15_10;
  assign t_r35_c15_12 = t_r35_c15_11 + p_36_16;
  assign out_35_15 = t_r35_c15_12 >> 4;

  assign t_r35_c16_0 = p_34_16 << 1;
  assign t_r35_c16_1 = p_35_15 << 1;
  assign t_r35_c16_2 = p_35_16 << 2;
  assign t_r35_c16_3 = p_35_17 << 1;
  assign t_r35_c16_4 = p_36_16 << 1;
  assign t_r35_c16_5 = t_r35_c16_0 + p_34_15;
  assign t_r35_c16_6 = t_r35_c16_1 + p_34_17;
  assign t_r35_c16_7 = t_r35_c16_2 + t_r35_c16_3;
  assign t_r35_c16_8 = t_r35_c16_4 + p_36_15;
  assign t_r35_c16_9 = t_r35_c16_5 + t_r35_c16_6;
  assign t_r35_c16_10 = t_r35_c16_7 + t_r35_c16_8;
  assign t_r35_c16_11 = t_r35_c16_9 + t_r35_c16_10;
  assign t_r35_c16_12 = t_r35_c16_11 + p_36_17;
  assign out_35_16 = t_r35_c16_12 >> 4;

  assign t_r35_c17_0 = p_34_17 << 1;
  assign t_r35_c17_1 = p_35_16 << 1;
  assign t_r35_c17_2 = p_35_17 << 2;
  assign t_r35_c17_3 = p_35_18 << 1;
  assign t_r35_c17_4 = p_36_17 << 1;
  assign t_r35_c17_5 = t_r35_c17_0 + p_34_16;
  assign t_r35_c17_6 = t_r35_c17_1 + p_34_18;
  assign t_r35_c17_7 = t_r35_c17_2 + t_r35_c17_3;
  assign t_r35_c17_8 = t_r35_c17_4 + p_36_16;
  assign t_r35_c17_9 = t_r35_c17_5 + t_r35_c17_6;
  assign t_r35_c17_10 = t_r35_c17_7 + t_r35_c17_8;
  assign t_r35_c17_11 = t_r35_c17_9 + t_r35_c17_10;
  assign t_r35_c17_12 = t_r35_c17_11 + p_36_18;
  assign out_35_17 = t_r35_c17_12 >> 4;

  assign t_r35_c18_0 = p_34_18 << 1;
  assign t_r35_c18_1 = p_35_17 << 1;
  assign t_r35_c18_2 = p_35_18 << 2;
  assign t_r35_c18_3 = p_35_19 << 1;
  assign t_r35_c18_4 = p_36_18 << 1;
  assign t_r35_c18_5 = t_r35_c18_0 + p_34_17;
  assign t_r35_c18_6 = t_r35_c18_1 + p_34_19;
  assign t_r35_c18_7 = t_r35_c18_2 + t_r35_c18_3;
  assign t_r35_c18_8 = t_r35_c18_4 + p_36_17;
  assign t_r35_c18_9 = t_r35_c18_5 + t_r35_c18_6;
  assign t_r35_c18_10 = t_r35_c18_7 + t_r35_c18_8;
  assign t_r35_c18_11 = t_r35_c18_9 + t_r35_c18_10;
  assign t_r35_c18_12 = t_r35_c18_11 + p_36_19;
  assign out_35_18 = t_r35_c18_12 >> 4;

  assign t_r35_c19_0 = p_34_19 << 1;
  assign t_r35_c19_1 = p_35_18 << 1;
  assign t_r35_c19_2 = p_35_19 << 2;
  assign t_r35_c19_3 = p_35_20 << 1;
  assign t_r35_c19_4 = p_36_19 << 1;
  assign t_r35_c19_5 = t_r35_c19_0 + p_34_18;
  assign t_r35_c19_6 = t_r35_c19_1 + p_34_20;
  assign t_r35_c19_7 = t_r35_c19_2 + t_r35_c19_3;
  assign t_r35_c19_8 = t_r35_c19_4 + p_36_18;
  assign t_r35_c19_9 = t_r35_c19_5 + t_r35_c19_6;
  assign t_r35_c19_10 = t_r35_c19_7 + t_r35_c19_8;
  assign t_r35_c19_11 = t_r35_c19_9 + t_r35_c19_10;
  assign t_r35_c19_12 = t_r35_c19_11 + p_36_20;
  assign out_35_19 = t_r35_c19_12 >> 4;

  assign t_r35_c20_0 = p_34_20 << 1;
  assign t_r35_c20_1 = p_35_19 << 1;
  assign t_r35_c20_2 = p_35_20 << 2;
  assign t_r35_c20_3 = p_35_21 << 1;
  assign t_r35_c20_4 = p_36_20 << 1;
  assign t_r35_c20_5 = t_r35_c20_0 + p_34_19;
  assign t_r35_c20_6 = t_r35_c20_1 + p_34_21;
  assign t_r35_c20_7 = t_r35_c20_2 + t_r35_c20_3;
  assign t_r35_c20_8 = t_r35_c20_4 + p_36_19;
  assign t_r35_c20_9 = t_r35_c20_5 + t_r35_c20_6;
  assign t_r35_c20_10 = t_r35_c20_7 + t_r35_c20_8;
  assign t_r35_c20_11 = t_r35_c20_9 + t_r35_c20_10;
  assign t_r35_c20_12 = t_r35_c20_11 + p_36_21;
  assign out_35_20 = t_r35_c20_12 >> 4;

  assign t_r35_c21_0 = p_34_21 << 1;
  assign t_r35_c21_1 = p_35_20 << 1;
  assign t_r35_c21_2 = p_35_21 << 2;
  assign t_r35_c21_3 = p_35_22 << 1;
  assign t_r35_c21_4 = p_36_21 << 1;
  assign t_r35_c21_5 = t_r35_c21_0 + p_34_20;
  assign t_r35_c21_6 = t_r35_c21_1 + p_34_22;
  assign t_r35_c21_7 = t_r35_c21_2 + t_r35_c21_3;
  assign t_r35_c21_8 = t_r35_c21_4 + p_36_20;
  assign t_r35_c21_9 = t_r35_c21_5 + t_r35_c21_6;
  assign t_r35_c21_10 = t_r35_c21_7 + t_r35_c21_8;
  assign t_r35_c21_11 = t_r35_c21_9 + t_r35_c21_10;
  assign t_r35_c21_12 = t_r35_c21_11 + p_36_22;
  assign out_35_21 = t_r35_c21_12 >> 4;

  assign t_r35_c22_0 = p_34_22 << 1;
  assign t_r35_c22_1 = p_35_21 << 1;
  assign t_r35_c22_2 = p_35_22 << 2;
  assign t_r35_c22_3 = p_35_23 << 1;
  assign t_r35_c22_4 = p_36_22 << 1;
  assign t_r35_c22_5 = t_r35_c22_0 + p_34_21;
  assign t_r35_c22_6 = t_r35_c22_1 + p_34_23;
  assign t_r35_c22_7 = t_r35_c22_2 + t_r35_c22_3;
  assign t_r35_c22_8 = t_r35_c22_4 + p_36_21;
  assign t_r35_c22_9 = t_r35_c22_5 + t_r35_c22_6;
  assign t_r35_c22_10 = t_r35_c22_7 + t_r35_c22_8;
  assign t_r35_c22_11 = t_r35_c22_9 + t_r35_c22_10;
  assign t_r35_c22_12 = t_r35_c22_11 + p_36_23;
  assign out_35_22 = t_r35_c22_12 >> 4;

  assign t_r35_c23_0 = p_34_23 << 1;
  assign t_r35_c23_1 = p_35_22 << 1;
  assign t_r35_c23_2 = p_35_23 << 2;
  assign t_r35_c23_3 = p_35_24 << 1;
  assign t_r35_c23_4 = p_36_23 << 1;
  assign t_r35_c23_5 = t_r35_c23_0 + p_34_22;
  assign t_r35_c23_6 = t_r35_c23_1 + p_34_24;
  assign t_r35_c23_7 = t_r35_c23_2 + t_r35_c23_3;
  assign t_r35_c23_8 = t_r35_c23_4 + p_36_22;
  assign t_r35_c23_9 = t_r35_c23_5 + t_r35_c23_6;
  assign t_r35_c23_10 = t_r35_c23_7 + t_r35_c23_8;
  assign t_r35_c23_11 = t_r35_c23_9 + t_r35_c23_10;
  assign t_r35_c23_12 = t_r35_c23_11 + p_36_24;
  assign out_35_23 = t_r35_c23_12 >> 4;

  assign t_r35_c24_0 = p_34_24 << 1;
  assign t_r35_c24_1 = p_35_23 << 1;
  assign t_r35_c24_2 = p_35_24 << 2;
  assign t_r35_c24_3 = p_35_25 << 1;
  assign t_r35_c24_4 = p_36_24 << 1;
  assign t_r35_c24_5 = t_r35_c24_0 + p_34_23;
  assign t_r35_c24_6 = t_r35_c24_1 + p_34_25;
  assign t_r35_c24_7 = t_r35_c24_2 + t_r35_c24_3;
  assign t_r35_c24_8 = t_r35_c24_4 + p_36_23;
  assign t_r35_c24_9 = t_r35_c24_5 + t_r35_c24_6;
  assign t_r35_c24_10 = t_r35_c24_7 + t_r35_c24_8;
  assign t_r35_c24_11 = t_r35_c24_9 + t_r35_c24_10;
  assign t_r35_c24_12 = t_r35_c24_11 + p_36_25;
  assign out_35_24 = t_r35_c24_12 >> 4;

  assign t_r35_c25_0 = p_34_25 << 1;
  assign t_r35_c25_1 = p_35_24 << 1;
  assign t_r35_c25_2 = p_35_25 << 2;
  assign t_r35_c25_3 = p_35_26 << 1;
  assign t_r35_c25_4 = p_36_25 << 1;
  assign t_r35_c25_5 = t_r35_c25_0 + p_34_24;
  assign t_r35_c25_6 = t_r35_c25_1 + p_34_26;
  assign t_r35_c25_7 = t_r35_c25_2 + t_r35_c25_3;
  assign t_r35_c25_8 = t_r35_c25_4 + p_36_24;
  assign t_r35_c25_9 = t_r35_c25_5 + t_r35_c25_6;
  assign t_r35_c25_10 = t_r35_c25_7 + t_r35_c25_8;
  assign t_r35_c25_11 = t_r35_c25_9 + t_r35_c25_10;
  assign t_r35_c25_12 = t_r35_c25_11 + p_36_26;
  assign out_35_25 = t_r35_c25_12 >> 4;

  assign t_r35_c26_0 = p_34_26 << 1;
  assign t_r35_c26_1 = p_35_25 << 1;
  assign t_r35_c26_2 = p_35_26 << 2;
  assign t_r35_c26_3 = p_35_27 << 1;
  assign t_r35_c26_4 = p_36_26 << 1;
  assign t_r35_c26_5 = t_r35_c26_0 + p_34_25;
  assign t_r35_c26_6 = t_r35_c26_1 + p_34_27;
  assign t_r35_c26_7 = t_r35_c26_2 + t_r35_c26_3;
  assign t_r35_c26_8 = t_r35_c26_4 + p_36_25;
  assign t_r35_c26_9 = t_r35_c26_5 + t_r35_c26_6;
  assign t_r35_c26_10 = t_r35_c26_7 + t_r35_c26_8;
  assign t_r35_c26_11 = t_r35_c26_9 + t_r35_c26_10;
  assign t_r35_c26_12 = t_r35_c26_11 + p_36_27;
  assign out_35_26 = t_r35_c26_12 >> 4;

  assign t_r35_c27_0 = p_34_27 << 1;
  assign t_r35_c27_1 = p_35_26 << 1;
  assign t_r35_c27_2 = p_35_27 << 2;
  assign t_r35_c27_3 = p_35_28 << 1;
  assign t_r35_c27_4 = p_36_27 << 1;
  assign t_r35_c27_5 = t_r35_c27_0 + p_34_26;
  assign t_r35_c27_6 = t_r35_c27_1 + p_34_28;
  assign t_r35_c27_7 = t_r35_c27_2 + t_r35_c27_3;
  assign t_r35_c27_8 = t_r35_c27_4 + p_36_26;
  assign t_r35_c27_9 = t_r35_c27_5 + t_r35_c27_6;
  assign t_r35_c27_10 = t_r35_c27_7 + t_r35_c27_8;
  assign t_r35_c27_11 = t_r35_c27_9 + t_r35_c27_10;
  assign t_r35_c27_12 = t_r35_c27_11 + p_36_28;
  assign out_35_27 = t_r35_c27_12 >> 4;

  assign t_r35_c28_0 = p_34_28 << 1;
  assign t_r35_c28_1 = p_35_27 << 1;
  assign t_r35_c28_2 = p_35_28 << 2;
  assign t_r35_c28_3 = p_35_29 << 1;
  assign t_r35_c28_4 = p_36_28 << 1;
  assign t_r35_c28_5 = t_r35_c28_0 + p_34_27;
  assign t_r35_c28_6 = t_r35_c28_1 + p_34_29;
  assign t_r35_c28_7 = t_r35_c28_2 + t_r35_c28_3;
  assign t_r35_c28_8 = t_r35_c28_4 + p_36_27;
  assign t_r35_c28_9 = t_r35_c28_5 + t_r35_c28_6;
  assign t_r35_c28_10 = t_r35_c28_7 + t_r35_c28_8;
  assign t_r35_c28_11 = t_r35_c28_9 + t_r35_c28_10;
  assign t_r35_c28_12 = t_r35_c28_11 + p_36_29;
  assign out_35_28 = t_r35_c28_12 >> 4;

  assign t_r35_c29_0 = p_34_29 << 1;
  assign t_r35_c29_1 = p_35_28 << 1;
  assign t_r35_c29_2 = p_35_29 << 2;
  assign t_r35_c29_3 = p_35_30 << 1;
  assign t_r35_c29_4 = p_36_29 << 1;
  assign t_r35_c29_5 = t_r35_c29_0 + p_34_28;
  assign t_r35_c29_6 = t_r35_c29_1 + p_34_30;
  assign t_r35_c29_7 = t_r35_c29_2 + t_r35_c29_3;
  assign t_r35_c29_8 = t_r35_c29_4 + p_36_28;
  assign t_r35_c29_9 = t_r35_c29_5 + t_r35_c29_6;
  assign t_r35_c29_10 = t_r35_c29_7 + t_r35_c29_8;
  assign t_r35_c29_11 = t_r35_c29_9 + t_r35_c29_10;
  assign t_r35_c29_12 = t_r35_c29_11 + p_36_30;
  assign out_35_29 = t_r35_c29_12 >> 4;

  assign t_r35_c30_0 = p_34_30 << 1;
  assign t_r35_c30_1 = p_35_29 << 1;
  assign t_r35_c30_2 = p_35_30 << 2;
  assign t_r35_c30_3 = p_35_31 << 1;
  assign t_r35_c30_4 = p_36_30 << 1;
  assign t_r35_c30_5 = t_r35_c30_0 + p_34_29;
  assign t_r35_c30_6 = t_r35_c30_1 + p_34_31;
  assign t_r35_c30_7 = t_r35_c30_2 + t_r35_c30_3;
  assign t_r35_c30_8 = t_r35_c30_4 + p_36_29;
  assign t_r35_c30_9 = t_r35_c30_5 + t_r35_c30_6;
  assign t_r35_c30_10 = t_r35_c30_7 + t_r35_c30_8;
  assign t_r35_c30_11 = t_r35_c30_9 + t_r35_c30_10;
  assign t_r35_c30_12 = t_r35_c30_11 + p_36_31;
  assign out_35_30 = t_r35_c30_12 >> 4;

  assign t_r35_c31_0 = p_34_31 << 1;
  assign t_r35_c31_1 = p_35_30 << 1;
  assign t_r35_c31_2 = p_35_31 << 2;
  assign t_r35_c31_3 = p_35_32 << 1;
  assign t_r35_c31_4 = p_36_31 << 1;
  assign t_r35_c31_5 = t_r35_c31_0 + p_34_30;
  assign t_r35_c31_6 = t_r35_c31_1 + p_34_32;
  assign t_r35_c31_7 = t_r35_c31_2 + t_r35_c31_3;
  assign t_r35_c31_8 = t_r35_c31_4 + p_36_30;
  assign t_r35_c31_9 = t_r35_c31_5 + t_r35_c31_6;
  assign t_r35_c31_10 = t_r35_c31_7 + t_r35_c31_8;
  assign t_r35_c31_11 = t_r35_c31_9 + t_r35_c31_10;
  assign t_r35_c31_12 = t_r35_c31_11 + p_36_32;
  assign out_35_31 = t_r35_c31_12 >> 4;

  assign t_r35_c32_0 = p_34_32 << 1;
  assign t_r35_c32_1 = p_35_31 << 1;
  assign t_r35_c32_2 = p_35_32 << 2;
  assign t_r35_c32_3 = p_35_33 << 1;
  assign t_r35_c32_4 = p_36_32 << 1;
  assign t_r35_c32_5 = t_r35_c32_0 + p_34_31;
  assign t_r35_c32_6 = t_r35_c32_1 + p_34_33;
  assign t_r35_c32_7 = t_r35_c32_2 + t_r35_c32_3;
  assign t_r35_c32_8 = t_r35_c32_4 + p_36_31;
  assign t_r35_c32_9 = t_r35_c32_5 + t_r35_c32_6;
  assign t_r35_c32_10 = t_r35_c32_7 + t_r35_c32_8;
  assign t_r35_c32_11 = t_r35_c32_9 + t_r35_c32_10;
  assign t_r35_c32_12 = t_r35_c32_11 + p_36_33;
  assign out_35_32 = t_r35_c32_12 >> 4;

  assign t_r35_c33_0 = p_34_33 << 1;
  assign t_r35_c33_1 = p_35_32 << 1;
  assign t_r35_c33_2 = p_35_33 << 2;
  assign t_r35_c33_3 = p_35_34 << 1;
  assign t_r35_c33_4 = p_36_33 << 1;
  assign t_r35_c33_5 = t_r35_c33_0 + p_34_32;
  assign t_r35_c33_6 = t_r35_c33_1 + p_34_34;
  assign t_r35_c33_7 = t_r35_c33_2 + t_r35_c33_3;
  assign t_r35_c33_8 = t_r35_c33_4 + p_36_32;
  assign t_r35_c33_9 = t_r35_c33_5 + t_r35_c33_6;
  assign t_r35_c33_10 = t_r35_c33_7 + t_r35_c33_8;
  assign t_r35_c33_11 = t_r35_c33_9 + t_r35_c33_10;
  assign t_r35_c33_12 = t_r35_c33_11 + p_36_34;
  assign out_35_33 = t_r35_c33_12 >> 4;

  assign t_r35_c34_0 = p_34_34 << 1;
  assign t_r35_c34_1 = p_35_33 << 1;
  assign t_r35_c34_2 = p_35_34 << 2;
  assign t_r35_c34_3 = p_35_35 << 1;
  assign t_r35_c34_4 = p_36_34 << 1;
  assign t_r35_c34_5 = t_r35_c34_0 + p_34_33;
  assign t_r35_c34_6 = t_r35_c34_1 + p_34_35;
  assign t_r35_c34_7 = t_r35_c34_2 + t_r35_c34_3;
  assign t_r35_c34_8 = t_r35_c34_4 + p_36_33;
  assign t_r35_c34_9 = t_r35_c34_5 + t_r35_c34_6;
  assign t_r35_c34_10 = t_r35_c34_7 + t_r35_c34_8;
  assign t_r35_c34_11 = t_r35_c34_9 + t_r35_c34_10;
  assign t_r35_c34_12 = t_r35_c34_11 + p_36_35;
  assign out_35_34 = t_r35_c34_12 >> 4;

  assign t_r35_c35_0 = p_34_35 << 1;
  assign t_r35_c35_1 = p_35_34 << 1;
  assign t_r35_c35_2 = p_35_35 << 2;
  assign t_r35_c35_3 = p_35_36 << 1;
  assign t_r35_c35_4 = p_36_35 << 1;
  assign t_r35_c35_5 = t_r35_c35_0 + p_34_34;
  assign t_r35_c35_6 = t_r35_c35_1 + p_34_36;
  assign t_r35_c35_7 = t_r35_c35_2 + t_r35_c35_3;
  assign t_r35_c35_8 = t_r35_c35_4 + p_36_34;
  assign t_r35_c35_9 = t_r35_c35_5 + t_r35_c35_6;
  assign t_r35_c35_10 = t_r35_c35_7 + t_r35_c35_8;
  assign t_r35_c35_11 = t_r35_c35_9 + t_r35_c35_10;
  assign t_r35_c35_12 = t_r35_c35_11 + p_36_36;
  assign out_35_35 = t_r35_c35_12 >> 4;

  assign t_r35_c36_0 = p_34_36 << 1;
  assign t_r35_c36_1 = p_35_35 << 1;
  assign t_r35_c36_2 = p_35_36 << 2;
  assign t_r35_c36_3 = p_35_37 << 1;
  assign t_r35_c36_4 = p_36_36 << 1;
  assign t_r35_c36_5 = t_r35_c36_0 + p_34_35;
  assign t_r35_c36_6 = t_r35_c36_1 + p_34_37;
  assign t_r35_c36_7 = t_r35_c36_2 + t_r35_c36_3;
  assign t_r35_c36_8 = t_r35_c36_4 + p_36_35;
  assign t_r35_c36_9 = t_r35_c36_5 + t_r35_c36_6;
  assign t_r35_c36_10 = t_r35_c36_7 + t_r35_c36_8;
  assign t_r35_c36_11 = t_r35_c36_9 + t_r35_c36_10;
  assign t_r35_c36_12 = t_r35_c36_11 + p_36_37;
  assign out_35_36 = t_r35_c36_12 >> 4;

  assign t_r35_c37_0 = p_34_37 << 1;
  assign t_r35_c37_1 = p_35_36 << 1;
  assign t_r35_c37_2 = p_35_37 << 2;
  assign t_r35_c37_3 = p_35_38 << 1;
  assign t_r35_c37_4 = p_36_37 << 1;
  assign t_r35_c37_5 = t_r35_c37_0 + p_34_36;
  assign t_r35_c37_6 = t_r35_c37_1 + p_34_38;
  assign t_r35_c37_7 = t_r35_c37_2 + t_r35_c37_3;
  assign t_r35_c37_8 = t_r35_c37_4 + p_36_36;
  assign t_r35_c37_9 = t_r35_c37_5 + t_r35_c37_6;
  assign t_r35_c37_10 = t_r35_c37_7 + t_r35_c37_8;
  assign t_r35_c37_11 = t_r35_c37_9 + t_r35_c37_10;
  assign t_r35_c37_12 = t_r35_c37_11 + p_36_38;
  assign out_35_37 = t_r35_c37_12 >> 4;

  assign t_r35_c38_0 = p_34_38 << 1;
  assign t_r35_c38_1 = p_35_37 << 1;
  assign t_r35_c38_2 = p_35_38 << 2;
  assign t_r35_c38_3 = p_35_39 << 1;
  assign t_r35_c38_4 = p_36_38 << 1;
  assign t_r35_c38_5 = t_r35_c38_0 + p_34_37;
  assign t_r35_c38_6 = t_r35_c38_1 + p_34_39;
  assign t_r35_c38_7 = t_r35_c38_2 + t_r35_c38_3;
  assign t_r35_c38_8 = t_r35_c38_4 + p_36_37;
  assign t_r35_c38_9 = t_r35_c38_5 + t_r35_c38_6;
  assign t_r35_c38_10 = t_r35_c38_7 + t_r35_c38_8;
  assign t_r35_c38_11 = t_r35_c38_9 + t_r35_c38_10;
  assign t_r35_c38_12 = t_r35_c38_11 + p_36_39;
  assign out_35_38 = t_r35_c38_12 >> 4;

  assign t_r35_c39_0 = p_34_39 << 1;
  assign t_r35_c39_1 = p_35_38 << 1;
  assign t_r35_c39_2 = p_35_39 << 2;
  assign t_r35_c39_3 = p_35_40 << 1;
  assign t_r35_c39_4 = p_36_39 << 1;
  assign t_r35_c39_5 = t_r35_c39_0 + p_34_38;
  assign t_r35_c39_6 = t_r35_c39_1 + p_34_40;
  assign t_r35_c39_7 = t_r35_c39_2 + t_r35_c39_3;
  assign t_r35_c39_8 = t_r35_c39_4 + p_36_38;
  assign t_r35_c39_9 = t_r35_c39_5 + t_r35_c39_6;
  assign t_r35_c39_10 = t_r35_c39_7 + t_r35_c39_8;
  assign t_r35_c39_11 = t_r35_c39_9 + t_r35_c39_10;
  assign t_r35_c39_12 = t_r35_c39_11 + p_36_40;
  assign out_35_39 = t_r35_c39_12 >> 4;

  assign t_r35_c40_0 = p_34_40 << 1;
  assign t_r35_c40_1 = p_35_39 << 1;
  assign t_r35_c40_2 = p_35_40 << 2;
  assign t_r35_c40_3 = p_35_41 << 1;
  assign t_r35_c40_4 = p_36_40 << 1;
  assign t_r35_c40_5 = t_r35_c40_0 + p_34_39;
  assign t_r35_c40_6 = t_r35_c40_1 + p_34_41;
  assign t_r35_c40_7 = t_r35_c40_2 + t_r35_c40_3;
  assign t_r35_c40_8 = t_r35_c40_4 + p_36_39;
  assign t_r35_c40_9 = t_r35_c40_5 + t_r35_c40_6;
  assign t_r35_c40_10 = t_r35_c40_7 + t_r35_c40_8;
  assign t_r35_c40_11 = t_r35_c40_9 + t_r35_c40_10;
  assign t_r35_c40_12 = t_r35_c40_11 + p_36_41;
  assign out_35_40 = t_r35_c40_12 >> 4;

  assign t_r35_c41_0 = p_34_41 << 1;
  assign t_r35_c41_1 = p_35_40 << 1;
  assign t_r35_c41_2 = p_35_41 << 2;
  assign t_r35_c41_3 = p_35_42 << 1;
  assign t_r35_c41_4 = p_36_41 << 1;
  assign t_r35_c41_5 = t_r35_c41_0 + p_34_40;
  assign t_r35_c41_6 = t_r35_c41_1 + p_34_42;
  assign t_r35_c41_7 = t_r35_c41_2 + t_r35_c41_3;
  assign t_r35_c41_8 = t_r35_c41_4 + p_36_40;
  assign t_r35_c41_9 = t_r35_c41_5 + t_r35_c41_6;
  assign t_r35_c41_10 = t_r35_c41_7 + t_r35_c41_8;
  assign t_r35_c41_11 = t_r35_c41_9 + t_r35_c41_10;
  assign t_r35_c41_12 = t_r35_c41_11 + p_36_42;
  assign out_35_41 = t_r35_c41_12 >> 4;

  assign t_r35_c42_0 = p_34_42 << 1;
  assign t_r35_c42_1 = p_35_41 << 1;
  assign t_r35_c42_2 = p_35_42 << 2;
  assign t_r35_c42_3 = p_35_43 << 1;
  assign t_r35_c42_4 = p_36_42 << 1;
  assign t_r35_c42_5 = t_r35_c42_0 + p_34_41;
  assign t_r35_c42_6 = t_r35_c42_1 + p_34_43;
  assign t_r35_c42_7 = t_r35_c42_2 + t_r35_c42_3;
  assign t_r35_c42_8 = t_r35_c42_4 + p_36_41;
  assign t_r35_c42_9 = t_r35_c42_5 + t_r35_c42_6;
  assign t_r35_c42_10 = t_r35_c42_7 + t_r35_c42_8;
  assign t_r35_c42_11 = t_r35_c42_9 + t_r35_c42_10;
  assign t_r35_c42_12 = t_r35_c42_11 + p_36_43;
  assign out_35_42 = t_r35_c42_12 >> 4;

  assign t_r35_c43_0 = p_34_43 << 1;
  assign t_r35_c43_1 = p_35_42 << 1;
  assign t_r35_c43_2 = p_35_43 << 2;
  assign t_r35_c43_3 = p_35_44 << 1;
  assign t_r35_c43_4 = p_36_43 << 1;
  assign t_r35_c43_5 = t_r35_c43_0 + p_34_42;
  assign t_r35_c43_6 = t_r35_c43_1 + p_34_44;
  assign t_r35_c43_7 = t_r35_c43_2 + t_r35_c43_3;
  assign t_r35_c43_8 = t_r35_c43_4 + p_36_42;
  assign t_r35_c43_9 = t_r35_c43_5 + t_r35_c43_6;
  assign t_r35_c43_10 = t_r35_c43_7 + t_r35_c43_8;
  assign t_r35_c43_11 = t_r35_c43_9 + t_r35_c43_10;
  assign t_r35_c43_12 = t_r35_c43_11 + p_36_44;
  assign out_35_43 = t_r35_c43_12 >> 4;

  assign t_r35_c44_0 = p_34_44 << 1;
  assign t_r35_c44_1 = p_35_43 << 1;
  assign t_r35_c44_2 = p_35_44 << 2;
  assign t_r35_c44_3 = p_35_45 << 1;
  assign t_r35_c44_4 = p_36_44 << 1;
  assign t_r35_c44_5 = t_r35_c44_0 + p_34_43;
  assign t_r35_c44_6 = t_r35_c44_1 + p_34_45;
  assign t_r35_c44_7 = t_r35_c44_2 + t_r35_c44_3;
  assign t_r35_c44_8 = t_r35_c44_4 + p_36_43;
  assign t_r35_c44_9 = t_r35_c44_5 + t_r35_c44_6;
  assign t_r35_c44_10 = t_r35_c44_7 + t_r35_c44_8;
  assign t_r35_c44_11 = t_r35_c44_9 + t_r35_c44_10;
  assign t_r35_c44_12 = t_r35_c44_11 + p_36_45;
  assign out_35_44 = t_r35_c44_12 >> 4;

  assign t_r35_c45_0 = p_34_45 << 1;
  assign t_r35_c45_1 = p_35_44 << 1;
  assign t_r35_c45_2 = p_35_45 << 2;
  assign t_r35_c45_3 = p_35_46 << 1;
  assign t_r35_c45_4 = p_36_45 << 1;
  assign t_r35_c45_5 = t_r35_c45_0 + p_34_44;
  assign t_r35_c45_6 = t_r35_c45_1 + p_34_46;
  assign t_r35_c45_7 = t_r35_c45_2 + t_r35_c45_3;
  assign t_r35_c45_8 = t_r35_c45_4 + p_36_44;
  assign t_r35_c45_9 = t_r35_c45_5 + t_r35_c45_6;
  assign t_r35_c45_10 = t_r35_c45_7 + t_r35_c45_8;
  assign t_r35_c45_11 = t_r35_c45_9 + t_r35_c45_10;
  assign t_r35_c45_12 = t_r35_c45_11 + p_36_46;
  assign out_35_45 = t_r35_c45_12 >> 4;

  assign t_r35_c46_0 = p_34_46 << 1;
  assign t_r35_c46_1 = p_35_45 << 1;
  assign t_r35_c46_2 = p_35_46 << 2;
  assign t_r35_c46_3 = p_35_47 << 1;
  assign t_r35_c46_4 = p_36_46 << 1;
  assign t_r35_c46_5 = t_r35_c46_0 + p_34_45;
  assign t_r35_c46_6 = t_r35_c46_1 + p_34_47;
  assign t_r35_c46_7 = t_r35_c46_2 + t_r35_c46_3;
  assign t_r35_c46_8 = t_r35_c46_4 + p_36_45;
  assign t_r35_c46_9 = t_r35_c46_5 + t_r35_c46_6;
  assign t_r35_c46_10 = t_r35_c46_7 + t_r35_c46_8;
  assign t_r35_c46_11 = t_r35_c46_9 + t_r35_c46_10;
  assign t_r35_c46_12 = t_r35_c46_11 + p_36_47;
  assign out_35_46 = t_r35_c46_12 >> 4;

  assign t_r35_c47_0 = p_34_47 << 1;
  assign t_r35_c47_1 = p_35_46 << 1;
  assign t_r35_c47_2 = p_35_47 << 2;
  assign t_r35_c47_3 = p_35_48 << 1;
  assign t_r35_c47_4 = p_36_47 << 1;
  assign t_r35_c47_5 = t_r35_c47_0 + p_34_46;
  assign t_r35_c47_6 = t_r35_c47_1 + p_34_48;
  assign t_r35_c47_7 = t_r35_c47_2 + t_r35_c47_3;
  assign t_r35_c47_8 = t_r35_c47_4 + p_36_46;
  assign t_r35_c47_9 = t_r35_c47_5 + t_r35_c47_6;
  assign t_r35_c47_10 = t_r35_c47_7 + t_r35_c47_8;
  assign t_r35_c47_11 = t_r35_c47_9 + t_r35_c47_10;
  assign t_r35_c47_12 = t_r35_c47_11 + p_36_48;
  assign out_35_47 = t_r35_c47_12 >> 4;

  assign t_r35_c48_0 = p_34_48 << 1;
  assign t_r35_c48_1 = p_35_47 << 1;
  assign t_r35_c48_2 = p_35_48 << 2;
  assign t_r35_c48_3 = p_35_49 << 1;
  assign t_r35_c48_4 = p_36_48 << 1;
  assign t_r35_c48_5 = t_r35_c48_0 + p_34_47;
  assign t_r35_c48_6 = t_r35_c48_1 + p_34_49;
  assign t_r35_c48_7 = t_r35_c48_2 + t_r35_c48_3;
  assign t_r35_c48_8 = t_r35_c48_4 + p_36_47;
  assign t_r35_c48_9 = t_r35_c48_5 + t_r35_c48_6;
  assign t_r35_c48_10 = t_r35_c48_7 + t_r35_c48_8;
  assign t_r35_c48_11 = t_r35_c48_9 + t_r35_c48_10;
  assign t_r35_c48_12 = t_r35_c48_11 + p_36_49;
  assign out_35_48 = t_r35_c48_12 >> 4;

  assign t_r35_c49_0 = p_34_49 << 1;
  assign t_r35_c49_1 = p_35_48 << 1;
  assign t_r35_c49_2 = p_35_49 << 2;
  assign t_r35_c49_3 = p_35_50 << 1;
  assign t_r35_c49_4 = p_36_49 << 1;
  assign t_r35_c49_5 = t_r35_c49_0 + p_34_48;
  assign t_r35_c49_6 = t_r35_c49_1 + p_34_50;
  assign t_r35_c49_7 = t_r35_c49_2 + t_r35_c49_3;
  assign t_r35_c49_8 = t_r35_c49_4 + p_36_48;
  assign t_r35_c49_9 = t_r35_c49_5 + t_r35_c49_6;
  assign t_r35_c49_10 = t_r35_c49_7 + t_r35_c49_8;
  assign t_r35_c49_11 = t_r35_c49_9 + t_r35_c49_10;
  assign t_r35_c49_12 = t_r35_c49_11 + p_36_50;
  assign out_35_49 = t_r35_c49_12 >> 4;

  assign t_r35_c50_0 = p_34_50 << 1;
  assign t_r35_c50_1 = p_35_49 << 1;
  assign t_r35_c50_2 = p_35_50 << 2;
  assign t_r35_c50_3 = p_35_51 << 1;
  assign t_r35_c50_4 = p_36_50 << 1;
  assign t_r35_c50_5 = t_r35_c50_0 + p_34_49;
  assign t_r35_c50_6 = t_r35_c50_1 + p_34_51;
  assign t_r35_c50_7 = t_r35_c50_2 + t_r35_c50_3;
  assign t_r35_c50_8 = t_r35_c50_4 + p_36_49;
  assign t_r35_c50_9 = t_r35_c50_5 + t_r35_c50_6;
  assign t_r35_c50_10 = t_r35_c50_7 + t_r35_c50_8;
  assign t_r35_c50_11 = t_r35_c50_9 + t_r35_c50_10;
  assign t_r35_c50_12 = t_r35_c50_11 + p_36_51;
  assign out_35_50 = t_r35_c50_12 >> 4;

  assign t_r35_c51_0 = p_34_51 << 1;
  assign t_r35_c51_1 = p_35_50 << 1;
  assign t_r35_c51_2 = p_35_51 << 2;
  assign t_r35_c51_3 = p_35_52 << 1;
  assign t_r35_c51_4 = p_36_51 << 1;
  assign t_r35_c51_5 = t_r35_c51_0 + p_34_50;
  assign t_r35_c51_6 = t_r35_c51_1 + p_34_52;
  assign t_r35_c51_7 = t_r35_c51_2 + t_r35_c51_3;
  assign t_r35_c51_8 = t_r35_c51_4 + p_36_50;
  assign t_r35_c51_9 = t_r35_c51_5 + t_r35_c51_6;
  assign t_r35_c51_10 = t_r35_c51_7 + t_r35_c51_8;
  assign t_r35_c51_11 = t_r35_c51_9 + t_r35_c51_10;
  assign t_r35_c51_12 = t_r35_c51_11 + p_36_52;
  assign out_35_51 = t_r35_c51_12 >> 4;

  assign t_r35_c52_0 = p_34_52 << 1;
  assign t_r35_c52_1 = p_35_51 << 1;
  assign t_r35_c52_2 = p_35_52 << 2;
  assign t_r35_c52_3 = p_35_53 << 1;
  assign t_r35_c52_4 = p_36_52 << 1;
  assign t_r35_c52_5 = t_r35_c52_0 + p_34_51;
  assign t_r35_c52_6 = t_r35_c52_1 + p_34_53;
  assign t_r35_c52_7 = t_r35_c52_2 + t_r35_c52_3;
  assign t_r35_c52_8 = t_r35_c52_4 + p_36_51;
  assign t_r35_c52_9 = t_r35_c52_5 + t_r35_c52_6;
  assign t_r35_c52_10 = t_r35_c52_7 + t_r35_c52_8;
  assign t_r35_c52_11 = t_r35_c52_9 + t_r35_c52_10;
  assign t_r35_c52_12 = t_r35_c52_11 + p_36_53;
  assign out_35_52 = t_r35_c52_12 >> 4;

  assign t_r35_c53_0 = p_34_53 << 1;
  assign t_r35_c53_1 = p_35_52 << 1;
  assign t_r35_c53_2 = p_35_53 << 2;
  assign t_r35_c53_3 = p_35_54 << 1;
  assign t_r35_c53_4 = p_36_53 << 1;
  assign t_r35_c53_5 = t_r35_c53_0 + p_34_52;
  assign t_r35_c53_6 = t_r35_c53_1 + p_34_54;
  assign t_r35_c53_7 = t_r35_c53_2 + t_r35_c53_3;
  assign t_r35_c53_8 = t_r35_c53_4 + p_36_52;
  assign t_r35_c53_9 = t_r35_c53_5 + t_r35_c53_6;
  assign t_r35_c53_10 = t_r35_c53_7 + t_r35_c53_8;
  assign t_r35_c53_11 = t_r35_c53_9 + t_r35_c53_10;
  assign t_r35_c53_12 = t_r35_c53_11 + p_36_54;
  assign out_35_53 = t_r35_c53_12 >> 4;

  assign t_r35_c54_0 = p_34_54 << 1;
  assign t_r35_c54_1 = p_35_53 << 1;
  assign t_r35_c54_2 = p_35_54 << 2;
  assign t_r35_c54_3 = p_35_55 << 1;
  assign t_r35_c54_4 = p_36_54 << 1;
  assign t_r35_c54_5 = t_r35_c54_0 + p_34_53;
  assign t_r35_c54_6 = t_r35_c54_1 + p_34_55;
  assign t_r35_c54_7 = t_r35_c54_2 + t_r35_c54_3;
  assign t_r35_c54_8 = t_r35_c54_4 + p_36_53;
  assign t_r35_c54_9 = t_r35_c54_5 + t_r35_c54_6;
  assign t_r35_c54_10 = t_r35_c54_7 + t_r35_c54_8;
  assign t_r35_c54_11 = t_r35_c54_9 + t_r35_c54_10;
  assign t_r35_c54_12 = t_r35_c54_11 + p_36_55;
  assign out_35_54 = t_r35_c54_12 >> 4;

  assign t_r35_c55_0 = p_34_55 << 1;
  assign t_r35_c55_1 = p_35_54 << 1;
  assign t_r35_c55_2 = p_35_55 << 2;
  assign t_r35_c55_3 = p_35_56 << 1;
  assign t_r35_c55_4 = p_36_55 << 1;
  assign t_r35_c55_5 = t_r35_c55_0 + p_34_54;
  assign t_r35_c55_6 = t_r35_c55_1 + p_34_56;
  assign t_r35_c55_7 = t_r35_c55_2 + t_r35_c55_3;
  assign t_r35_c55_8 = t_r35_c55_4 + p_36_54;
  assign t_r35_c55_9 = t_r35_c55_5 + t_r35_c55_6;
  assign t_r35_c55_10 = t_r35_c55_7 + t_r35_c55_8;
  assign t_r35_c55_11 = t_r35_c55_9 + t_r35_c55_10;
  assign t_r35_c55_12 = t_r35_c55_11 + p_36_56;
  assign out_35_55 = t_r35_c55_12 >> 4;

  assign t_r35_c56_0 = p_34_56 << 1;
  assign t_r35_c56_1 = p_35_55 << 1;
  assign t_r35_c56_2 = p_35_56 << 2;
  assign t_r35_c56_3 = p_35_57 << 1;
  assign t_r35_c56_4 = p_36_56 << 1;
  assign t_r35_c56_5 = t_r35_c56_0 + p_34_55;
  assign t_r35_c56_6 = t_r35_c56_1 + p_34_57;
  assign t_r35_c56_7 = t_r35_c56_2 + t_r35_c56_3;
  assign t_r35_c56_8 = t_r35_c56_4 + p_36_55;
  assign t_r35_c56_9 = t_r35_c56_5 + t_r35_c56_6;
  assign t_r35_c56_10 = t_r35_c56_7 + t_r35_c56_8;
  assign t_r35_c56_11 = t_r35_c56_9 + t_r35_c56_10;
  assign t_r35_c56_12 = t_r35_c56_11 + p_36_57;
  assign out_35_56 = t_r35_c56_12 >> 4;

  assign t_r35_c57_0 = p_34_57 << 1;
  assign t_r35_c57_1 = p_35_56 << 1;
  assign t_r35_c57_2 = p_35_57 << 2;
  assign t_r35_c57_3 = p_35_58 << 1;
  assign t_r35_c57_4 = p_36_57 << 1;
  assign t_r35_c57_5 = t_r35_c57_0 + p_34_56;
  assign t_r35_c57_6 = t_r35_c57_1 + p_34_58;
  assign t_r35_c57_7 = t_r35_c57_2 + t_r35_c57_3;
  assign t_r35_c57_8 = t_r35_c57_4 + p_36_56;
  assign t_r35_c57_9 = t_r35_c57_5 + t_r35_c57_6;
  assign t_r35_c57_10 = t_r35_c57_7 + t_r35_c57_8;
  assign t_r35_c57_11 = t_r35_c57_9 + t_r35_c57_10;
  assign t_r35_c57_12 = t_r35_c57_11 + p_36_58;
  assign out_35_57 = t_r35_c57_12 >> 4;

  assign t_r35_c58_0 = p_34_58 << 1;
  assign t_r35_c58_1 = p_35_57 << 1;
  assign t_r35_c58_2 = p_35_58 << 2;
  assign t_r35_c58_3 = p_35_59 << 1;
  assign t_r35_c58_4 = p_36_58 << 1;
  assign t_r35_c58_5 = t_r35_c58_0 + p_34_57;
  assign t_r35_c58_6 = t_r35_c58_1 + p_34_59;
  assign t_r35_c58_7 = t_r35_c58_2 + t_r35_c58_3;
  assign t_r35_c58_8 = t_r35_c58_4 + p_36_57;
  assign t_r35_c58_9 = t_r35_c58_5 + t_r35_c58_6;
  assign t_r35_c58_10 = t_r35_c58_7 + t_r35_c58_8;
  assign t_r35_c58_11 = t_r35_c58_9 + t_r35_c58_10;
  assign t_r35_c58_12 = t_r35_c58_11 + p_36_59;
  assign out_35_58 = t_r35_c58_12 >> 4;

  assign t_r35_c59_0 = p_34_59 << 1;
  assign t_r35_c59_1 = p_35_58 << 1;
  assign t_r35_c59_2 = p_35_59 << 2;
  assign t_r35_c59_3 = p_35_60 << 1;
  assign t_r35_c59_4 = p_36_59 << 1;
  assign t_r35_c59_5 = t_r35_c59_0 + p_34_58;
  assign t_r35_c59_6 = t_r35_c59_1 + p_34_60;
  assign t_r35_c59_7 = t_r35_c59_2 + t_r35_c59_3;
  assign t_r35_c59_8 = t_r35_c59_4 + p_36_58;
  assign t_r35_c59_9 = t_r35_c59_5 + t_r35_c59_6;
  assign t_r35_c59_10 = t_r35_c59_7 + t_r35_c59_8;
  assign t_r35_c59_11 = t_r35_c59_9 + t_r35_c59_10;
  assign t_r35_c59_12 = t_r35_c59_11 + p_36_60;
  assign out_35_59 = t_r35_c59_12 >> 4;

  assign t_r35_c60_0 = p_34_60 << 1;
  assign t_r35_c60_1 = p_35_59 << 1;
  assign t_r35_c60_2 = p_35_60 << 2;
  assign t_r35_c60_3 = p_35_61 << 1;
  assign t_r35_c60_4 = p_36_60 << 1;
  assign t_r35_c60_5 = t_r35_c60_0 + p_34_59;
  assign t_r35_c60_6 = t_r35_c60_1 + p_34_61;
  assign t_r35_c60_7 = t_r35_c60_2 + t_r35_c60_3;
  assign t_r35_c60_8 = t_r35_c60_4 + p_36_59;
  assign t_r35_c60_9 = t_r35_c60_5 + t_r35_c60_6;
  assign t_r35_c60_10 = t_r35_c60_7 + t_r35_c60_8;
  assign t_r35_c60_11 = t_r35_c60_9 + t_r35_c60_10;
  assign t_r35_c60_12 = t_r35_c60_11 + p_36_61;
  assign out_35_60 = t_r35_c60_12 >> 4;

  assign t_r35_c61_0 = p_34_61 << 1;
  assign t_r35_c61_1 = p_35_60 << 1;
  assign t_r35_c61_2 = p_35_61 << 2;
  assign t_r35_c61_3 = p_35_62 << 1;
  assign t_r35_c61_4 = p_36_61 << 1;
  assign t_r35_c61_5 = t_r35_c61_0 + p_34_60;
  assign t_r35_c61_6 = t_r35_c61_1 + p_34_62;
  assign t_r35_c61_7 = t_r35_c61_2 + t_r35_c61_3;
  assign t_r35_c61_8 = t_r35_c61_4 + p_36_60;
  assign t_r35_c61_9 = t_r35_c61_5 + t_r35_c61_6;
  assign t_r35_c61_10 = t_r35_c61_7 + t_r35_c61_8;
  assign t_r35_c61_11 = t_r35_c61_9 + t_r35_c61_10;
  assign t_r35_c61_12 = t_r35_c61_11 + p_36_62;
  assign out_35_61 = t_r35_c61_12 >> 4;

  assign t_r35_c62_0 = p_34_62 << 1;
  assign t_r35_c62_1 = p_35_61 << 1;
  assign t_r35_c62_2 = p_35_62 << 2;
  assign t_r35_c62_3 = p_35_63 << 1;
  assign t_r35_c62_4 = p_36_62 << 1;
  assign t_r35_c62_5 = t_r35_c62_0 + p_34_61;
  assign t_r35_c62_6 = t_r35_c62_1 + p_34_63;
  assign t_r35_c62_7 = t_r35_c62_2 + t_r35_c62_3;
  assign t_r35_c62_8 = t_r35_c62_4 + p_36_61;
  assign t_r35_c62_9 = t_r35_c62_5 + t_r35_c62_6;
  assign t_r35_c62_10 = t_r35_c62_7 + t_r35_c62_8;
  assign t_r35_c62_11 = t_r35_c62_9 + t_r35_c62_10;
  assign t_r35_c62_12 = t_r35_c62_11 + p_36_63;
  assign out_35_62 = t_r35_c62_12 >> 4;

  assign t_r35_c63_0 = p_34_63 << 1;
  assign t_r35_c63_1 = p_35_62 << 1;
  assign t_r35_c63_2 = p_35_63 << 2;
  assign t_r35_c63_3 = p_35_64 << 1;
  assign t_r35_c63_4 = p_36_63 << 1;
  assign t_r35_c63_5 = t_r35_c63_0 + p_34_62;
  assign t_r35_c63_6 = t_r35_c63_1 + p_34_64;
  assign t_r35_c63_7 = t_r35_c63_2 + t_r35_c63_3;
  assign t_r35_c63_8 = t_r35_c63_4 + p_36_62;
  assign t_r35_c63_9 = t_r35_c63_5 + t_r35_c63_6;
  assign t_r35_c63_10 = t_r35_c63_7 + t_r35_c63_8;
  assign t_r35_c63_11 = t_r35_c63_9 + t_r35_c63_10;
  assign t_r35_c63_12 = t_r35_c63_11 + p_36_64;
  assign out_35_63 = t_r35_c63_12 >> 4;

  assign t_r35_c64_0 = p_34_64 << 1;
  assign t_r35_c64_1 = p_35_63 << 1;
  assign t_r35_c64_2 = p_35_64 << 2;
  assign t_r35_c64_3 = p_35_65 << 1;
  assign t_r35_c64_4 = p_36_64 << 1;
  assign t_r35_c64_5 = t_r35_c64_0 + p_34_63;
  assign t_r35_c64_6 = t_r35_c64_1 + p_34_65;
  assign t_r35_c64_7 = t_r35_c64_2 + t_r35_c64_3;
  assign t_r35_c64_8 = t_r35_c64_4 + p_36_63;
  assign t_r35_c64_9 = t_r35_c64_5 + t_r35_c64_6;
  assign t_r35_c64_10 = t_r35_c64_7 + t_r35_c64_8;
  assign t_r35_c64_11 = t_r35_c64_9 + t_r35_c64_10;
  assign t_r35_c64_12 = t_r35_c64_11 + p_36_65;
  assign out_35_64 = t_r35_c64_12 >> 4;

  assign t_r36_c1_0 = p_35_1 << 1;
  assign t_r36_c1_1 = p_36_0 << 1;
  assign t_r36_c1_2 = p_36_1 << 2;
  assign t_r36_c1_3 = p_36_2 << 1;
  assign t_r36_c1_4 = p_37_1 << 1;
  assign t_r36_c1_5 = t_r36_c1_0 + p_35_0;
  assign t_r36_c1_6 = t_r36_c1_1 + p_35_2;
  assign t_r36_c1_7 = t_r36_c1_2 + t_r36_c1_3;
  assign t_r36_c1_8 = t_r36_c1_4 + p_37_0;
  assign t_r36_c1_9 = t_r36_c1_5 + t_r36_c1_6;
  assign t_r36_c1_10 = t_r36_c1_7 + t_r36_c1_8;
  assign t_r36_c1_11 = t_r36_c1_9 + t_r36_c1_10;
  assign t_r36_c1_12 = t_r36_c1_11 + p_37_2;
  assign out_36_1 = t_r36_c1_12 >> 4;

  assign t_r36_c2_0 = p_35_2 << 1;
  assign t_r36_c2_1 = p_36_1 << 1;
  assign t_r36_c2_2 = p_36_2 << 2;
  assign t_r36_c2_3 = p_36_3 << 1;
  assign t_r36_c2_4 = p_37_2 << 1;
  assign t_r36_c2_5 = t_r36_c2_0 + p_35_1;
  assign t_r36_c2_6 = t_r36_c2_1 + p_35_3;
  assign t_r36_c2_7 = t_r36_c2_2 + t_r36_c2_3;
  assign t_r36_c2_8 = t_r36_c2_4 + p_37_1;
  assign t_r36_c2_9 = t_r36_c2_5 + t_r36_c2_6;
  assign t_r36_c2_10 = t_r36_c2_7 + t_r36_c2_8;
  assign t_r36_c2_11 = t_r36_c2_9 + t_r36_c2_10;
  assign t_r36_c2_12 = t_r36_c2_11 + p_37_3;
  assign out_36_2 = t_r36_c2_12 >> 4;

  assign t_r36_c3_0 = p_35_3 << 1;
  assign t_r36_c3_1 = p_36_2 << 1;
  assign t_r36_c3_2 = p_36_3 << 2;
  assign t_r36_c3_3 = p_36_4 << 1;
  assign t_r36_c3_4 = p_37_3 << 1;
  assign t_r36_c3_5 = t_r36_c3_0 + p_35_2;
  assign t_r36_c3_6 = t_r36_c3_1 + p_35_4;
  assign t_r36_c3_7 = t_r36_c3_2 + t_r36_c3_3;
  assign t_r36_c3_8 = t_r36_c3_4 + p_37_2;
  assign t_r36_c3_9 = t_r36_c3_5 + t_r36_c3_6;
  assign t_r36_c3_10 = t_r36_c3_7 + t_r36_c3_8;
  assign t_r36_c3_11 = t_r36_c3_9 + t_r36_c3_10;
  assign t_r36_c3_12 = t_r36_c3_11 + p_37_4;
  assign out_36_3 = t_r36_c3_12 >> 4;

  assign t_r36_c4_0 = p_35_4 << 1;
  assign t_r36_c4_1 = p_36_3 << 1;
  assign t_r36_c4_2 = p_36_4 << 2;
  assign t_r36_c4_3 = p_36_5 << 1;
  assign t_r36_c4_4 = p_37_4 << 1;
  assign t_r36_c4_5 = t_r36_c4_0 + p_35_3;
  assign t_r36_c4_6 = t_r36_c4_1 + p_35_5;
  assign t_r36_c4_7 = t_r36_c4_2 + t_r36_c4_3;
  assign t_r36_c4_8 = t_r36_c4_4 + p_37_3;
  assign t_r36_c4_9 = t_r36_c4_5 + t_r36_c4_6;
  assign t_r36_c4_10 = t_r36_c4_7 + t_r36_c4_8;
  assign t_r36_c4_11 = t_r36_c4_9 + t_r36_c4_10;
  assign t_r36_c4_12 = t_r36_c4_11 + p_37_5;
  assign out_36_4 = t_r36_c4_12 >> 4;

  assign t_r36_c5_0 = p_35_5 << 1;
  assign t_r36_c5_1 = p_36_4 << 1;
  assign t_r36_c5_2 = p_36_5 << 2;
  assign t_r36_c5_3 = p_36_6 << 1;
  assign t_r36_c5_4 = p_37_5 << 1;
  assign t_r36_c5_5 = t_r36_c5_0 + p_35_4;
  assign t_r36_c5_6 = t_r36_c5_1 + p_35_6;
  assign t_r36_c5_7 = t_r36_c5_2 + t_r36_c5_3;
  assign t_r36_c5_8 = t_r36_c5_4 + p_37_4;
  assign t_r36_c5_9 = t_r36_c5_5 + t_r36_c5_6;
  assign t_r36_c5_10 = t_r36_c5_7 + t_r36_c5_8;
  assign t_r36_c5_11 = t_r36_c5_9 + t_r36_c5_10;
  assign t_r36_c5_12 = t_r36_c5_11 + p_37_6;
  assign out_36_5 = t_r36_c5_12 >> 4;

  assign t_r36_c6_0 = p_35_6 << 1;
  assign t_r36_c6_1 = p_36_5 << 1;
  assign t_r36_c6_2 = p_36_6 << 2;
  assign t_r36_c6_3 = p_36_7 << 1;
  assign t_r36_c6_4 = p_37_6 << 1;
  assign t_r36_c6_5 = t_r36_c6_0 + p_35_5;
  assign t_r36_c6_6 = t_r36_c6_1 + p_35_7;
  assign t_r36_c6_7 = t_r36_c6_2 + t_r36_c6_3;
  assign t_r36_c6_8 = t_r36_c6_4 + p_37_5;
  assign t_r36_c6_9 = t_r36_c6_5 + t_r36_c6_6;
  assign t_r36_c6_10 = t_r36_c6_7 + t_r36_c6_8;
  assign t_r36_c6_11 = t_r36_c6_9 + t_r36_c6_10;
  assign t_r36_c6_12 = t_r36_c6_11 + p_37_7;
  assign out_36_6 = t_r36_c6_12 >> 4;

  assign t_r36_c7_0 = p_35_7 << 1;
  assign t_r36_c7_1 = p_36_6 << 1;
  assign t_r36_c7_2 = p_36_7 << 2;
  assign t_r36_c7_3 = p_36_8 << 1;
  assign t_r36_c7_4 = p_37_7 << 1;
  assign t_r36_c7_5 = t_r36_c7_0 + p_35_6;
  assign t_r36_c7_6 = t_r36_c7_1 + p_35_8;
  assign t_r36_c7_7 = t_r36_c7_2 + t_r36_c7_3;
  assign t_r36_c7_8 = t_r36_c7_4 + p_37_6;
  assign t_r36_c7_9 = t_r36_c7_5 + t_r36_c7_6;
  assign t_r36_c7_10 = t_r36_c7_7 + t_r36_c7_8;
  assign t_r36_c7_11 = t_r36_c7_9 + t_r36_c7_10;
  assign t_r36_c7_12 = t_r36_c7_11 + p_37_8;
  assign out_36_7 = t_r36_c7_12 >> 4;

  assign t_r36_c8_0 = p_35_8 << 1;
  assign t_r36_c8_1 = p_36_7 << 1;
  assign t_r36_c8_2 = p_36_8 << 2;
  assign t_r36_c8_3 = p_36_9 << 1;
  assign t_r36_c8_4 = p_37_8 << 1;
  assign t_r36_c8_5 = t_r36_c8_0 + p_35_7;
  assign t_r36_c8_6 = t_r36_c8_1 + p_35_9;
  assign t_r36_c8_7 = t_r36_c8_2 + t_r36_c8_3;
  assign t_r36_c8_8 = t_r36_c8_4 + p_37_7;
  assign t_r36_c8_9 = t_r36_c8_5 + t_r36_c8_6;
  assign t_r36_c8_10 = t_r36_c8_7 + t_r36_c8_8;
  assign t_r36_c8_11 = t_r36_c8_9 + t_r36_c8_10;
  assign t_r36_c8_12 = t_r36_c8_11 + p_37_9;
  assign out_36_8 = t_r36_c8_12 >> 4;

  assign t_r36_c9_0 = p_35_9 << 1;
  assign t_r36_c9_1 = p_36_8 << 1;
  assign t_r36_c9_2 = p_36_9 << 2;
  assign t_r36_c9_3 = p_36_10 << 1;
  assign t_r36_c9_4 = p_37_9 << 1;
  assign t_r36_c9_5 = t_r36_c9_0 + p_35_8;
  assign t_r36_c9_6 = t_r36_c9_1 + p_35_10;
  assign t_r36_c9_7 = t_r36_c9_2 + t_r36_c9_3;
  assign t_r36_c9_8 = t_r36_c9_4 + p_37_8;
  assign t_r36_c9_9 = t_r36_c9_5 + t_r36_c9_6;
  assign t_r36_c9_10 = t_r36_c9_7 + t_r36_c9_8;
  assign t_r36_c9_11 = t_r36_c9_9 + t_r36_c9_10;
  assign t_r36_c9_12 = t_r36_c9_11 + p_37_10;
  assign out_36_9 = t_r36_c9_12 >> 4;

  assign t_r36_c10_0 = p_35_10 << 1;
  assign t_r36_c10_1 = p_36_9 << 1;
  assign t_r36_c10_2 = p_36_10 << 2;
  assign t_r36_c10_3 = p_36_11 << 1;
  assign t_r36_c10_4 = p_37_10 << 1;
  assign t_r36_c10_5 = t_r36_c10_0 + p_35_9;
  assign t_r36_c10_6 = t_r36_c10_1 + p_35_11;
  assign t_r36_c10_7 = t_r36_c10_2 + t_r36_c10_3;
  assign t_r36_c10_8 = t_r36_c10_4 + p_37_9;
  assign t_r36_c10_9 = t_r36_c10_5 + t_r36_c10_6;
  assign t_r36_c10_10 = t_r36_c10_7 + t_r36_c10_8;
  assign t_r36_c10_11 = t_r36_c10_9 + t_r36_c10_10;
  assign t_r36_c10_12 = t_r36_c10_11 + p_37_11;
  assign out_36_10 = t_r36_c10_12 >> 4;

  assign t_r36_c11_0 = p_35_11 << 1;
  assign t_r36_c11_1 = p_36_10 << 1;
  assign t_r36_c11_2 = p_36_11 << 2;
  assign t_r36_c11_3 = p_36_12 << 1;
  assign t_r36_c11_4 = p_37_11 << 1;
  assign t_r36_c11_5 = t_r36_c11_0 + p_35_10;
  assign t_r36_c11_6 = t_r36_c11_1 + p_35_12;
  assign t_r36_c11_7 = t_r36_c11_2 + t_r36_c11_3;
  assign t_r36_c11_8 = t_r36_c11_4 + p_37_10;
  assign t_r36_c11_9 = t_r36_c11_5 + t_r36_c11_6;
  assign t_r36_c11_10 = t_r36_c11_7 + t_r36_c11_8;
  assign t_r36_c11_11 = t_r36_c11_9 + t_r36_c11_10;
  assign t_r36_c11_12 = t_r36_c11_11 + p_37_12;
  assign out_36_11 = t_r36_c11_12 >> 4;

  assign t_r36_c12_0 = p_35_12 << 1;
  assign t_r36_c12_1 = p_36_11 << 1;
  assign t_r36_c12_2 = p_36_12 << 2;
  assign t_r36_c12_3 = p_36_13 << 1;
  assign t_r36_c12_4 = p_37_12 << 1;
  assign t_r36_c12_5 = t_r36_c12_0 + p_35_11;
  assign t_r36_c12_6 = t_r36_c12_1 + p_35_13;
  assign t_r36_c12_7 = t_r36_c12_2 + t_r36_c12_3;
  assign t_r36_c12_8 = t_r36_c12_4 + p_37_11;
  assign t_r36_c12_9 = t_r36_c12_5 + t_r36_c12_6;
  assign t_r36_c12_10 = t_r36_c12_7 + t_r36_c12_8;
  assign t_r36_c12_11 = t_r36_c12_9 + t_r36_c12_10;
  assign t_r36_c12_12 = t_r36_c12_11 + p_37_13;
  assign out_36_12 = t_r36_c12_12 >> 4;

  assign t_r36_c13_0 = p_35_13 << 1;
  assign t_r36_c13_1 = p_36_12 << 1;
  assign t_r36_c13_2 = p_36_13 << 2;
  assign t_r36_c13_3 = p_36_14 << 1;
  assign t_r36_c13_4 = p_37_13 << 1;
  assign t_r36_c13_5 = t_r36_c13_0 + p_35_12;
  assign t_r36_c13_6 = t_r36_c13_1 + p_35_14;
  assign t_r36_c13_7 = t_r36_c13_2 + t_r36_c13_3;
  assign t_r36_c13_8 = t_r36_c13_4 + p_37_12;
  assign t_r36_c13_9 = t_r36_c13_5 + t_r36_c13_6;
  assign t_r36_c13_10 = t_r36_c13_7 + t_r36_c13_8;
  assign t_r36_c13_11 = t_r36_c13_9 + t_r36_c13_10;
  assign t_r36_c13_12 = t_r36_c13_11 + p_37_14;
  assign out_36_13 = t_r36_c13_12 >> 4;

  assign t_r36_c14_0 = p_35_14 << 1;
  assign t_r36_c14_1 = p_36_13 << 1;
  assign t_r36_c14_2 = p_36_14 << 2;
  assign t_r36_c14_3 = p_36_15 << 1;
  assign t_r36_c14_4 = p_37_14 << 1;
  assign t_r36_c14_5 = t_r36_c14_0 + p_35_13;
  assign t_r36_c14_6 = t_r36_c14_1 + p_35_15;
  assign t_r36_c14_7 = t_r36_c14_2 + t_r36_c14_3;
  assign t_r36_c14_8 = t_r36_c14_4 + p_37_13;
  assign t_r36_c14_9 = t_r36_c14_5 + t_r36_c14_6;
  assign t_r36_c14_10 = t_r36_c14_7 + t_r36_c14_8;
  assign t_r36_c14_11 = t_r36_c14_9 + t_r36_c14_10;
  assign t_r36_c14_12 = t_r36_c14_11 + p_37_15;
  assign out_36_14 = t_r36_c14_12 >> 4;

  assign t_r36_c15_0 = p_35_15 << 1;
  assign t_r36_c15_1 = p_36_14 << 1;
  assign t_r36_c15_2 = p_36_15 << 2;
  assign t_r36_c15_3 = p_36_16 << 1;
  assign t_r36_c15_4 = p_37_15 << 1;
  assign t_r36_c15_5 = t_r36_c15_0 + p_35_14;
  assign t_r36_c15_6 = t_r36_c15_1 + p_35_16;
  assign t_r36_c15_7 = t_r36_c15_2 + t_r36_c15_3;
  assign t_r36_c15_8 = t_r36_c15_4 + p_37_14;
  assign t_r36_c15_9 = t_r36_c15_5 + t_r36_c15_6;
  assign t_r36_c15_10 = t_r36_c15_7 + t_r36_c15_8;
  assign t_r36_c15_11 = t_r36_c15_9 + t_r36_c15_10;
  assign t_r36_c15_12 = t_r36_c15_11 + p_37_16;
  assign out_36_15 = t_r36_c15_12 >> 4;

  assign t_r36_c16_0 = p_35_16 << 1;
  assign t_r36_c16_1 = p_36_15 << 1;
  assign t_r36_c16_2 = p_36_16 << 2;
  assign t_r36_c16_3 = p_36_17 << 1;
  assign t_r36_c16_4 = p_37_16 << 1;
  assign t_r36_c16_5 = t_r36_c16_0 + p_35_15;
  assign t_r36_c16_6 = t_r36_c16_1 + p_35_17;
  assign t_r36_c16_7 = t_r36_c16_2 + t_r36_c16_3;
  assign t_r36_c16_8 = t_r36_c16_4 + p_37_15;
  assign t_r36_c16_9 = t_r36_c16_5 + t_r36_c16_6;
  assign t_r36_c16_10 = t_r36_c16_7 + t_r36_c16_8;
  assign t_r36_c16_11 = t_r36_c16_9 + t_r36_c16_10;
  assign t_r36_c16_12 = t_r36_c16_11 + p_37_17;
  assign out_36_16 = t_r36_c16_12 >> 4;

  assign t_r36_c17_0 = p_35_17 << 1;
  assign t_r36_c17_1 = p_36_16 << 1;
  assign t_r36_c17_2 = p_36_17 << 2;
  assign t_r36_c17_3 = p_36_18 << 1;
  assign t_r36_c17_4 = p_37_17 << 1;
  assign t_r36_c17_5 = t_r36_c17_0 + p_35_16;
  assign t_r36_c17_6 = t_r36_c17_1 + p_35_18;
  assign t_r36_c17_7 = t_r36_c17_2 + t_r36_c17_3;
  assign t_r36_c17_8 = t_r36_c17_4 + p_37_16;
  assign t_r36_c17_9 = t_r36_c17_5 + t_r36_c17_6;
  assign t_r36_c17_10 = t_r36_c17_7 + t_r36_c17_8;
  assign t_r36_c17_11 = t_r36_c17_9 + t_r36_c17_10;
  assign t_r36_c17_12 = t_r36_c17_11 + p_37_18;
  assign out_36_17 = t_r36_c17_12 >> 4;

  assign t_r36_c18_0 = p_35_18 << 1;
  assign t_r36_c18_1 = p_36_17 << 1;
  assign t_r36_c18_2 = p_36_18 << 2;
  assign t_r36_c18_3 = p_36_19 << 1;
  assign t_r36_c18_4 = p_37_18 << 1;
  assign t_r36_c18_5 = t_r36_c18_0 + p_35_17;
  assign t_r36_c18_6 = t_r36_c18_1 + p_35_19;
  assign t_r36_c18_7 = t_r36_c18_2 + t_r36_c18_3;
  assign t_r36_c18_8 = t_r36_c18_4 + p_37_17;
  assign t_r36_c18_9 = t_r36_c18_5 + t_r36_c18_6;
  assign t_r36_c18_10 = t_r36_c18_7 + t_r36_c18_8;
  assign t_r36_c18_11 = t_r36_c18_9 + t_r36_c18_10;
  assign t_r36_c18_12 = t_r36_c18_11 + p_37_19;
  assign out_36_18 = t_r36_c18_12 >> 4;

  assign t_r36_c19_0 = p_35_19 << 1;
  assign t_r36_c19_1 = p_36_18 << 1;
  assign t_r36_c19_2 = p_36_19 << 2;
  assign t_r36_c19_3 = p_36_20 << 1;
  assign t_r36_c19_4 = p_37_19 << 1;
  assign t_r36_c19_5 = t_r36_c19_0 + p_35_18;
  assign t_r36_c19_6 = t_r36_c19_1 + p_35_20;
  assign t_r36_c19_7 = t_r36_c19_2 + t_r36_c19_3;
  assign t_r36_c19_8 = t_r36_c19_4 + p_37_18;
  assign t_r36_c19_9 = t_r36_c19_5 + t_r36_c19_6;
  assign t_r36_c19_10 = t_r36_c19_7 + t_r36_c19_8;
  assign t_r36_c19_11 = t_r36_c19_9 + t_r36_c19_10;
  assign t_r36_c19_12 = t_r36_c19_11 + p_37_20;
  assign out_36_19 = t_r36_c19_12 >> 4;

  assign t_r36_c20_0 = p_35_20 << 1;
  assign t_r36_c20_1 = p_36_19 << 1;
  assign t_r36_c20_2 = p_36_20 << 2;
  assign t_r36_c20_3 = p_36_21 << 1;
  assign t_r36_c20_4 = p_37_20 << 1;
  assign t_r36_c20_5 = t_r36_c20_0 + p_35_19;
  assign t_r36_c20_6 = t_r36_c20_1 + p_35_21;
  assign t_r36_c20_7 = t_r36_c20_2 + t_r36_c20_3;
  assign t_r36_c20_8 = t_r36_c20_4 + p_37_19;
  assign t_r36_c20_9 = t_r36_c20_5 + t_r36_c20_6;
  assign t_r36_c20_10 = t_r36_c20_7 + t_r36_c20_8;
  assign t_r36_c20_11 = t_r36_c20_9 + t_r36_c20_10;
  assign t_r36_c20_12 = t_r36_c20_11 + p_37_21;
  assign out_36_20 = t_r36_c20_12 >> 4;

  assign t_r36_c21_0 = p_35_21 << 1;
  assign t_r36_c21_1 = p_36_20 << 1;
  assign t_r36_c21_2 = p_36_21 << 2;
  assign t_r36_c21_3 = p_36_22 << 1;
  assign t_r36_c21_4 = p_37_21 << 1;
  assign t_r36_c21_5 = t_r36_c21_0 + p_35_20;
  assign t_r36_c21_6 = t_r36_c21_1 + p_35_22;
  assign t_r36_c21_7 = t_r36_c21_2 + t_r36_c21_3;
  assign t_r36_c21_8 = t_r36_c21_4 + p_37_20;
  assign t_r36_c21_9 = t_r36_c21_5 + t_r36_c21_6;
  assign t_r36_c21_10 = t_r36_c21_7 + t_r36_c21_8;
  assign t_r36_c21_11 = t_r36_c21_9 + t_r36_c21_10;
  assign t_r36_c21_12 = t_r36_c21_11 + p_37_22;
  assign out_36_21 = t_r36_c21_12 >> 4;

  assign t_r36_c22_0 = p_35_22 << 1;
  assign t_r36_c22_1 = p_36_21 << 1;
  assign t_r36_c22_2 = p_36_22 << 2;
  assign t_r36_c22_3 = p_36_23 << 1;
  assign t_r36_c22_4 = p_37_22 << 1;
  assign t_r36_c22_5 = t_r36_c22_0 + p_35_21;
  assign t_r36_c22_6 = t_r36_c22_1 + p_35_23;
  assign t_r36_c22_7 = t_r36_c22_2 + t_r36_c22_3;
  assign t_r36_c22_8 = t_r36_c22_4 + p_37_21;
  assign t_r36_c22_9 = t_r36_c22_5 + t_r36_c22_6;
  assign t_r36_c22_10 = t_r36_c22_7 + t_r36_c22_8;
  assign t_r36_c22_11 = t_r36_c22_9 + t_r36_c22_10;
  assign t_r36_c22_12 = t_r36_c22_11 + p_37_23;
  assign out_36_22 = t_r36_c22_12 >> 4;

  assign t_r36_c23_0 = p_35_23 << 1;
  assign t_r36_c23_1 = p_36_22 << 1;
  assign t_r36_c23_2 = p_36_23 << 2;
  assign t_r36_c23_3 = p_36_24 << 1;
  assign t_r36_c23_4 = p_37_23 << 1;
  assign t_r36_c23_5 = t_r36_c23_0 + p_35_22;
  assign t_r36_c23_6 = t_r36_c23_1 + p_35_24;
  assign t_r36_c23_7 = t_r36_c23_2 + t_r36_c23_3;
  assign t_r36_c23_8 = t_r36_c23_4 + p_37_22;
  assign t_r36_c23_9 = t_r36_c23_5 + t_r36_c23_6;
  assign t_r36_c23_10 = t_r36_c23_7 + t_r36_c23_8;
  assign t_r36_c23_11 = t_r36_c23_9 + t_r36_c23_10;
  assign t_r36_c23_12 = t_r36_c23_11 + p_37_24;
  assign out_36_23 = t_r36_c23_12 >> 4;

  assign t_r36_c24_0 = p_35_24 << 1;
  assign t_r36_c24_1 = p_36_23 << 1;
  assign t_r36_c24_2 = p_36_24 << 2;
  assign t_r36_c24_3 = p_36_25 << 1;
  assign t_r36_c24_4 = p_37_24 << 1;
  assign t_r36_c24_5 = t_r36_c24_0 + p_35_23;
  assign t_r36_c24_6 = t_r36_c24_1 + p_35_25;
  assign t_r36_c24_7 = t_r36_c24_2 + t_r36_c24_3;
  assign t_r36_c24_8 = t_r36_c24_4 + p_37_23;
  assign t_r36_c24_9 = t_r36_c24_5 + t_r36_c24_6;
  assign t_r36_c24_10 = t_r36_c24_7 + t_r36_c24_8;
  assign t_r36_c24_11 = t_r36_c24_9 + t_r36_c24_10;
  assign t_r36_c24_12 = t_r36_c24_11 + p_37_25;
  assign out_36_24 = t_r36_c24_12 >> 4;

  assign t_r36_c25_0 = p_35_25 << 1;
  assign t_r36_c25_1 = p_36_24 << 1;
  assign t_r36_c25_2 = p_36_25 << 2;
  assign t_r36_c25_3 = p_36_26 << 1;
  assign t_r36_c25_4 = p_37_25 << 1;
  assign t_r36_c25_5 = t_r36_c25_0 + p_35_24;
  assign t_r36_c25_6 = t_r36_c25_1 + p_35_26;
  assign t_r36_c25_7 = t_r36_c25_2 + t_r36_c25_3;
  assign t_r36_c25_8 = t_r36_c25_4 + p_37_24;
  assign t_r36_c25_9 = t_r36_c25_5 + t_r36_c25_6;
  assign t_r36_c25_10 = t_r36_c25_7 + t_r36_c25_8;
  assign t_r36_c25_11 = t_r36_c25_9 + t_r36_c25_10;
  assign t_r36_c25_12 = t_r36_c25_11 + p_37_26;
  assign out_36_25 = t_r36_c25_12 >> 4;

  assign t_r36_c26_0 = p_35_26 << 1;
  assign t_r36_c26_1 = p_36_25 << 1;
  assign t_r36_c26_2 = p_36_26 << 2;
  assign t_r36_c26_3 = p_36_27 << 1;
  assign t_r36_c26_4 = p_37_26 << 1;
  assign t_r36_c26_5 = t_r36_c26_0 + p_35_25;
  assign t_r36_c26_6 = t_r36_c26_1 + p_35_27;
  assign t_r36_c26_7 = t_r36_c26_2 + t_r36_c26_3;
  assign t_r36_c26_8 = t_r36_c26_4 + p_37_25;
  assign t_r36_c26_9 = t_r36_c26_5 + t_r36_c26_6;
  assign t_r36_c26_10 = t_r36_c26_7 + t_r36_c26_8;
  assign t_r36_c26_11 = t_r36_c26_9 + t_r36_c26_10;
  assign t_r36_c26_12 = t_r36_c26_11 + p_37_27;
  assign out_36_26 = t_r36_c26_12 >> 4;

  assign t_r36_c27_0 = p_35_27 << 1;
  assign t_r36_c27_1 = p_36_26 << 1;
  assign t_r36_c27_2 = p_36_27 << 2;
  assign t_r36_c27_3 = p_36_28 << 1;
  assign t_r36_c27_4 = p_37_27 << 1;
  assign t_r36_c27_5 = t_r36_c27_0 + p_35_26;
  assign t_r36_c27_6 = t_r36_c27_1 + p_35_28;
  assign t_r36_c27_7 = t_r36_c27_2 + t_r36_c27_3;
  assign t_r36_c27_8 = t_r36_c27_4 + p_37_26;
  assign t_r36_c27_9 = t_r36_c27_5 + t_r36_c27_6;
  assign t_r36_c27_10 = t_r36_c27_7 + t_r36_c27_8;
  assign t_r36_c27_11 = t_r36_c27_9 + t_r36_c27_10;
  assign t_r36_c27_12 = t_r36_c27_11 + p_37_28;
  assign out_36_27 = t_r36_c27_12 >> 4;

  assign t_r36_c28_0 = p_35_28 << 1;
  assign t_r36_c28_1 = p_36_27 << 1;
  assign t_r36_c28_2 = p_36_28 << 2;
  assign t_r36_c28_3 = p_36_29 << 1;
  assign t_r36_c28_4 = p_37_28 << 1;
  assign t_r36_c28_5 = t_r36_c28_0 + p_35_27;
  assign t_r36_c28_6 = t_r36_c28_1 + p_35_29;
  assign t_r36_c28_7 = t_r36_c28_2 + t_r36_c28_3;
  assign t_r36_c28_8 = t_r36_c28_4 + p_37_27;
  assign t_r36_c28_9 = t_r36_c28_5 + t_r36_c28_6;
  assign t_r36_c28_10 = t_r36_c28_7 + t_r36_c28_8;
  assign t_r36_c28_11 = t_r36_c28_9 + t_r36_c28_10;
  assign t_r36_c28_12 = t_r36_c28_11 + p_37_29;
  assign out_36_28 = t_r36_c28_12 >> 4;

  assign t_r36_c29_0 = p_35_29 << 1;
  assign t_r36_c29_1 = p_36_28 << 1;
  assign t_r36_c29_2 = p_36_29 << 2;
  assign t_r36_c29_3 = p_36_30 << 1;
  assign t_r36_c29_4 = p_37_29 << 1;
  assign t_r36_c29_5 = t_r36_c29_0 + p_35_28;
  assign t_r36_c29_6 = t_r36_c29_1 + p_35_30;
  assign t_r36_c29_7 = t_r36_c29_2 + t_r36_c29_3;
  assign t_r36_c29_8 = t_r36_c29_4 + p_37_28;
  assign t_r36_c29_9 = t_r36_c29_5 + t_r36_c29_6;
  assign t_r36_c29_10 = t_r36_c29_7 + t_r36_c29_8;
  assign t_r36_c29_11 = t_r36_c29_9 + t_r36_c29_10;
  assign t_r36_c29_12 = t_r36_c29_11 + p_37_30;
  assign out_36_29 = t_r36_c29_12 >> 4;

  assign t_r36_c30_0 = p_35_30 << 1;
  assign t_r36_c30_1 = p_36_29 << 1;
  assign t_r36_c30_2 = p_36_30 << 2;
  assign t_r36_c30_3 = p_36_31 << 1;
  assign t_r36_c30_4 = p_37_30 << 1;
  assign t_r36_c30_5 = t_r36_c30_0 + p_35_29;
  assign t_r36_c30_6 = t_r36_c30_1 + p_35_31;
  assign t_r36_c30_7 = t_r36_c30_2 + t_r36_c30_3;
  assign t_r36_c30_8 = t_r36_c30_4 + p_37_29;
  assign t_r36_c30_9 = t_r36_c30_5 + t_r36_c30_6;
  assign t_r36_c30_10 = t_r36_c30_7 + t_r36_c30_8;
  assign t_r36_c30_11 = t_r36_c30_9 + t_r36_c30_10;
  assign t_r36_c30_12 = t_r36_c30_11 + p_37_31;
  assign out_36_30 = t_r36_c30_12 >> 4;

  assign t_r36_c31_0 = p_35_31 << 1;
  assign t_r36_c31_1 = p_36_30 << 1;
  assign t_r36_c31_2 = p_36_31 << 2;
  assign t_r36_c31_3 = p_36_32 << 1;
  assign t_r36_c31_4 = p_37_31 << 1;
  assign t_r36_c31_5 = t_r36_c31_0 + p_35_30;
  assign t_r36_c31_6 = t_r36_c31_1 + p_35_32;
  assign t_r36_c31_7 = t_r36_c31_2 + t_r36_c31_3;
  assign t_r36_c31_8 = t_r36_c31_4 + p_37_30;
  assign t_r36_c31_9 = t_r36_c31_5 + t_r36_c31_6;
  assign t_r36_c31_10 = t_r36_c31_7 + t_r36_c31_8;
  assign t_r36_c31_11 = t_r36_c31_9 + t_r36_c31_10;
  assign t_r36_c31_12 = t_r36_c31_11 + p_37_32;
  assign out_36_31 = t_r36_c31_12 >> 4;

  assign t_r36_c32_0 = p_35_32 << 1;
  assign t_r36_c32_1 = p_36_31 << 1;
  assign t_r36_c32_2 = p_36_32 << 2;
  assign t_r36_c32_3 = p_36_33 << 1;
  assign t_r36_c32_4 = p_37_32 << 1;
  assign t_r36_c32_5 = t_r36_c32_0 + p_35_31;
  assign t_r36_c32_6 = t_r36_c32_1 + p_35_33;
  assign t_r36_c32_7 = t_r36_c32_2 + t_r36_c32_3;
  assign t_r36_c32_8 = t_r36_c32_4 + p_37_31;
  assign t_r36_c32_9 = t_r36_c32_5 + t_r36_c32_6;
  assign t_r36_c32_10 = t_r36_c32_7 + t_r36_c32_8;
  assign t_r36_c32_11 = t_r36_c32_9 + t_r36_c32_10;
  assign t_r36_c32_12 = t_r36_c32_11 + p_37_33;
  assign out_36_32 = t_r36_c32_12 >> 4;

  assign t_r36_c33_0 = p_35_33 << 1;
  assign t_r36_c33_1 = p_36_32 << 1;
  assign t_r36_c33_2 = p_36_33 << 2;
  assign t_r36_c33_3 = p_36_34 << 1;
  assign t_r36_c33_4 = p_37_33 << 1;
  assign t_r36_c33_5 = t_r36_c33_0 + p_35_32;
  assign t_r36_c33_6 = t_r36_c33_1 + p_35_34;
  assign t_r36_c33_7 = t_r36_c33_2 + t_r36_c33_3;
  assign t_r36_c33_8 = t_r36_c33_4 + p_37_32;
  assign t_r36_c33_9 = t_r36_c33_5 + t_r36_c33_6;
  assign t_r36_c33_10 = t_r36_c33_7 + t_r36_c33_8;
  assign t_r36_c33_11 = t_r36_c33_9 + t_r36_c33_10;
  assign t_r36_c33_12 = t_r36_c33_11 + p_37_34;
  assign out_36_33 = t_r36_c33_12 >> 4;

  assign t_r36_c34_0 = p_35_34 << 1;
  assign t_r36_c34_1 = p_36_33 << 1;
  assign t_r36_c34_2 = p_36_34 << 2;
  assign t_r36_c34_3 = p_36_35 << 1;
  assign t_r36_c34_4 = p_37_34 << 1;
  assign t_r36_c34_5 = t_r36_c34_0 + p_35_33;
  assign t_r36_c34_6 = t_r36_c34_1 + p_35_35;
  assign t_r36_c34_7 = t_r36_c34_2 + t_r36_c34_3;
  assign t_r36_c34_8 = t_r36_c34_4 + p_37_33;
  assign t_r36_c34_9 = t_r36_c34_5 + t_r36_c34_6;
  assign t_r36_c34_10 = t_r36_c34_7 + t_r36_c34_8;
  assign t_r36_c34_11 = t_r36_c34_9 + t_r36_c34_10;
  assign t_r36_c34_12 = t_r36_c34_11 + p_37_35;
  assign out_36_34 = t_r36_c34_12 >> 4;

  assign t_r36_c35_0 = p_35_35 << 1;
  assign t_r36_c35_1 = p_36_34 << 1;
  assign t_r36_c35_2 = p_36_35 << 2;
  assign t_r36_c35_3 = p_36_36 << 1;
  assign t_r36_c35_4 = p_37_35 << 1;
  assign t_r36_c35_5 = t_r36_c35_0 + p_35_34;
  assign t_r36_c35_6 = t_r36_c35_1 + p_35_36;
  assign t_r36_c35_7 = t_r36_c35_2 + t_r36_c35_3;
  assign t_r36_c35_8 = t_r36_c35_4 + p_37_34;
  assign t_r36_c35_9 = t_r36_c35_5 + t_r36_c35_6;
  assign t_r36_c35_10 = t_r36_c35_7 + t_r36_c35_8;
  assign t_r36_c35_11 = t_r36_c35_9 + t_r36_c35_10;
  assign t_r36_c35_12 = t_r36_c35_11 + p_37_36;
  assign out_36_35 = t_r36_c35_12 >> 4;

  assign t_r36_c36_0 = p_35_36 << 1;
  assign t_r36_c36_1 = p_36_35 << 1;
  assign t_r36_c36_2 = p_36_36 << 2;
  assign t_r36_c36_3 = p_36_37 << 1;
  assign t_r36_c36_4 = p_37_36 << 1;
  assign t_r36_c36_5 = t_r36_c36_0 + p_35_35;
  assign t_r36_c36_6 = t_r36_c36_1 + p_35_37;
  assign t_r36_c36_7 = t_r36_c36_2 + t_r36_c36_3;
  assign t_r36_c36_8 = t_r36_c36_4 + p_37_35;
  assign t_r36_c36_9 = t_r36_c36_5 + t_r36_c36_6;
  assign t_r36_c36_10 = t_r36_c36_7 + t_r36_c36_8;
  assign t_r36_c36_11 = t_r36_c36_9 + t_r36_c36_10;
  assign t_r36_c36_12 = t_r36_c36_11 + p_37_37;
  assign out_36_36 = t_r36_c36_12 >> 4;

  assign t_r36_c37_0 = p_35_37 << 1;
  assign t_r36_c37_1 = p_36_36 << 1;
  assign t_r36_c37_2 = p_36_37 << 2;
  assign t_r36_c37_3 = p_36_38 << 1;
  assign t_r36_c37_4 = p_37_37 << 1;
  assign t_r36_c37_5 = t_r36_c37_0 + p_35_36;
  assign t_r36_c37_6 = t_r36_c37_1 + p_35_38;
  assign t_r36_c37_7 = t_r36_c37_2 + t_r36_c37_3;
  assign t_r36_c37_8 = t_r36_c37_4 + p_37_36;
  assign t_r36_c37_9 = t_r36_c37_5 + t_r36_c37_6;
  assign t_r36_c37_10 = t_r36_c37_7 + t_r36_c37_8;
  assign t_r36_c37_11 = t_r36_c37_9 + t_r36_c37_10;
  assign t_r36_c37_12 = t_r36_c37_11 + p_37_38;
  assign out_36_37 = t_r36_c37_12 >> 4;

  assign t_r36_c38_0 = p_35_38 << 1;
  assign t_r36_c38_1 = p_36_37 << 1;
  assign t_r36_c38_2 = p_36_38 << 2;
  assign t_r36_c38_3 = p_36_39 << 1;
  assign t_r36_c38_4 = p_37_38 << 1;
  assign t_r36_c38_5 = t_r36_c38_0 + p_35_37;
  assign t_r36_c38_6 = t_r36_c38_1 + p_35_39;
  assign t_r36_c38_7 = t_r36_c38_2 + t_r36_c38_3;
  assign t_r36_c38_8 = t_r36_c38_4 + p_37_37;
  assign t_r36_c38_9 = t_r36_c38_5 + t_r36_c38_6;
  assign t_r36_c38_10 = t_r36_c38_7 + t_r36_c38_8;
  assign t_r36_c38_11 = t_r36_c38_9 + t_r36_c38_10;
  assign t_r36_c38_12 = t_r36_c38_11 + p_37_39;
  assign out_36_38 = t_r36_c38_12 >> 4;

  assign t_r36_c39_0 = p_35_39 << 1;
  assign t_r36_c39_1 = p_36_38 << 1;
  assign t_r36_c39_2 = p_36_39 << 2;
  assign t_r36_c39_3 = p_36_40 << 1;
  assign t_r36_c39_4 = p_37_39 << 1;
  assign t_r36_c39_5 = t_r36_c39_0 + p_35_38;
  assign t_r36_c39_6 = t_r36_c39_1 + p_35_40;
  assign t_r36_c39_7 = t_r36_c39_2 + t_r36_c39_3;
  assign t_r36_c39_8 = t_r36_c39_4 + p_37_38;
  assign t_r36_c39_9 = t_r36_c39_5 + t_r36_c39_6;
  assign t_r36_c39_10 = t_r36_c39_7 + t_r36_c39_8;
  assign t_r36_c39_11 = t_r36_c39_9 + t_r36_c39_10;
  assign t_r36_c39_12 = t_r36_c39_11 + p_37_40;
  assign out_36_39 = t_r36_c39_12 >> 4;

  assign t_r36_c40_0 = p_35_40 << 1;
  assign t_r36_c40_1 = p_36_39 << 1;
  assign t_r36_c40_2 = p_36_40 << 2;
  assign t_r36_c40_3 = p_36_41 << 1;
  assign t_r36_c40_4 = p_37_40 << 1;
  assign t_r36_c40_5 = t_r36_c40_0 + p_35_39;
  assign t_r36_c40_6 = t_r36_c40_1 + p_35_41;
  assign t_r36_c40_7 = t_r36_c40_2 + t_r36_c40_3;
  assign t_r36_c40_8 = t_r36_c40_4 + p_37_39;
  assign t_r36_c40_9 = t_r36_c40_5 + t_r36_c40_6;
  assign t_r36_c40_10 = t_r36_c40_7 + t_r36_c40_8;
  assign t_r36_c40_11 = t_r36_c40_9 + t_r36_c40_10;
  assign t_r36_c40_12 = t_r36_c40_11 + p_37_41;
  assign out_36_40 = t_r36_c40_12 >> 4;

  assign t_r36_c41_0 = p_35_41 << 1;
  assign t_r36_c41_1 = p_36_40 << 1;
  assign t_r36_c41_2 = p_36_41 << 2;
  assign t_r36_c41_3 = p_36_42 << 1;
  assign t_r36_c41_4 = p_37_41 << 1;
  assign t_r36_c41_5 = t_r36_c41_0 + p_35_40;
  assign t_r36_c41_6 = t_r36_c41_1 + p_35_42;
  assign t_r36_c41_7 = t_r36_c41_2 + t_r36_c41_3;
  assign t_r36_c41_8 = t_r36_c41_4 + p_37_40;
  assign t_r36_c41_9 = t_r36_c41_5 + t_r36_c41_6;
  assign t_r36_c41_10 = t_r36_c41_7 + t_r36_c41_8;
  assign t_r36_c41_11 = t_r36_c41_9 + t_r36_c41_10;
  assign t_r36_c41_12 = t_r36_c41_11 + p_37_42;
  assign out_36_41 = t_r36_c41_12 >> 4;

  assign t_r36_c42_0 = p_35_42 << 1;
  assign t_r36_c42_1 = p_36_41 << 1;
  assign t_r36_c42_2 = p_36_42 << 2;
  assign t_r36_c42_3 = p_36_43 << 1;
  assign t_r36_c42_4 = p_37_42 << 1;
  assign t_r36_c42_5 = t_r36_c42_0 + p_35_41;
  assign t_r36_c42_6 = t_r36_c42_1 + p_35_43;
  assign t_r36_c42_7 = t_r36_c42_2 + t_r36_c42_3;
  assign t_r36_c42_8 = t_r36_c42_4 + p_37_41;
  assign t_r36_c42_9 = t_r36_c42_5 + t_r36_c42_6;
  assign t_r36_c42_10 = t_r36_c42_7 + t_r36_c42_8;
  assign t_r36_c42_11 = t_r36_c42_9 + t_r36_c42_10;
  assign t_r36_c42_12 = t_r36_c42_11 + p_37_43;
  assign out_36_42 = t_r36_c42_12 >> 4;

  assign t_r36_c43_0 = p_35_43 << 1;
  assign t_r36_c43_1 = p_36_42 << 1;
  assign t_r36_c43_2 = p_36_43 << 2;
  assign t_r36_c43_3 = p_36_44 << 1;
  assign t_r36_c43_4 = p_37_43 << 1;
  assign t_r36_c43_5 = t_r36_c43_0 + p_35_42;
  assign t_r36_c43_6 = t_r36_c43_1 + p_35_44;
  assign t_r36_c43_7 = t_r36_c43_2 + t_r36_c43_3;
  assign t_r36_c43_8 = t_r36_c43_4 + p_37_42;
  assign t_r36_c43_9 = t_r36_c43_5 + t_r36_c43_6;
  assign t_r36_c43_10 = t_r36_c43_7 + t_r36_c43_8;
  assign t_r36_c43_11 = t_r36_c43_9 + t_r36_c43_10;
  assign t_r36_c43_12 = t_r36_c43_11 + p_37_44;
  assign out_36_43 = t_r36_c43_12 >> 4;

  assign t_r36_c44_0 = p_35_44 << 1;
  assign t_r36_c44_1 = p_36_43 << 1;
  assign t_r36_c44_2 = p_36_44 << 2;
  assign t_r36_c44_3 = p_36_45 << 1;
  assign t_r36_c44_4 = p_37_44 << 1;
  assign t_r36_c44_5 = t_r36_c44_0 + p_35_43;
  assign t_r36_c44_6 = t_r36_c44_1 + p_35_45;
  assign t_r36_c44_7 = t_r36_c44_2 + t_r36_c44_3;
  assign t_r36_c44_8 = t_r36_c44_4 + p_37_43;
  assign t_r36_c44_9 = t_r36_c44_5 + t_r36_c44_6;
  assign t_r36_c44_10 = t_r36_c44_7 + t_r36_c44_8;
  assign t_r36_c44_11 = t_r36_c44_9 + t_r36_c44_10;
  assign t_r36_c44_12 = t_r36_c44_11 + p_37_45;
  assign out_36_44 = t_r36_c44_12 >> 4;

  assign t_r36_c45_0 = p_35_45 << 1;
  assign t_r36_c45_1 = p_36_44 << 1;
  assign t_r36_c45_2 = p_36_45 << 2;
  assign t_r36_c45_3 = p_36_46 << 1;
  assign t_r36_c45_4 = p_37_45 << 1;
  assign t_r36_c45_5 = t_r36_c45_0 + p_35_44;
  assign t_r36_c45_6 = t_r36_c45_1 + p_35_46;
  assign t_r36_c45_7 = t_r36_c45_2 + t_r36_c45_3;
  assign t_r36_c45_8 = t_r36_c45_4 + p_37_44;
  assign t_r36_c45_9 = t_r36_c45_5 + t_r36_c45_6;
  assign t_r36_c45_10 = t_r36_c45_7 + t_r36_c45_8;
  assign t_r36_c45_11 = t_r36_c45_9 + t_r36_c45_10;
  assign t_r36_c45_12 = t_r36_c45_11 + p_37_46;
  assign out_36_45 = t_r36_c45_12 >> 4;

  assign t_r36_c46_0 = p_35_46 << 1;
  assign t_r36_c46_1 = p_36_45 << 1;
  assign t_r36_c46_2 = p_36_46 << 2;
  assign t_r36_c46_3 = p_36_47 << 1;
  assign t_r36_c46_4 = p_37_46 << 1;
  assign t_r36_c46_5 = t_r36_c46_0 + p_35_45;
  assign t_r36_c46_6 = t_r36_c46_1 + p_35_47;
  assign t_r36_c46_7 = t_r36_c46_2 + t_r36_c46_3;
  assign t_r36_c46_8 = t_r36_c46_4 + p_37_45;
  assign t_r36_c46_9 = t_r36_c46_5 + t_r36_c46_6;
  assign t_r36_c46_10 = t_r36_c46_7 + t_r36_c46_8;
  assign t_r36_c46_11 = t_r36_c46_9 + t_r36_c46_10;
  assign t_r36_c46_12 = t_r36_c46_11 + p_37_47;
  assign out_36_46 = t_r36_c46_12 >> 4;

  assign t_r36_c47_0 = p_35_47 << 1;
  assign t_r36_c47_1 = p_36_46 << 1;
  assign t_r36_c47_2 = p_36_47 << 2;
  assign t_r36_c47_3 = p_36_48 << 1;
  assign t_r36_c47_4 = p_37_47 << 1;
  assign t_r36_c47_5 = t_r36_c47_0 + p_35_46;
  assign t_r36_c47_6 = t_r36_c47_1 + p_35_48;
  assign t_r36_c47_7 = t_r36_c47_2 + t_r36_c47_3;
  assign t_r36_c47_8 = t_r36_c47_4 + p_37_46;
  assign t_r36_c47_9 = t_r36_c47_5 + t_r36_c47_6;
  assign t_r36_c47_10 = t_r36_c47_7 + t_r36_c47_8;
  assign t_r36_c47_11 = t_r36_c47_9 + t_r36_c47_10;
  assign t_r36_c47_12 = t_r36_c47_11 + p_37_48;
  assign out_36_47 = t_r36_c47_12 >> 4;

  assign t_r36_c48_0 = p_35_48 << 1;
  assign t_r36_c48_1 = p_36_47 << 1;
  assign t_r36_c48_2 = p_36_48 << 2;
  assign t_r36_c48_3 = p_36_49 << 1;
  assign t_r36_c48_4 = p_37_48 << 1;
  assign t_r36_c48_5 = t_r36_c48_0 + p_35_47;
  assign t_r36_c48_6 = t_r36_c48_1 + p_35_49;
  assign t_r36_c48_7 = t_r36_c48_2 + t_r36_c48_3;
  assign t_r36_c48_8 = t_r36_c48_4 + p_37_47;
  assign t_r36_c48_9 = t_r36_c48_5 + t_r36_c48_6;
  assign t_r36_c48_10 = t_r36_c48_7 + t_r36_c48_8;
  assign t_r36_c48_11 = t_r36_c48_9 + t_r36_c48_10;
  assign t_r36_c48_12 = t_r36_c48_11 + p_37_49;
  assign out_36_48 = t_r36_c48_12 >> 4;

  assign t_r36_c49_0 = p_35_49 << 1;
  assign t_r36_c49_1 = p_36_48 << 1;
  assign t_r36_c49_2 = p_36_49 << 2;
  assign t_r36_c49_3 = p_36_50 << 1;
  assign t_r36_c49_4 = p_37_49 << 1;
  assign t_r36_c49_5 = t_r36_c49_0 + p_35_48;
  assign t_r36_c49_6 = t_r36_c49_1 + p_35_50;
  assign t_r36_c49_7 = t_r36_c49_2 + t_r36_c49_3;
  assign t_r36_c49_8 = t_r36_c49_4 + p_37_48;
  assign t_r36_c49_9 = t_r36_c49_5 + t_r36_c49_6;
  assign t_r36_c49_10 = t_r36_c49_7 + t_r36_c49_8;
  assign t_r36_c49_11 = t_r36_c49_9 + t_r36_c49_10;
  assign t_r36_c49_12 = t_r36_c49_11 + p_37_50;
  assign out_36_49 = t_r36_c49_12 >> 4;

  assign t_r36_c50_0 = p_35_50 << 1;
  assign t_r36_c50_1 = p_36_49 << 1;
  assign t_r36_c50_2 = p_36_50 << 2;
  assign t_r36_c50_3 = p_36_51 << 1;
  assign t_r36_c50_4 = p_37_50 << 1;
  assign t_r36_c50_5 = t_r36_c50_0 + p_35_49;
  assign t_r36_c50_6 = t_r36_c50_1 + p_35_51;
  assign t_r36_c50_7 = t_r36_c50_2 + t_r36_c50_3;
  assign t_r36_c50_8 = t_r36_c50_4 + p_37_49;
  assign t_r36_c50_9 = t_r36_c50_5 + t_r36_c50_6;
  assign t_r36_c50_10 = t_r36_c50_7 + t_r36_c50_8;
  assign t_r36_c50_11 = t_r36_c50_9 + t_r36_c50_10;
  assign t_r36_c50_12 = t_r36_c50_11 + p_37_51;
  assign out_36_50 = t_r36_c50_12 >> 4;

  assign t_r36_c51_0 = p_35_51 << 1;
  assign t_r36_c51_1 = p_36_50 << 1;
  assign t_r36_c51_2 = p_36_51 << 2;
  assign t_r36_c51_3 = p_36_52 << 1;
  assign t_r36_c51_4 = p_37_51 << 1;
  assign t_r36_c51_5 = t_r36_c51_0 + p_35_50;
  assign t_r36_c51_6 = t_r36_c51_1 + p_35_52;
  assign t_r36_c51_7 = t_r36_c51_2 + t_r36_c51_3;
  assign t_r36_c51_8 = t_r36_c51_4 + p_37_50;
  assign t_r36_c51_9 = t_r36_c51_5 + t_r36_c51_6;
  assign t_r36_c51_10 = t_r36_c51_7 + t_r36_c51_8;
  assign t_r36_c51_11 = t_r36_c51_9 + t_r36_c51_10;
  assign t_r36_c51_12 = t_r36_c51_11 + p_37_52;
  assign out_36_51 = t_r36_c51_12 >> 4;

  assign t_r36_c52_0 = p_35_52 << 1;
  assign t_r36_c52_1 = p_36_51 << 1;
  assign t_r36_c52_2 = p_36_52 << 2;
  assign t_r36_c52_3 = p_36_53 << 1;
  assign t_r36_c52_4 = p_37_52 << 1;
  assign t_r36_c52_5 = t_r36_c52_0 + p_35_51;
  assign t_r36_c52_6 = t_r36_c52_1 + p_35_53;
  assign t_r36_c52_7 = t_r36_c52_2 + t_r36_c52_3;
  assign t_r36_c52_8 = t_r36_c52_4 + p_37_51;
  assign t_r36_c52_9 = t_r36_c52_5 + t_r36_c52_6;
  assign t_r36_c52_10 = t_r36_c52_7 + t_r36_c52_8;
  assign t_r36_c52_11 = t_r36_c52_9 + t_r36_c52_10;
  assign t_r36_c52_12 = t_r36_c52_11 + p_37_53;
  assign out_36_52 = t_r36_c52_12 >> 4;

  assign t_r36_c53_0 = p_35_53 << 1;
  assign t_r36_c53_1 = p_36_52 << 1;
  assign t_r36_c53_2 = p_36_53 << 2;
  assign t_r36_c53_3 = p_36_54 << 1;
  assign t_r36_c53_4 = p_37_53 << 1;
  assign t_r36_c53_5 = t_r36_c53_0 + p_35_52;
  assign t_r36_c53_6 = t_r36_c53_1 + p_35_54;
  assign t_r36_c53_7 = t_r36_c53_2 + t_r36_c53_3;
  assign t_r36_c53_8 = t_r36_c53_4 + p_37_52;
  assign t_r36_c53_9 = t_r36_c53_5 + t_r36_c53_6;
  assign t_r36_c53_10 = t_r36_c53_7 + t_r36_c53_8;
  assign t_r36_c53_11 = t_r36_c53_9 + t_r36_c53_10;
  assign t_r36_c53_12 = t_r36_c53_11 + p_37_54;
  assign out_36_53 = t_r36_c53_12 >> 4;

  assign t_r36_c54_0 = p_35_54 << 1;
  assign t_r36_c54_1 = p_36_53 << 1;
  assign t_r36_c54_2 = p_36_54 << 2;
  assign t_r36_c54_3 = p_36_55 << 1;
  assign t_r36_c54_4 = p_37_54 << 1;
  assign t_r36_c54_5 = t_r36_c54_0 + p_35_53;
  assign t_r36_c54_6 = t_r36_c54_1 + p_35_55;
  assign t_r36_c54_7 = t_r36_c54_2 + t_r36_c54_3;
  assign t_r36_c54_8 = t_r36_c54_4 + p_37_53;
  assign t_r36_c54_9 = t_r36_c54_5 + t_r36_c54_6;
  assign t_r36_c54_10 = t_r36_c54_7 + t_r36_c54_8;
  assign t_r36_c54_11 = t_r36_c54_9 + t_r36_c54_10;
  assign t_r36_c54_12 = t_r36_c54_11 + p_37_55;
  assign out_36_54 = t_r36_c54_12 >> 4;

  assign t_r36_c55_0 = p_35_55 << 1;
  assign t_r36_c55_1 = p_36_54 << 1;
  assign t_r36_c55_2 = p_36_55 << 2;
  assign t_r36_c55_3 = p_36_56 << 1;
  assign t_r36_c55_4 = p_37_55 << 1;
  assign t_r36_c55_5 = t_r36_c55_0 + p_35_54;
  assign t_r36_c55_6 = t_r36_c55_1 + p_35_56;
  assign t_r36_c55_7 = t_r36_c55_2 + t_r36_c55_3;
  assign t_r36_c55_8 = t_r36_c55_4 + p_37_54;
  assign t_r36_c55_9 = t_r36_c55_5 + t_r36_c55_6;
  assign t_r36_c55_10 = t_r36_c55_7 + t_r36_c55_8;
  assign t_r36_c55_11 = t_r36_c55_9 + t_r36_c55_10;
  assign t_r36_c55_12 = t_r36_c55_11 + p_37_56;
  assign out_36_55 = t_r36_c55_12 >> 4;

  assign t_r36_c56_0 = p_35_56 << 1;
  assign t_r36_c56_1 = p_36_55 << 1;
  assign t_r36_c56_2 = p_36_56 << 2;
  assign t_r36_c56_3 = p_36_57 << 1;
  assign t_r36_c56_4 = p_37_56 << 1;
  assign t_r36_c56_5 = t_r36_c56_0 + p_35_55;
  assign t_r36_c56_6 = t_r36_c56_1 + p_35_57;
  assign t_r36_c56_7 = t_r36_c56_2 + t_r36_c56_3;
  assign t_r36_c56_8 = t_r36_c56_4 + p_37_55;
  assign t_r36_c56_9 = t_r36_c56_5 + t_r36_c56_6;
  assign t_r36_c56_10 = t_r36_c56_7 + t_r36_c56_8;
  assign t_r36_c56_11 = t_r36_c56_9 + t_r36_c56_10;
  assign t_r36_c56_12 = t_r36_c56_11 + p_37_57;
  assign out_36_56 = t_r36_c56_12 >> 4;

  assign t_r36_c57_0 = p_35_57 << 1;
  assign t_r36_c57_1 = p_36_56 << 1;
  assign t_r36_c57_2 = p_36_57 << 2;
  assign t_r36_c57_3 = p_36_58 << 1;
  assign t_r36_c57_4 = p_37_57 << 1;
  assign t_r36_c57_5 = t_r36_c57_0 + p_35_56;
  assign t_r36_c57_6 = t_r36_c57_1 + p_35_58;
  assign t_r36_c57_7 = t_r36_c57_2 + t_r36_c57_3;
  assign t_r36_c57_8 = t_r36_c57_4 + p_37_56;
  assign t_r36_c57_9 = t_r36_c57_5 + t_r36_c57_6;
  assign t_r36_c57_10 = t_r36_c57_7 + t_r36_c57_8;
  assign t_r36_c57_11 = t_r36_c57_9 + t_r36_c57_10;
  assign t_r36_c57_12 = t_r36_c57_11 + p_37_58;
  assign out_36_57 = t_r36_c57_12 >> 4;

  assign t_r36_c58_0 = p_35_58 << 1;
  assign t_r36_c58_1 = p_36_57 << 1;
  assign t_r36_c58_2 = p_36_58 << 2;
  assign t_r36_c58_3 = p_36_59 << 1;
  assign t_r36_c58_4 = p_37_58 << 1;
  assign t_r36_c58_5 = t_r36_c58_0 + p_35_57;
  assign t_r36_c58_6 = t_r36_c58_1 + p_35_59;
  assign t_r36_c58_7 = t_r36_c58_2 + t_r36_c58_3;
  assign t_r36_c58_8 = t_r36_c58_4 + p_37_57;
  assign t_r36_c58_9 = t_r36_c58_5 + t_r36_c58_6;
  assign t_r36_c58_10 = t_r36_c58_7 + t_r36_c58_8;
  assign t_r36_c58_11 = t_r36_c58_9 + t_r36_c58_10;
  assign t_r36_c58_12 = t_r36_c58_11 + p_37_59;
  assign out_36_58 = t_r36_c58_12 >> 4;

  assign t_r36_c59_0 = p_35_59 << 1;
  assign t_r36_c59_1 = p_36_58 << 1;
  assign t_r36_c59_2 = p_36_59 << 2;
  assign t_r36_c59_3 = p_36_60 << 1;
  assign t_r36_c59_4 = p_37_59 << 1;
  assign t_r36_c59_5 = t_r36_c59_0 + p_35_58;
  assign t_r36_c59_6 = t_r36_c59_1 + p_35_60;
  assign t_r36_c59_7 = t_r36_c59_2 + t_r36_c59_3;
  assign t_r36_c59_8 = t_r36_c59_4 + p_37_58;
  assign t_r36_c59_9 = t_r36_c59_5 + t_r36_c59_6;
  assign t_r36_c59_10 = t_r36_c59_7 + t_r36_c59_8;
  assign t_r36_c59_11 = t_r36_c59_9 + t_r36_c59_10;
  assign t_r36_c59_12 = t_r36_c59_11 + p_37_60;
  assign out_36_59 = t_r36_c59_12 >> 4;

  assign t_r36_c60_0 = p_35_60 << 1;
  assign t_r36_c60_1 = p_36_59 << 1;
  assign t_r36_c60_2 = p_36_60 << 2;
  assign t_r36_c60_3 = p_36_61 << 1;
  assign t_r36_c60_4 = p_37_60 << 1;
  assign t_r36_c60_5 = t_r36_c60_0 + p_35_59;
  assign t_r36_c60_6 = t_r36_c60_1 + p_35_61;
  assign t_r36_c60_7 = t_r36_c60_2 + t_r36_c60_3;
  assign t_r36_c60_8 = t_r36_c60_4 + p_37_59;
  assign t_r36_c60_9 = t_r36_c60_5 + t_r36_c60_6;
  assign t_r36_c60_10 = t_r36_c60_7 + t_r36_c60_8;
  assign t_r36_c60_11 = t_r36_c60_9 + t_r36_c60_10;
  assign t_r36_c60_12 = t_r36_c60_11 + p_37_61;
  assign out_36_60 = t_r36_c60_12 >> 4;

  assign t_r36_c61_0 = p_35_61 << 1;
  assign t_r36_c61_1 = p_36_60 << 1;
  assign t_r36_c61_2 = p_36_61 << 2;
  assign t_r36_c61_3 = p_36_62 << 1;
  assign t_r36_c61_4 = p_37_61 << 1;
  assign t_r36_c61_5 = t_r36_c61_0 + p_35_60;
  assign t_r36_c61_6 = t_r36_c61_1 + p_35_62;
  assign t_r36_c61_7 = t_r36_c61_2 + t_r36_c61_3;
  assign t_r36_c61_8 = t_r36_c61_4 + p_37_60;
  assign t_r36_c61_9 = t_r36_c61_5 + t_r36_c61_6;
  assign t_r36_c61_10 = t_r36_c61_7 + t_r36_c61_8;
  assign t_r36_c61_11 = t_r36_c61_9 + t_r36_c61_10;
  assign t_r36_c61_12 = t_r36_c61_11 + p_37_62;
  assign out_36_61 = t_r36_c61_12 >> 4;

  assign t_r36_c62_0 = p_35_62 << 1;
  assign t_r36_c62_1 = p_36_61 << 1;
  assign t_r36_c62_2 = p_36_62 << 2;
  assign t_r36_c62_3 = p_36_63 << 1;
  assign t_r36_c62_4 = p_37_62 << 1;
  assign t_r36_c62_5 = t_r36_c62_0 + p_35_61;
  assign t_r36_c62_6 = t_r36_c62_1 + p_35_63;
  assign t_r36_c62_7 = t_r36_c62_2 + t_r36_c62_3;
  assign t_r36_c62_8 = t_r36_c62_4 + p_37_61;
  assign t_r36_c62_9 = t_r36_c62_5 + t_r36_c62_6;
  assign t_r36_c62_10 = t_r36_c62_7 + t_r36_c62_8;
  assign t_r36_c62_11 = t_r36_c62_9 + t_r36_c62_10;
  assign t_r36_c62_12 = t_r36_c62_11 + p_37_63;
  assign out_36_62 = t_r36_c62_12 >> 4;

  assign t_r36_c63_0 = p_35_63 << 1;
  assign t_r36_c63_1 = p_36_62 << 1;
  assign t_r36_c63_2 = p_36_63 << 2;
  assign t_r36_c63_3 = p_36_64 << 1;
  assign t_r36_c63_4 = p_37_63 << 1;
  assign t_r36_c63_5 = t_r36_c63_0 + p_35_62;
  assign t_r36_c63_6 = t_r36_c63_1 + p_35_64;
  assign t_r36_c63_7 = t_r36_c63_2 + t_r36_c63_3;
  assign t_r36_c63_8 = t_r36_c63_4 + p_37_62;
  assign t_r36_c63_9 = t_r36_c63_5 + t_r36_c63_6;
  assign t_r36_c63_10 = t_r36_c63_7 + t_r36_c63_8;
  assign t_r36_c63_11 = t_r36_c63_9 + t_r36_c63_10;
  assign t_r36_c63_12 = t_r36_c63_11 + p_37_64;
  assign out_36_63 = t_r36_c63_12 >> 4;

  assign t_r36_c64_0 = p_35_64 << 1;
  assign t_r36_c64_1 = p_36_63 << 1;
  assign t_r36_c64_2 = p_36_64 << 2;
  assign t_r36_c64_3 = p_36_65 << 1;
  assign t_r36_c64_4 = p_37_64 << 1;
  assign t_r36_c64_5 = t_r36_c64_0 + p_35_63;
  assign t_r36_c64_6 = t_r36_c64_1 + p_35_65;
  assign t_r36_c64_7 = t_r36_c64_2 + t_r36_c64_3;
  assign t_r36_c64_8 = t_r36_c64_4 + p_37_63;
  assign t_r36_c64_9 = t_r36_c64_5 + t_r36_c64_6;
  assign t_r36_c64_10 = t_r36_c64_7 + t_r36_c64_8;
  assign t_r36_c64_11 = t_r36_c64_9 + t_r36_c64_10;
  assign t_r36_c64_12 = t_r36_c64_11 + p_37_65;
  assign out_36_64 = t_r36_c64_12 >> 4;

  assign t_r37_c1_0 = p_36_1 << 1;
  assign t_r37_c1_1 = p_37_0 << 1;
  assign t_r37_c1_2 = p_37_1 << 2;
  assign t_r37_c1_3 = p_37_2 << 1;
  assign t_r37_c1_4 = p_38_1 << 1;
  assign t_r37_c1_5 = t_r37_c1_0 + p_36_0;
  assign t_r37_c1_6 = t_r37_c1_1 + p_36_2;
  assign t_r37_c1_7 = t_r37_c1_2 + t_r37_c1_3;
  assign t_r37_c1_8 = t_r37_c1_4 + p_38_0;
  assign t_r37_c1_9 = t_r37_c1_5 + t_r37_c1_6;
  assign t_r37_c1_10 = t_r37_c1_7 + t_r37_c1_8;
  assign t_r37_c1_11 = t_r37_c1_9 + t_r37_c1_10;
  assign t_r37_c1_12 = t_r37_c1_11 + p_38_2;
  assign out_37_1 = t_r37_c1_12 >> 4;

  assign t_r37_c2_0 = p_36_2 << 1;
  assign t_r37_c2_1 = p_37_1 << 1;
  assign t_r37_c2_2 = p_37_2 << 2;
  assign t_r37_c2_3 = p_37_3 << 1;
  assign t_r37_c2_4 = p_38_2 << 1;
  assign t_r37_c2_5 = t_r37_c2_0 + p_36_1;
  assign t_r37_c2_6 = t_r37_c2_1 + p_36_3;
  assign t_r37_c2_7 = t_r37_c2_2 + t_r37_c2_3;
  assign t_r37_c2_8 = t_r37_c2_4 + p_38_1;
  assign t_r37_c2_9 = t_r37_c2_5 + t_r37_c2_6;
  assign t_r37_c2_10 = t_r37_c2_7 + t_r37_c2_8;
  assign t_r37_c2_11 = t_r37_c2_9 + t_r37_c2_10;
  assign t_r37_c2_12 = t_r37_c2_11 + p_38_3;
  assign out_37_2 = t_r37_c2_12 >> 4;

  assign t_r37_c3_0 = p_36_3 << 1;
  assign t_r37_c3_1 = p_37_2 << 1;
  assign t_r37_c3_2 = p_37_3 << 2;
  assign t_r37_c3_3 = p_37_4 << 1;
  assign t_r37_c3_4 = p_38_3 << 1;
  assign t_r37_c3_5 = t_r37_c3_0 + p_36_2;
  assign t_r37_c3_6 = t_r37_c3_1 + p_36_4;
  assign t_r37_c3_7 = t_r37_c3_2 + t_r37_c3_3;
  assign t_r37_c3_8 = t_r37_c3_4 + p_38_2;
  assign t_r37_c3_9 = t_r37_c3_5 + t_r37_c3_6;
  assign t_r37_c3_10 = t_r37_c3_7 + t_r37_c3_8;
  assign t_r37_c3_11 = t_r37_c3_9 + t_r37_c3_10;
  assign t_r37_c3_12 = t_r37_c3_11 + p_38_4;
  assign out_37_3 = t_r37_c3_12 >> 4;

  assign t_r37_c4_0 = p_36_4 << 1;
  assign t_r37_c4_1 = p_37_3 << 1;
  assign t_r37_c4_2 = p_37_4 << 2;
  assign t_r37_c4_3 = p_37_5 << 1;
  assign t_r37_c4_4 = p_38_4 << 1;
  assign t_r37_c4_5 = t_r37_c4_0 + p_36_3;
  assign t_r37_c4_6 = t_r37_c4_1 + p_36_5;
  assign t_r37_c4_7 = t_r37_c4_2 + t_r37_c4_3;
  assign t_r37_c4_8 = t_r37_c4_4 + p_38_3;
  assign t_r37_c4_9 = t_r37_c4_5 + t_r37_c4_6;
  assign t_r37_c4_10 = t_r37_c4_7 + t_r37_c4_8;
  assign t_r37_c4_11 = t_r37_c4_9 + t_r37_c4_10;
  assign t_r37_c4_12 = t_r37_c4_11 + p_38_5;
  assign out_37_4 = t_r37_c4_12 >> 4;

  assign t_r37_c5_0 = p_36_5 << 1;
  assign t_r37_c5_1 = p_37_4 << 1;
  assign t_r37_c5_2 = p_37_5 << 2;
  assign t_r37_c5_3 = p_37_6 << 1;
  assign t_r37_c5_4 = p_38_5 << 1;
  assign t_r37_c5_5 = t_r37_c5_0 + p_36_4;
  assign t_r37_c5_6 = t_r37_c5_1 + p_36_6;
  assign t_r37_c5_7 = t_r37_c5_2 + t_r37_c5_3;
  assign t_r37_c5_8 = t_r37_c5_4 + p_38_4;
  assign t_r37_c5_9 = t_r37_c5_5 + t_r37_c5_6;
  assign t_r37_c5_10 = t_r37_c5_7 + t_r37_c5_8;
  assign t_r37_c5_11 = t_r37_c5_9 + t_r37_c5_10;
  assign t_r37_c5_12 = t_r37_c5_11 + p_38_6;
  assign out_37_5 = t_r37_c5_12 >> 4;

  assign t_r37_c6_0 = p_36_6 << 1;
  assign t_r37_c6_1 = p_37_5 << 1;
  assign t_r37_c6_2 = p_37_6 << 2;
  assign t_r37_c6_3 = p_37_7 << 1;
  assign t_r37_c6_4 = p_38_6 << 1;
  assign t_r37_c6_5 = t_r37_c6_0 + p_36_5;
  assign t_r37_c6_6 = t_r37_c6_1 + p_36_7;
  assign t_r37_c6_7 = t_r37_c6_2 + t_r37_c6_3;
  assign t_r37_c6_8 = t_r37_c6_4 + p_38_5;
  assign t_r37_c6_9 = t_r37_c6_5 + t_r37_c6_6;
  assign t_r37_c6_10 = t_r37_c6_7 + t_r37_c6_8;
  assign t_r37_c6_11 = t_r37_c6_9 + t_r37_c6_10;
  assign t_r37_c6_12 = t_r37_c6_11 + p_38_7;
  assign out_37_6 = t_r37_c6_12 >> 4;

  assign t_r37_c7_0 = p_36_7 << 1;
  assign t_r37_c7_1 = p_37_6 << 1;
  assign t_r37_c7_2 = p_37_7 << 2;
  assign t_r37_c7_3 = p_37_8 << 1;
  assign t_r37_c7_4 = p_38_7 << 1;
  assign t_r37_c7_5 = t_r37_c7_0 + p_36_6;
  assign t_r37_c7_6 = t_r37_c7_1 + p_36_8;
  assign t_r37_c7_7 = t_r37_c7_2 + t_r37_c7_3;
  assign t_r37_c7_8 = t_r37_c7_4 + p_38_6;
  assign t_r37_c7_9 = t_r37_c7_5 + t_r37_c7_6;
  assign t_r37_c7_10 = t_r37_c7_7 + t_r37_c7_8;
  assign t_r37_c7_11 = t_r37_c7_9 + t_r37_c7_10;
  assign t_r37_c7_12 = t_r37_c7_11 + p_38_8;
  assign out_37_7 = t_r37_c7_12 >> 4;

  assign t_r37_c8_0 = p_36_8 << 1;
  assign t_r37_c8_1 = p_37_7 << 1;
  assign t_r37_c8_2 = p_37_8 << 2;
  assign t_r37_c8_3 = p_37_9 << 1;
  assign t_r37_c8_4 = p_38_8 << 1;
  assign t_r37_c8_5 = t_r37_c8_0 + p_36_7;
  assign t_r37_c8_6 = t_r37_c8_1 + p_36_9;
  assign t_r37_c8_7 = t_r37_c8_2 + t_r37_c8_3;
  assign t_r37_c8_8 = t_r37_c8_4 + p_38_7;
  assign t_r37_c8_9 = t_r37_c8_5 + t_r37_c8_6;
  assign t_r37_c8_10 = t_r37_c8_7 + t_r37_c8_8;
  assign t_r37_c8_11 = t_r37_c8_9 + t_r37_c8_10;
  assign t_r37_c8_12 = t_r37_c8_11 + p_38_9;
  assign out_37_8 = t_r37_c8_12 >> 4;

  assign t_r37_c9_0 = p_36_9 << 1;
  assign t_r37_c9_1 = p_37_8 << 1;
  assign t_r37_c9_2 = p_37_9 << 2;
  assign t_r37_c9_3 = p_37_10 << 1;
  assign t_r37_c9_4 = p_38_9 << 1;
  assign t_r37_c9_5 = t_r37_c9_0 + p_36_8;
  assign t_r37_c9_6 = t_r37_c9_1 + p_36_10;
  assign t_r37_c9_7 = t_r37_c9_2 + t_r37_c9_3;
  assign t_r37_c9_8 = t_r37_c9_4 + p_38_8;
  assign t_r37_c9_9 = t_r37_c9_5 + t_r37_c9_6;
  assign t_r37_c9_10 = t_r37_c9_7 + t_r37_c9_8;
  assign t_r37_c9_11 = t_r37_c9_9 + t_r37_c9_10;
  assign t_r37_c9_12 = t_r37_c9_11 + p_38_10;
  assign out_37_9 = t_r37_c9_12 >> 4;

  assign t_r37_c10_0 = p_36_10 << 1;
  assign t_r37_c10_1 = p_37_9 << 1;
  assign t_r37_c10_2 = p_37_10 << 2;
  assign t_r37_c10_3 = p_37_11 << 1;
  assign t_r37_c10_4 = p_38_10 << 1;
  assign t_r37_c10_5 = t_r37_c10_0 + p_36_9;
  assign t_r37_c10_6 = t_r37_c10_1 + p_36_11;
  assign t_r37_c10_7 = t_r37_c10_2 + t_r37_c10_3;
  assign t_r37_c10_8 = t_r37_c10_4 + p_38_9;
  assign t_r37_c10_9 = t_r37_c10_5 + t_r37_c10_6;
  assign t_r37_c10_10 = t_r37_c10_7 + t_r37_c10_8;
  assign t_r37_c10_11 = t_r37_c10_9 + t_r37_c10_10;
  assign t_r37_c10_12 = t_r37_c10_11 + p_38_11;
  assign out_37_10 = t_r37_c10_12 >> 4;

  assign t_r37_c11_0 = p_36_11 << 1;
  assign t_r37_c11_1 = p_37_10 << 1;
  assign t_r37_c11_2 = p_37_11 << 2;
  assign t_r37_c11_3 = p_37_12 << 1;
  assign t_r37_c11_4 = p_38_11 << 1;
  assign t_r37_c11_5 = t_r37_c11_0 + p_36_10;
  assign t_r37_c11_6 = t_r37_c11_1 + p_36_12;
  assign t_r37_c11_7 = t_r37_c11_2 + t_r37_c11_3;
  assign t_r37_c11_8 = t_r37_c11_4 + p_38_10;
  assign t_r37_c11_9 = t_r37_c11_5 + t_r37_c11_6;
  assign t_r37_c11_10 = t_r37_c11_7 + t_r37_c11_8;
  assign t_r37_c11_11 = t_r37_c11_9 + t_r37_c11_10;
  assign t_r37_c11_12 = t_r37_c11_11 + p_38_12;
  assign out_37_11 = t_r37_c11_12 >> 4;

  assign t_r37_c12_0 = p_36_12 << 1;
  assign t_r37_c12_1 = p_37_11 << 1;
  assign t_r37_c12_2 = p_37_12 << 2;
  assign t_r37_c12_3 = p_37_13 << 1;
  assign t_r37_c12_4 = p_38_12 << 1;
  assign t_r37_c12_5 = t_r37_c12_0 + p_36_11;
  assign t_r37_c12_6 = t_r37_c12_1 + p_36_13;
  assign t_r37_c12_7 = t_r37_c12_2 + t_r37_c12_3;
  assign t_r37_c12_8 = t_r37_c12_4 + p_38_11;
  assign t_r37_c12_9 = t_r37_c12_5 + t_r37_c12_6;
  assign t_r37_c12_10 = t_r37_c12_7 + t_r37_c12_8;
  assign t_r37_c12_11 = t_r37_c12_9 + t_r37_c12_10;
  assign t_r37_c12_12 = t_r37_c12_11 + p_38_13;
  assign out_37_12 = t_r37_c12_12 >> 4;

  assign t_r37_c13_0 = p_36_13 << 1;
  assign t_r37_c13_1 = p_37_12 << 1;
  assign t_r37_c13_2 = p_37_13 << 2;
  assign t_r37_c13_3 = p_37_14 << 1;
  assign t_r37_c13_4 = p_38_13 << 1;
  assign t_r37_c13_5 = t_r37_c13_0 + p_36_12;
  assign t_r37_c13_6 = t_r37_c13_1 + p_36_14;
  assign t_r37_c13_7 = t_r37_c13_2 + t_r37_c13_3;
  assign t_r37_c13_8 = t_r37_c13_4 + p_38_12;
  assign t_r37_c13_9 = t_r37_c13_5 + t_r37_c13_6;
  assign t_r37_c13_10 = t_r37_c13_7 + t_r37_c13_8;
  assign t_r37_c13_11 = t_r37_c13_9 + t_r37_c13_10;
  assign t_r37_c13_12 = t_r37_c13_11 + p_38_14;
  assign out_37_13 = t_r37_c13_12 >> 4;

  assign t_r37_c14_0 = p_36_14 << 1;
  assign t_r37_c14_1 = p_37_13 << 1;
  assign t_r37_c14_2 = p_37_14 << 2;
  assign t_r37_c14_3 = p_37_15 << 1;
  assign t_r37_c14_4 = p_38_14 << 1;
  assign t_r37_c14_5 = t_r37_c14_0 + p_36_13;
  assign t_r37_c14_6 = t_r37_c14_1 + p_36_15;
  assign t_r37_c14_7 = t_r37_c14_2 + t_r37_c14_3;
  assign t_r37_c14_8 = t_r37_c14_4 + p_38_13;
  assign t_r37_c14_9 = t_r37_c14_5 + t_r37_c14_6;
  assign t_r37_c14_10 = t_r37_c14_7 + t_r37_c14_8;
  assign t_r37_c14_11 = t_r37_c14_9 + t_r37_c14_10;
  assign t_r37_c14_12 = t_r37_c14_11 + p_38_15;
  assign out_37_14 = t_r37_c14_12 >> 4;

  assign t_r37_c15_0 = p_36_15 << 1;
  assign t_r37_c15_1 = p_37_14 << 1;
  assign t_r37_c15_2 = p_37_15 << 2;
  assign t_r37_c15_3 = p_37_16 << 1;
  assign t_r37_c15_4 = p_38_15 << 1;
  assign t_r37_c15_5 = t_r37_c15_0 + p_36_14;
  assign t_r37_c15_6 = t_r37_c15_1 + p_36_16;
  assign t_r37_c15_7 = t_r37_c15_2 + t_r37_c15_3;
  assign t_r37_c15_8 = t_r37_c15_4 + p_38_14;
  assign t_r37_c15_9 = t_r37_c15_5 + t_r37_c15_6;
  assign t_r37_c15_10 = t_r37_c15_7 + t_r37_c15_8;
  assign t_r37_c15_11 = t_r37_c15_9 + t_r37_c15_10;
  assign t_r37_c15_12 = t_r37_c15_11 + p_38_16;
  assign out_37_15 = t_r37_c15_12 >> 4;

  assign t_r37_c16_0 = p_36_16 << 1;
  assign t_r37_c16_1 = p_37_15 << 1;
  assign t_r37_c16_2 = p_37_16 << 2;
  assign t_r37_c16_3 = p_37_17 << 1;
  assign t_r37_c16_4 = p_38_16 << 1;
  assign t_r37_c16_5 = t_r37_c16_0 + p_36_15;
  assign t_r37_c16_6 = t_r37_c16_1 + p_36_17;
  assign t_r37_c16_7 = t_r37_c16_2 + t_r37_c16_3;
  assign t_r37_c16_8 = t_r37_c16_4 + p_38_15;
  assign t_r37_c16_9 = t_r37_c16_5 + t_r37_c16_6;
  assign t_r37_c16_10 = t_r37_c16_7 + t_r37_c16_8;
  assign t_r37_c16_11 = t_r37_c16_9 + t_r37_c16_10;
  assign t_r37_c16_12 = t_r37_c16_11 + p_38_17;
  assign out_37_16 = t_r37_c16_12 >> 4;

  assign t_r37_c17_0 = p_36_17 << 1;
  assign t_r37_c17_1 = p_37_16 << 1;
  assign t_r37_c17_2 = p_37_17 << 2;
  assign t_r37_c17_3 = p_37_18 << 1;
  assign t_r37_c17_4 = p_38_17 << 1;
  assign t_r37_c17_5 = t_r37_c17_0 + p_36_16;
  assign t_r37_c17_6 = t_r37_c17_1 + p_36_18;
  assign t_r37_c17_7 = t_r37_c17_2 + t_r37_c17_3;
  assign t_r37_c17_8 = t_r37_c17_4 + p_38_16;
  assign t_r37_c17_9 = t_r37_c17_5 + t_r37_c17_6;
  assign t_r37_c17_10 = t_r37_c17_7 + t_r37_c17_8;
  assign t_r37_c17_11 = t_r37_c17_9 + t_r37_c17_10;
  assign t_r37_c17_12 = t_r37_c17_11 + p_38_18;
  assign out_37_17 = t_r37_c17_12 >> 4;

  assign t_r37_c18_0 = p_36_18 << 1;
  assign t_r37_c18_1 = p_37_17 << 1;
  assign t_r37_c18_2 = p_37_18 << 2;
  assign t_r37_c18_3 = p_37_19 << 1;
  assign t_r37_c18_4 = p_38_18 << 1;
  assign t_r37_c18_5 = t_r37_c18_0 + p_36_17;
  assign t_r37_c18_6 = t_r37_c18_1 + p_36_19;
  assign t_r37_c18_7 = t_r37_c18_2 + t_r37_c18_3;
  assign t_r37_c18_8 = t_r37_c18_4 + p_38_17;
  assign t_r37_c18_9 = t_r37_c18_5 + t_r37_c18_6;
  assign t_r37_c18_10 = t_r37_c18_7 + t_r37_c18_8;
  assign t_r37_c18_11 = t_r37_c18_9 + t_r37_c18_10;
  assign t_r37_c18_12 = t_r37_c18_11 + p_38_19;
  assign out_37_18 = t_r37_c18_12 >> 4;

  assign t_r37_c19_0 = p_36_19 << 1;
  assign t_r37_c19_1 = p_37_18 << 1;
  assign t_r37_c19_2 = p_37_19 << 2;
  assign t_r37_c19_3 = p_37_20 << 1;
  assign t_r37_c19_4 = p_38_19 << 1;
  assign t_r37_c19_5 = t_r37_c19_0 + p_36_18;
  assign t_r37_c19_6 = t_r37_c19_1 + p_36_20;
  assign t_r37_c19_7 = t_r37_c19_2 + t_r37_c19_3;
  assign t_r37_c19_8 = t_r37_c19_4 + p_38_18;
  assign t_r37_c19_9 = t_r37_c19_5 + t_r37_c19_6;
  assign t_r37_c19_10 = t_r37_c19_7 + t_r37_c19_8;
  assign t_r37_c19_11 = t_r37_c19_9 + t_r37_c19_10;
  assign t_r37_c19_12 = t_r37_c19_11 + p_38_20;
  assign out_37_19 = t_r37_c19_12 >> 4;

  assign t_r37_c20_0 = p_36_20 << 1;
  assign t_r37_c20_1 = p_37_19 << 1;
  assign t_r37_c20_2 = p_37_20 << 2;
  assign t_r37_c20_3 = p_37_21 << 1;
  assign t_r37_c20_4 = p_38_20 << 1;
  assign t_r37_c20_5 = t_r37_c20_0 + p_36_19;
  assign t_r37_c20_6 = t_r37_c20_1 + p_36_21;
  assign t_r37_c20_7 = t_r37_c20_2 + t_r37_c20_3;
  assign t_r37_c20_8 = t_r37_c20_4 + p_38_19;
  assign t_r37_c20_9 = t_r37_c20_5 + t_r37_c20_6;
  assign t_r37_c20_10 = t_r37_c20_7 + t_r37_c20_8;
  assign t_r37_c20_11 = t_r37_c20_9 + t_r37_c20_10;
  assign t_r37_c20_12 = t_r37_c20_11 + p_38_21;
  assign out_37_20 = t_r37_c20_12 >> 4;

  assign t_r37_c21_0 = p_36_21 << 1;
  assign t_r37_c21_1 = p_37_20 << 1;
  assign t_r37_c21_2 = p_37_21 << 2;
  assign t_r37_c21_3 = p_37_22 << 1;
  assign t_r37_c21_4 = p_38_21 << 1;
  assign t_r37_c21_5 = t_r37_c21_0 + p_36_20;
  assign t_r37_c21_6 = t_r37_c21_1 + p_36_22;
  assign t_r37_c21_7 = t_r37_c21_2 + t_r37_c21_3;
  assign t_r37_c21_8 = t_r37_c21_4 + p_38_20;
  assign t_r37_c21_9 = t_r37_c21_5 + t_r37_c21_6;
  assign t_r37_c21_10 = t_r37_c21_7 + t_r37_c21_8;
  assign t_r37_c21_11 = t_r37_c21_9 + t_r37_c21_10;
  assign t_r37_c21_12 = t_r37_c21_11 + p_38_22;
  assign out_37_21 = t_r37_c21_12 >> 4;

  assign t_r37_c22_0 = p_36_22 << 1;
  assign t_r37_c22_1 = p_37_21 << 1;
  assign t_r37_c22_2 = p_37_22 << 2;
  assign t_r37_c22_3 = p_37_23 << 1;
  assign t_r37_c22_4 = p_38_22 << 1;
  assign t_r37_c22_5 = t_r37_c22_0 + p_36_21;
  assign t_r37_c22_6 = t_r37_c22_1 + p_36_23;
  assign t_r37_c22_7 = t_r37_c22_2 + t_r37_c22_3;
  assign t_r37_c22_8 = t_r37_c22_4 + p_38_21;
  assign t_r37_c22_9 = t_r37_c22_5 + t_r37_c22_6;
  assign t_r37_c22_10 = t_r37_c22_7 + t_r37_c22_8;
  assign t_r37_c22_11 = t_r37_c22_9 + t_r37_c22_10;
  assign t_r37_c22_12 = t_r37_c22_11 + p_38_23;
  assign out_37_22 = t_r37_c22_12 >> 4;

  assign t_r37_c23_0 = p_36_23 << 1;
  assign t_r37_c23_1 = p_37_22 << 1;
  assign t_r37_c23_2 = p_37_23 << 2;
  assign t_r37_c23_3 = p_37_24 << 1;
  assign t_r37_c23_4 = p_38_23 << 1;
  assign t_r37_c23_5 = t_r37_c23_0 + p_36_22;
  assign t_r37_c23_6 = t_r37_c23_1 + p_36_24;
  assign t_r37_c23_7 = t_r37_c23_2 + t_r37_c23_3;
  assign t_r37_c23_8 = t_r37_c23_4 + p_38_22;
  assign t_r37_c23_9 = t_r37_c23_5 + t_r37_c23_6;
  assign t_r37_c23_10 = t_r37_c23_7 + t_r37_c23_8;
  assign t_r37_c23_11 = t_r37_c23_9 + t_r37_c23_10;
  assign t_r37_c23_12 = t_r37_c23_11 + p_38_24;
  assign out_37_23 = t_r37_c23_12 >> 4;

  assign t_r37_c24_0 = p_36_24 << 1;
  assign t_r37_c24_1 = p_37_23 << 1;
  assign t_r37_c24_2 = p_37_24 << 2;
  assign t_r37_c24_3 = p_37_25 << 1;
  assign t_r37_c24_4 = p_38_24 << 1;
  assign t_r37_c24_5 = t_r37_c24_0 + p_36_23;
  assign t_r37_c24_6 = t_r37_c24_1 + p_36_25;
  assign t_r37_c24_7 = t_r37_c24_2 + t_r37_c24_3;
  assign t_r37_c24_8 = t_r37_c24_4 + p_38_23;
  assign t_r37_c24_9 = t_r37_c24_5 + t_r37_c24_6;
  assign t_r37_c24_10 = t_r37_c24_7 + t_r37_c24_8;
  assign t_r37_c24_11 = t_r37_c24_9 + t_r37_c24_10;
  assign t_r37_c24_12 = t_r37_c24_11 + p_38_25;
  assign out_37_24 = t_r37_c24_12 >> 4;

  assign t_r37_c25_0 = p_36_25 << 1;
  assign t_r37_c25_1 = p_37_24 << 1;
  assign t_r37_c25_2 = p_37_25 << 2;
  assign t_r37_c25_3 = p_37_26 << 1;
  assign t_r37_c25_4 = p_38_25 << 1;
  assign t_r37_c25_5 = t_r37_c25_0 + p_36_24;
  assign t_r37_c25_6 = t_r37_c25_1 + p_36_26;
  assign t_r37_c25_7 = t_r37_c25_2 + t_r37_c25_3;
  assign t_r37_c25_8 = t_r37_c25_4 + p_38_24;
  assign t_r37_c25_9 = t_r37_c25_5 + t_r37_c25_6;
  assign t_r37_c25_10 = t_r37_c25_7 + t_r37_c25_8;
  assign t_r37_c25_11 = t_r37_c25_9 + t_r37_c25_10;
  assign t_r37_c25_12 = t_r37_c25_11 + p_38_26;
  assign out_37_25 = t_r37_c25_12 >> 4;

  assign t_r37_c26_0 = p_36_26 << 1;
  assign t_r37_c26_1 = p_37_25 << 1;
  assign t_r37_c26_2 = p_37_26 << 2;
  assign t_r37_c26_3 = p_37_27 << 1;
  assign t_r37_c26_4 = p_38_26 << 1;
  assign t_r37_c26_5 = t_r37_c26_0 + p_36_25;
  assign t_r37_c26_6 = t_r37_c26_1 + p_36_27;
  assign t_r37_c26_7 = t_r37_c26_2 + t_r37_c26_3;
  assign t_r37_c26_8 = t_r37_c26_4 + p_38_25;
  assign t_r37_c26_9 = t_r37_c26_5 + t_r37_c26_6;
  assign t_r37_c26_10 = t_r37_c26_7 + t_r37_c26_8;
  assign t_r37_c26_11 = t_r37_c26_9 + t_r37_c26_10;
  assign t_r37_c26_12 = t_r37_c26_11 + p_38_27;
  assign out_37_26 = t_r37_c26_12 >> 4;

  assign t_r37_c27_0 = p_36_27 << 1;
  assign t_r37_c27_1 = p_37_26 << 1;
  assign t_r37_c27_2 = p_37_27 << 2;
  assign t_r37_c27_3 = p_37_28 << 1;
  assign t_r37_c27_4 = p_38_27 << 1;
  assign t_r37_c27_5 = t_r37_c27_0 + p_36_26;
  assign t_r37_c27_6 = t_r37_c27_1 + p_36_28;
  assign t_r37_c27_7 = t_r37_c27_2 + t_r37_c27_3;
  assign t_r37_c27_8 = t_r37_c27_4 + p_38_26;
  assign t_r37_c27_9 = t_r37_c27_5 + t_r37_c27_6;
  assign t_r37_c27_10 = t_r37_c27_7 + t_r37_c27_8;
  assign t_r37_c27_11 = t_r37_c27_9 + t_r37_c27_10;
  assign t_r37_c27_12 = t_r37_c27_11 + p_38_28;
  assign out_37_27 = t_r37_c27_12 >> 4;

  assign t_r37_c28_0 = p_36_28 << 1;
  assign t_r37_c28_1 = p_37_27 << 1;
  assign t_r37_c28_2 = p_37_28 << 2;
  assign t_r37_c28_3 = p_37_29 << 1;
  assign t_r37_c28_4 = p_38_28 << 1;
  assign t_r37_c28_5 = t_r37_c28_0 + p_36_27;
  assign t_r37_c28_6 = t_r37_c28_1 + p_36_29;
  assign t_r37_c28_7 = t_r37_c28_2 + t_r37_c28_3;
  assign t_r37_c28_8 = t_r37_c28_4 + p_38_27;
  assign t_r37_c28_9 = t_r37_c28_5 + t_r37_c28_6;
  assign t_r37_c28_10 = t_r37_c28_7 + t_r37_c28_8;
  assign t_r37_c28_11 = t_r37_c28_9 + t_r37_c28_10;
  assign t_r37_c28_12 = t_r37_c28_11 + p_38_29;
  assign out_37_28 = t_r37_c28_12 >> 4;

  assign t_r37_c29_0 = p_36_29 << 1;
  assign t_r37_c29_1 = p_37_28 << 1;
  assign t_r37_c29_2 = p_37_29 << 2;
  assign t_r37_c29_3 = p_37_30 << 1;
  assign t_r37_c29_4 = p_38_29 << 1;
  assign t_r37_c29_5 = t_r37_c29_0 + p_36_28;
  assign t_r37_c29_6 = t_r37_c29_1 + p_36_30;
  assign t_r37_c29_7 = t_r37_c29_2 + t_r37_c29_3;
  assign t_r37_c29_8 = t_r37_c29_4 + p_38_28;
  assign t_r37_c29_9 = t_r37_c29_5 + t_r37_c29_6;
  assign t_r37_c29_10 = t_r37_c29_7 + t_r37_c29_8;
  assign t_r37_c29_11 = t_r37_c29_9 + t_r37_c29_10;
  assign t_r37_c29_12 = t_r37_c29_11 + p_38_30;
  assign out_37_29 = t_r37_c29_12 >> 4;

  assign t_r37_c30_0 = p_36_30 << 1;
  assign t_r37_c30_1 = p_37_29 << 1;
  assign t_r37_c30_2 = p_37_30 << 2;
  assign t_r37_c30_3 = p_37_31 << 1;
  assign t_r37_c30_4 = p_38_30 << 1;
  assign t_r37_c30_5 = t_r37_c30_0 + p_36_29;
  assign t_r37_c30_6 = t_r37_c30_1 + p_36_31;
  assign t_r37_c30_7 = t_r37_c30_2 + t_r37_c30_3;
  assign t_r37_c30_8 = t_r37_c30_4 + p_38_29;
  assign t_r37_c30_9 = t_r37_c30_5 + t_r37_c30_6;
  assign t_r37_c30_10 = t_r37_c30_7 + t_r37_c30_8;
  assign t_r37_c30_11 = t_r37_c30_9 + t_r37_c30_10;
  assign t_r37_c30_12 = t_r37_c30_11 + p_38_31;
  assign out_37_30 = t_r37_c30_12 >> 4;

  assign t_r37_c31_0 = p_36_31 << 1;
  assign t_r37_c31_1 = p_37_30 << 1;
  assign t_r37_c31_2 = p_37_31 << 2;
  assign t_r37_c31_3 = p_37_32 << 1;
  assign t_r37_c31_4 = p_38_31 << 1;
  assign t_r37_c31_5 = t_r37_c31_0 + p_36_30;
  assign t_r37_c31_6 = t_r37_c31_1 + p_36_32;
  assign t_r37_c31_7 = t_r37_c31_2 + t_r37_c31_3;
  assign t_r37_c31_8 = t_r37_c31_4 + p_38_30;
  assign t_r37_c31_9 = t_r37_c31_5 + t_r37_c31_6;
  assign t_r37_c31_10 = t_r37_c31_7 + t_r37_c31_8;
  assign t_r37_c31_11 = t_r37_c31_9 + t_r37_c31_10;
  assign t_r37_c31_12 = t_r37_c31_11 + p_38_32;
  assign out_37_31 = t_r37_c31_12 >> 4;

  assign t_r37_c32_0 = p_36_32 << 1;
  assign t_r37_c32_1 = p_37_31 << 1;
  assign t_r37_c32_2 = p_37_32 << 2;
  assign t_r37_c32_3 = p_37_33 << 1;
  assign t_r37_c32_4 = p_38_32 << 1;
  assign t_r37_c32_5 = t_r37_c32_0 + p_36_31;
  assign t_r37_c32_6 = t_r37_c32_1 + p_36_33;
  assign t_r37_c32_7 = t_r37_c32_2 + t_r37_c32_3;
  assign t_r37_c32_8 = t_r37_c32_4 + p_38_31;
  assign t_r37_c32_9 = t_r37_c32_5 + t_r37_c32_6;
  assign t_r37_c32_10 = t_r37_c32_7 + t_r37_c32_8;
  assign t_r37_c32_11 = t_r37_c32_9 + t_r37_c32_10;
  assign t_r37_c32_12 = t_r37_c32_11 + p_38_33;
  assign out_37_32 = t_r37_c32_12 >> 4;

  assign t_r37_c33_0 = p_36_33 << 1;
  assign t_r37_c33_1 = p_37_32 << 1;
  assign t_r37_c33_2 = p_37_33 << 2;
  assign t_r37_c33_3 = p_37_34 << 1;
  assign t_r37_c33_4 = p_38_33 << 1;
  assign t_r37_c33_5 = t_r37_c33_0 + p_36_32;
  assign t_r37_c33_6 = t_r37_c33_1 + p_36_34;
  assign t_r37_c33_7 = t_r37_c33_2 + t_r37_c33_3;
  assign t_r37_c33_8 = t_r37_c33_4 + p_38_32;
  assign t_r37_c33_9 = t_r37_c33_5 + t_r37_c33_6;
  assign t_r37_c33_10 = t_r37_c33_7 + t_r37_c33_8;
  assign t_r37_c33_11 = t_r37_c33_9 + t_r37_c33_10;
  assign t_r37_c33_12 = t_r37_c33_11 + p_38_34;
  assign out_37_33 = t_r37_c33_12 >> 4;

  assign t_r37_c34_0 = p_36_34 << 1;
  assign t_r37_c34_1 = p_37_33 << 1;
  assign t_r37_c34_2 = p_37_34 << 2;
  assign t_r37_c34_3 = p_37_35 << 1;
  assign t_r37_c34_4 = p_38_34 << 1;
  assign t_r37_c34_5 = t_r37_c34_0 + p_36_33;
  assign t_r37_c34_6 = t_r37_c34_1 + p_36_35;
  assign t_r37_c34_7 = t_r37_c34_2 + t_r37_c34_3;
  assign t_r37_c34_8 = t_r37_c34_4 + p_38_33;
  assign t_r37_c34_9 = t_r37_c34_5 + t_r37_c34_6;
  assign t_r37_c34_10 = t_r37_c34_7 + t_r37_c34_8;
  assign t_r37_c34_11 = t_r37_c34_9 + t_r37_c34_10;
  assign t_r37_c34_12 = t_r37_c34_11 + p_38_35;
  assign out_37_34 = t_r37_c34_12 >> 4;

  assign t_r37_c35_0 = p_36_35 << 1;
  assign t_r37_c35_1 = p_37_34 << 1;
  assign t_r37_c35_2 = p_37_35 << 2;
  assign t_r37_c35_3 = p_37_36 << 1;
  assign t_r37_c35_4 = p_38_35 << 1;
  assign t_r37_c35_5 = t_r37_c35_0 + p_36_34;
  assign t_r37_c35_6 = t_r37_c35_1 + p_36_36;
  assign t_r37_c35_7 = t_r37_c35_2 + t_r37_c35_3;
  assign t_r37_c35_8 = t_r37_c35_4 + p_38_34;
  assign t_r37_c35_9 = t_r37_c35_5 + t_r37_c35_6;
  assign t_r37_c35_10 = t_r37_c35_7 + t_r37_c35_8;
  assign t_r37_c35_11 = t_r37_c35_9 + t_r37_c35_10;
  assign t_r37_c35_12 = t_r37_c35_11 + p_38_36;
  assign out_37_35 = t_r37_c35_12 >> 4;

  assign t_r37_c36_0 = p_36_36 << 1;
  assign t_r37_c36_1 = p_37_35 << 1;
  assign t_r37_c36_2 = p_37_36 << 2;
  assign t_r37_c36_3 = p_37_37 << 1;
  assign t_r37_c36_4 = p_38_36 << 1;
  assign t_r37_c36_5 = t_r37_c36_0 + p_36_35;
  assign t_r37_c36_6 = t_r37_c36_1 + p_36_37;
  assign t_r37_c36_7 = t_r37_c36_2 + t_r37_c36_3;
  assign t_r37_c36_8 = t_r37_c36_4 + p_38_35;
  assign t_r37_c36_9 = t_r37_c36_5 + t_r37_c36_6;
  assign t_r37_c36_10 = t_r37_c36_7 + t_r37_c36_8;
  assign t_r37_c36_11 = t_r37_c36_9 + t_r37_c36_10;
  assign t_r37_c36_12 = t_r37_c36_11 + p_38_37;
  assign out_37_36 = t_r37_c36_12 >> 4;

  assign t_r37_c37_0 = p_36_37 << 1;
  assign t_r37_c37_1 = p_37_36 << 1;
  assign t_r37_c37_2 = p_37_37 << 2;
  assign t_r37_c37_3 = p_37_38 << 1;
  assign t_r37_c37_4 = p_38_37 << 1;
  assign t_r37_c37_5 = t_r37_c37_0 + p_36_36;
  assign t_r37_c37_6 = t_r37_c37_1 + p_36_38;
  assign t_r37_c37_7 = t_r37_c37_2 + t_r37_c37_3;
  assign t_r37_c37_8 = t_r37_c37_4 + p_38_36;
  assign t_r37_c37_9 = t_r37_c37_5 + t_r37_c37_6;
  assign t_r37_c37_10 = t_r37_c37_7 + t_r37_c37_8;
  assign t_r37_c37_11 = t_r37_c37_9 + t_r37_c37_10;
  assign t_r37_c37_12 = t_r37_c37_11 + p_38_38;
  assign out_37_37 = t_r37_c37_12 >> 4;

  assign t_r37_c38_0 = p_36_38 << 1;
  assign t_r37_c38_1 = p_37_37 << 1;
  assign t_r37_c38_2 = p_37_38 << 2;
  assign t_r37_c38_3 = p_37_39 << 1;
  assign t_r37_c38_4 = p_38_38 << 1;
  assign t_r37_c38_5 = t_r37_c38_0 + p_36_37;
  assign t_r37_c38_6 = t_r37_c38_1 + p_36_39;
  assign t_r37_c38_7 = t_r37_c38_2 + t_r37_c38_3;
  assign t_r37_c38_8 = t_r37_c38_4 + p_38_37;
  assign t_r37_c38_9 = t_r37_c38_5 + t_r37_c38_6;
  assign t_r37_c38_10 = t_r37_c38_7 + t_r37_c38_8;
  assign t_r37_c38_11 = t_r37_c38_9 + t_r37_c38_10;
  assign t_r37_c38_12 = t_r37_c38_11 + p_38_39;
  assign out_37_38 = t_r37_c38_12 >> 4;

  assign t_r37_c39_0 = p_36_39 << 1;
  assign t_r37_c39_1 = p_37_38 << 1;
  assign t_r37_c39_2 = p_37_39 << 2;
  assign t_r37_c39_3 = p_37_40 << 1;
  assign t_r37_c39_4 = p_38_39 << 1;
  assign t_r37_c39_5 = t_r37_c39_0 + p_36_38;
  assign t_r37_c39_6 = t_r37_c39_1 + p_36_40;
  assign t_r37_c39_7 = t_r37_c39_2 + t_r37_c39_3;
  assign t_r37_c39_8 = t_r37_c39_4 + p_38_38;
  assign t_r37_c39_9 = t_r37_c39_5 + t_r37_c39_6;
  assign t_r37_c39_10 = t_r37_c39_7 + t_r37_c39_8;
  assign t_r37_c39_11 = t_r37_c39_9 + t_r37_c39_10;
  assign t_r37_c39_12 = t_r37_c39_11 + p_38_40;
  assign out_37_39 = t_r37_c39_12 >> 4;

  assign t_r37_c40_0 = p_36_40 << 1;
  assign t_r37_c40_1 = p_37_39 << 1;
  assign t_r37_c40_2 = p_37_40 << 2;
  assign t_r37_c40_3 = p_37_41 << 1;
  assign t_r37_c40_4 = p_38_40 << 1;
  assign t_r37_c40_5 = t_r37_c40_0 + p_36_39;
  assign t_r37_c40_6 = t_r37_c40_1 + p_36_41;
  assign t_r37_c40_7 = t_r37_c40_2 + t_r37_c40_3;
  assign t_r37_c40_8 = t_r37_c40_4 + p_38_39;
  assign t_r37_c40_9 = t_r37_c40_5 + t_r37_c40_6;
  assign t_r37_c40_10 = t_r37_c40_7 + t_r37_c40_8;
  assign t_r37_c40_11 = t_r37_c40_9 + t_r37_c40_10;
  assign t_r37_c40_12 = t_r37_c40_11 + p_38_41;
  assign out_37_40 = t_r37_c40_12 >> 4;

  assign t_r37_c41_0 = p_36_41 << 1;
  assign t_r37_c41_1 = p_37_40 << 1;
  assign t_r37_c41_2 = p_37_41 << 2;
  assign t_r37_c41_3 = p_37_42 << 1;
  assign t_r37_c41_4 = p_38_41 << 1;
  assign t_r37_c41_5 = t_r37_c41_0 + p_36_40;
  assign t_r37_c41_6 = t_r37_c41_1 + p_36_42;
  assign t_r37_c41_7 = t_r37_c41_2 + t_r37_c41_3;
  assign t_r37_c41_8 = t_r37_c41_4 + p_38_40;
  assign t_r37_c41_9 = t_r37_c41_5 + t_r37_c41_6;
  assign t_r37_c41_10 = t_r37_c41_7 + t_r37_c41_8;
  assign t_r37_c41_11 = t_r37_c41_9 + t_r37_c41_10;
  assign t_r37_c41_12 = t_r37_c41_11 + p_38_42;
  assign out_37_41 = t_r37_c41_12 >> 4;

  assign t_r37_c42_0 = p_36_42 << 1;
  assign t_r37_c42_1 = p_37_41 << 1;
  assign t_r37_c42_2 = p_37_42 << 2;
  assign t_r37_c42_3 = p_37_43 << 1;
  assign t_r37_c42_4 = p_38_42 << 1;
  assign t_r37_c42_5 = t_r37_c42_0 + p_36_41;
  assign t_r37_c42_6 = t_r37_c42_1 + p_36_43;
  assign t_r37_c42_7 = t_r37_c42_2 + t_r37_c42_3;
  assign t_r37_c42_8 = t_r37_c42_4 + p_38_41;
  assign t_r37_c42_9 = t_r37_c42_5 + t_r37_c42_6;
  assign t_r37_c42_10 = t_r37_c42_7 + t_r37_c42_8;
  assign t_r37_c42_11 = t_r37_c42_9 + t_r37_c42_10;
  assign t_r37_c42_12 = t_r37_c42_11 + p_38_43;
  assign out_37_42 = t_r37_c42_12 >> 4;

  assign t_r37_c43_0 = p_36_43 << 1;
  assign t_r37_c43_1 = p_37_42 << 1;
  assign t_r37_c43_2 = p_37_43 << 2;
  assign t_r37_c43_3 = p_37_44 << 1;
  assign t_r37_c43_4 = p_38_43 << 1;
  assign t_r37_c43_5 = t_r37_c43_0 + p_36_42;
  assign t_r37_c43_6 = t_r37_c43_1 + p_36_44;
  assign t_r37_c43_7 = t_r37_c43_2 + t_r37_c43_3;
  assign t_r37_c43_8 = t_r37_c43_4 + p_38_42;
  assign t_r37_c43_9 = t_r37_c43_5 + t_r37_c43_6;
  assign t_r37_c43_10 = t_r37_c43_7 + t_r37_c43_8;
  assign t_r37_c43_11 = t_r37_c43_9 + t_r37_c43_10;
  assign t_r37_c43_12 = t_r37_c43_11 + p_38_44;
  assign out_37_43 = t_r37_c43_12 >> 4;

  assign t_r37_c44_0 = p_36_44 << 1;
  assign t_r37_c44_1 = p_37_43 << 1;
  assign t_r37_c44_2 = p_37_44 << 2;
  assign t_r37_c44_3 = p_37_45 << 1;
  assign t_r37_c44_4 = p_38_44 << 1;
  assign t_r37_c44_5 = t_r37_c44_0 + p_36_43;
  assign t_r37_c44_6 = t_r37_c44_1 + p_36_45;
  assign t_r37_c44_7 = t_r37_c44_2 + t_r37_c44_3;
  assign t_r37_c44_8 = t_r37_c44_4 + p_38_43;
  assign t_r37_c44_9 = t_r37_c44_5 + t_r37_c44_6;
  assign t_r37_c44_10 = t_r37_c44_7 + t_r37_c44_8;
  assign t_r37_c44_11 = t_r37_c44_9 + t_r37_c44_10;
  assign t_r37_c44_12 = t_r37_c44_11 + p_38_45;
  assign out_37_44 = t_r37_c44_12 >> 4;

  assign t_r37_c45_0 = p_36_45 << 1;
  assign t_r37_c45_1 = p_37_44 << 1;
  assign t_r37_c45_2 = p_37_45 << 2;
  assign t_r37_c45_3 = p_37_46 << 1;
  assign t_r37_c45_4 = p_38_45 << 1;
  assign t_r37_c45_5 = t_r37_c45_0 + p_36_44;
  assign t_r37_c45_6 = t_r37_c45_1 + p_36_46;
  assign t_r37_c45_7 = t_r37_c45_2 + t_r37_c45_3;
  assign t_r37_c45_8 = t_r37_c45_4 + p_38_44;
  assign t_r37_c45_9 = t_r37_c45_5 + t_r37_c45_6;
  assign t_r37_c45_10 = t_r37_c45_7 + t_r37_c45_8;
  assign t_r37_c45_11 = t_r37_c45_9 + t_r37_c45_10;
  assign t_r37_c45_12 = t_r37_c45_11 + p_38_46;
  assign out_37_45 = t_r37_c45_12 >> 4;

  assign t_r37_c46_0 = p_36_46 << 1;
  assign t_r37_c46_1 = p_37_45 << 1;
  assign t_r37_c46_2 = p_37_46 << 2;
  assign t_r37_c46_3 = p_37_47 << 1;
  assign t_r37_c46_4 = p_38_46 << 1;
  assign t_r37_c46_5 = t_r37_c46_0 + p_36_45;
  assign t_r37_c46_6 = t_r37_c46_1 + p_36_47;
  assign t_r37_c46_7 = t_r37_c46_2 + t_r37_c46_3;
  assign t_r37_c46_8 = t_r37_c46_4 + p_38_45;
  assign t_r37_c46_9 = t_r37_c46_5 + t_r37_c46_6;
  assign t_r37_c46_10 = t_r37_c46_7 + t_r37_c46_8;
  assign t_r37_c46_11 = t_r37_c46_9 + t_r37_c46_10;
  assign t_r37_c46_12 = t_r37_c46_11 + p_38_47;
  assign out_37_46 = t_r37_c46_12 >> 4;

  assign t_r37_c47_0 = p_36_47 << 1;
  assign t_r37_c47_1 = p_37_46 << 1;
  assign t_r37_c47_2 = p_37_47 << 2;
  assign t_r37_c47_3 = p_37_48 << 1;
  assign t_r37_c47_4 = p_38_47 << 1;
  assign t_r37_c47_5 = t_r37_c47_0 + p_36_46;
  assign t_r37_c47_6 = t_r37_c47_1 + p_36_48;
  assign t_r37_c47_7 = t_r37_c47_2 + t_r37_c47_3;
  assign t_r37_c47_8 = t_r37_c47_4 + p_38_46;
  assign t_r37_c47_9 = t_r37_c47_5 + t_r37_c47_6;
  assign t_r37_c47_10 = t_r37_c47_7 + t_r37_c47_8;
  assign t_r37_c47_11 = t_r37_c47_9 + t_r37_c47_10;
  assign t_r37_c47_12 = t_r37_c47_11 + p_38_48;
  assign out_37_47 = t_r37_c47_12 >> 4;

  assign t_r37_c48_0 = p_36_48 << 1;
  assign t_r37_c48_1 = p_37_47 << 1;
  assign t_r37_c48_2 = p_37_48 << 2;
  assign t_r37_c48_3 = p_37_49 << 1;
  assign t_r37_c48_4 = p_38_48 << 1;
  assign t_r37_c48_5 = t_r37_c48_0 + p_36_47;
  assign t_r37_c48_6 = t_r37_c48_1 + p_36_49;
  assign t_r37_c48_7 = t_r37_c48_2 + t_r37_c48_3;
  assign t_r37_c48_8 = t_r37_c48_4 + p_38_47;
  assign t_r37_c48_9 = t_r37_c48_5 + t_r37_c48_6;
  assign t_r37_c48_10 = t_r37_c48_7 + t_r37_c48_8;
  assign t_r37_c48_11 = t_r37_c48_9 + t_r37_c48_10;
  assign t_r37_c48_12 = t_r37_c48_11 + p_38_49;
  assign out_37_48 = t_r37_c48_12 >> 4;

  assign t_r37_c49_0 = p_36_49 << 1;
  assign t_r37_c49_1 = p_37_48 << 1;
  assign t_r37_c49_2 = p_37_49 << 2;
  assign t_r37_c49_3 = p_37_50 << 1;
  assign t_r37_c49_4 = p_38_49 << 1;
  assign t_r37_c49_5 = t_r37_c49_0 + p_36_48;
  assign t_r37_c49_6 = t_r37_c49_1 + p_36_50;
  assign t_r37_c49_7 = t_r37_c49_2 + t_r37_c49_3;
  assign t_r37_c49_8 = t_r37_c49_4 + p_38_48;
  assign t_r37_c49_9 = t_r37_c49_5 + t_r37_c49_6;
  assign t_r37_c49_10 = t_r37_c49_7 + t_r37_c49_8;
  assign t_r37_c49_11 = t_r37_c49_9 + t_r37_c49_10;
  assign t_r37_c49_12 = t_r37_c49_11 + p_38_50;
  assign out_37_49 = t_r37_c49_12 >> 4;

  assign t_r37_c50_0 = p_36_50 << 1;
  assign t_r37_c50_1 = p_37_49 << 1;
  assign t_r37_c50_2 = p_37_50 << 2;
  assign t_r37_c50_3 = p_37_51 << 1;
  assign t_r37_c50_4 = p_38_50 << 1;
  assign t_r37_c50_5 = t_r37_c50_0 + p_36_49;
  assign t_r37_c50_6 = t_r37_c50_1 + p_36_51;
  assign t_r37_c50_7 = t_r37_c50_2 + t_r37_c50_3;
  assign t_r37_c50_8 = t_r37_c50_4 + p_38_49;
  assign t_r37_c50_9 = t_r37_c50_5 + t_r37_c50_6;
  assign t_r37_c50_10 = t_r37_c50_7 + t_r37_c50_8;
  assign t_r37_c50_11 = t_r37_c50_9 + t_r37_c50_10;
  assign t_r37_c50_12 = t_r37_c50_11 + p_38_51;
  assign out_37_50 = t_r37_c50_12 >> 4;

  assign t_r37_c51_0 = p_36_51 << 1;
  assign t_r37_c51_1 = p_37_50 << 1;
  assign t_r37_c51_2 = p_37_51 << 2;
  assign t_r37_c51_3 = p_37_52 << 1;
  assign t_r37_c51_4 = p_38_51 << 1;
  assign t_r37_c51_5 = t_r37_c51_0 + p_36_50;
  assign t_r37_c51_6 = t_r37_c51_1 + p_36_52;
  assign t_r37_c51_7 = t_r37_c51_2 + t_r37_c51_3;
  assign t_r37_c51_8 = t_r37_c51_4 + p_38_50;
  assign t_r37_c51_9 = t_r37_c51_5 + t_r37_c51_6;
  assign t_r37_c51_10 = t_r37_c51_7 + t_r37_c51_8;
  assign t_r37_c51_11 = t_r37_c51_9 + t_r37_c51_10;
  assign t_r37_c51_12 = t_r37_c51_11 + p_38_52;
  assign out_37_51 = t_r37_c51_12 >> 4;

  assign t_r37_c52_0 = p_36_52 << 1;
  assign t_r37_c52_1 = p_37_51 << 1;
  assign t_r37_c52_2 = p_37_52 << 2;
  assign t_r37_c52_3 = p_37_53 << 1;
  assign t_r37_c52_4 = p_38_52 << 1;
  assign t_r37_c52_5 = t_r37_c52_0 + p_36_51;
  assign t_r37_c52_6 = t_r37_c52_1 + p_36_53;
  assign t_r37_c52_7 = t_r37_c52_2 + t_r37_c52_3;
  assign t_r37_c52_8 = t_r37_c52_4 + p_38_51;
  assign t_r37_c52_9 = t_r37_c52_5 + t_r37_c52_6;
  assign t_r37_c52_10 = t_r37_c52_7 + t_r37_c52_8;
  assign t_r37_c52_11 = t_r37_c52_9 + t_r37_c52_10;
  assign t_r37_c52_12 = t_r37_c52_11 + p_38_53;
  assign out_37_52 = t_r37_c52_12 >> 4;

  assign t_r37_c53_0 = p_36_53 << 1;
  assign t_r37_c53_1 = p_37_52 << 1;
  assign t_r37_c53_2 = p_37_53 << 2;
  assign t_r37_c53_3 = p_37_54 << 1;
  assign t_r37_c53_4 = p_38_53 << 1;
  assign t_r37_c53_5 = t_r37_c53_0 + p_36_52;
  assign t_r37_c53_6 = t_r37_c53_1 + p_36_54;
  assign t_r37_c53_7 = t_r37_c53_2 + t_r37_c53_3;
  assign t_r37_c53_8 = t_r37_c53_4 + p_38_52;
  assign t_r37_c53_9 = t_r37_c53_5 + t_r37_c53_6;
  assign t_r37_c53_10 = t_r37_c53_7 + t_r37_c53_8;
  assign t_r37_c53_11 = t_r37_c53_9 + t_r37_c53_10;
  assign t_r37_c53_12 = t_r37_c53_11 + p_38_54;
  assign out_37_53 = t_r37_c53_12 >> 4;

  assign t_r37_c54_0 = p_36_54 << 1;
  assign t_r37_c54_1 = p_37_53 << 1;
  assign t_r37_c54_2 = p_37_54 << 2;
  assign t_r37_c54_3 = p_37_55 << 1;
  assign t_r37_c54_4 = p_38_54 << 1;
  assign t_r37_c54_5 = t_r37_c54_0 + p_36_53;
  assign t_r37_c54_6 = t_r37_c54_1 + p_36_55;
  assign t_r37_c54_7 = t_r37_c54_2 + t_r37_c54_3;
  assign t_r37_c54_8 = t_r37_c54_4 + p_38_53;
  assign t_r37_c54_9 = t_r37_c54_5 + t_r37_c54_6;
  assign t_r37_c54_10 = t_r37_c54_7 + t_r37_c54_8;
  assign t_r37_c54_11 = t_r37_c54_9 + t_r37_c54_10;
  assign t_r37_c54_12 = t_r37_c54_11 + p_38_55;
  assign out_37_54 = t_r37_c54_12 >> 4;

  assign t_r37_c55_0 = p_36_55 << 1;
  assign t_r37_c55_1 = p_37_54 << 1;
  assign t_r37_c55_2 = p_37_55 << 2;
  assign t_r37_c55_3 = p_37_56 << 1;
  assign t_r37_c55_4 = p_38_55 << 1;
  assign t_r37_c55_5 = t_r37_c55_0 + p_36_54;
  assign t_r37_c55_6 = t_r37_c55_1 + p_36_56;
  assign t_r37_c55_7 = t_r37_c55_2 + t_r37_c55_3;
  assign t_r37_c55_8 = t_r37_c55_4 + p_38_54;
  assign t_r37_c55_9 = t_r37_c55_5 + t_r37_c55_6;
  assign t_r37_c55_10 = t_r37_c55_7 + t_r37_c55_8;
  assign t_r37_c55_11 = t_r37_c55_9 + t_r37_c55_10;
  assign t_r37_c55_12 = t_r37_c55_11 + p_38_56;
  assign out_37_55 = t_r37_c55_12 >> 4;

  assign t_r37_c56_0 = p_36_56 << 1;
  assign t_r37_c56_1 = p_37_55 << 1;
  assign t_r37_c56_2 = p_37_56 << 2;
  assign t_r37_c56_3 = p_37_57 << 1;
  assign t_r37_c56_4 = p_38_56 << 1;
  assign t_r37_c56_5 = t_r37_c56_0 + p_36_55;
  assign t_r37_c56_6 = t_r37_c56_1 + p_36_57;
  assign t_r37_c56_7 = t_r37_c56_2 + t_r37_c56_3;
  assign t_r37_c56_8 = t_r37_c56_4 + p_38_55;
  assign t_r37_c56_9 = t_r37_c56_5 + t_r37_c56_6;
  assign t_r37_c56_10 = t_r37_c56_7 + t_r37_c56_8;
  assign t_r37_c56_11 = t_r37_c56_9 + t_r37_c56_10;
  assign t_r37_c56_12 = t_r37_c56_11 + p_38_57;
  assign out_37_56 = t_r37_c56_12 >> 4;

  assign t_r37_c57_0 = p_36_57 << 1;
  assign t_r37_c57_1 = p_37_56 << 1;
  assign t_r37_c57_2 = p_37_57 << 2;
  assign t_r37_c57_3 = p_37_58 << 1;
  assign t_r37_c57_4 = p_38_57 << 1;
  assign t_r37_c57_5 = t_r37_c57_0 + p_36_56;
  assign t_r37_c57_6 = t_r37_c57_1 + p_36_58;
  assign t_r37_c57_7 = t_r37_c57_2 + t_r37_c57_3;
  assign t_r37_c57_8 = t_r37_c57_4 + p_38_56;
  assign t_r37_c57_9 = t_r37_c57_5 + t_r37_c57_6;
  assign t_r37_c57_10 = t_r37_c57_7 + t_r37_c57_8;
  assign t_r37_c57_11 = t_r37_c57_9 + t_r37_c57_10;
  assign t_r37_c57_12 = t_r37_c57_11 + p_38_58;
  assign out_37_57 = t_r37_c57_12 >> 4;

  assign t_r37_c58_0 = p_36_58 << 1;
  assign t_r37_c58_1 = p_37_57 << 1;
  assign t_r37_c58_2 = p_37_58 << 2;
  assign t_r37_c58_3 = p_37_59 << 1;
  assign t_r37_c58_4 = p_38_58 << 1;
  assign t_r37_c58_5 = t_r37_c58_0 + p_36_57;
  assign t_r37_c58_6 = t_r37_c58_1 + p_36_59;
  assign t_r37_c58_7 = t_r37_c58_2 + t_r37_c58_3;
  assign t_r37_c58_8 = t_r37_c58_4 + p_38_57;
  assign t_r37_c58_9 = t_r37_c58_5 + t_r37_c58_6;
  assign t_r37_c58_10 = t_r37_c58_7 + t_r37_c58_8;
  assign t_r37_c58_11 = t_r37_c58_9 + t_r37_c58_10;
  assign t_r37_c58_12 = t_r37_c58_11 + p_38_59;
  assign out_37_58 = t_r37_c58_12 >> 4;

  assign t_r37_c59_0 = p_36_59 << 1;
  assign t_r37_c59_1 = p_37_58 << 1;
  assign t_r37_c59_2 = p_37_59 << 2;
  assign t_r37_c59_3 = p_37_60 << 1;
  assign t_r37_c59_4 = p_38_59 << 1;
  assign t_r37_c59_5 = t_r37_c59_0 + p_36_58;
  assign t_r37_c59_6 = t_r37_c59_1 + p_36_60;
  assign t_r37_c59_7 = t_r37_c59_2 + t_r37_c59_3;
  assign t_r37_c59_8 = t_r37_c59_4 + p_38_58;
  assign t_r37_c59_9 = t_r37_c59_5 + t_r37_c59_6;
  assign t_r37_c59_10 = t_r37_c59_7 + t_r37_c59_8;
  assign t_r37_c59_11 = t_r37_c59_9 + t_r37_c59_10;
  assign t_r37_c59_12 = t_r37_c59_11 + p_38_60;
  assign out_37_59 = t_r37_c59_12 >> 4;

  assign t_r37_c60_0 = p_36_60 << 1;
  assign t_r37_c60_1 = p_37_59 << 1;
  assign t_r37_c60_2 = p_37_60 << 2;
  assign t_r37_c60_3 = p_37_61 << 1;
  assign t_r37_c60_4 = p_38_60 << 1;
  assign t_r37_c60_5 = t_r37_c60_0 + p_36_59;
  assign t_r37_c60_6 = t_r37_c60_1 + p_36_61;
  assign t_r37_c60_7 = t_r37_c60_2 + t_r37_c60_3;
  assign t_r37_c60_8 = t_r37_c60_4 + p_38_59;
  assign t_r37_c60_9 = t_r37_c60_5 + t_r37_c60_6;
  assign t_r37_c60_10 = t_r37_c60_7 + t_r37_c60_8;
  assign t_r37_c60_11 = t_r37_c60_9 + t_r37_c60_10;
  assign t_r37_c60_12 = t_r37_c60_11 + p_38_61;
  assign out_37_60 = t_r37_c60_12 >> 4;

  assign t_r37_c61_0 = p_36_61 << 1;
  assign t_r37_c61_1 = p_37_60 << 1;
  assign t_r37_c61_2 = p_37_61 << 2;
  assign t_r37_c61_3 = p_37_62 << 1;
  assign t_r37_c61_4 = p_38_61 << 1;
  assign t_r37_c61_5 = t_r37_c61_0 + p_36_60;
  assign t_r37_c61_6 = t_r37_c61_1 + p_36_62;
  assign t_r37_c61_7 = t_r37_c61_2 + t_r37_c61_3;
  assign t_r37_c61_8 = t_r37_c61_4 + p_38_60;
  assign t_r37_c61_9 = t_r37_c61_5 + t_r37_c61_6;
  assign t_r37_c61_10 = t_r37_c61_7 + t_r37_c61_8;
  assign t_r37_c61_11 = t_r37_c61_9 + t_r37_c61_10;
  assign t_r37_c61_12 = t_r37_c61_11 + p_38_62;
  assign out_37_61 = t_r37_c61_12 >> 4;

  assign t_r37_c62_0 = p_36_62 << 1;
  assign t_r37_c62_1 = p_37_61 << 1;
  assign t_r37_c62_2 = p_37_62 << 2;
  assign t_r37_c62_3 = p_37_63 << 1;
  assign t_r37_c62_4 = p_38_62 << 1;
  assign t_r37_c62_5 = t_r37_c62_0 + p_36_61;
  assign t_r37_c62_6 = t_r37_c62_1 + p_36_63;
  assign t_r37_c62_7 = t_r37_c62_2 + t_r37_c62_3;
  assign t_r37_c62_8 = t_r37_c62_4 + p_38_61;
  assign t_r37_c62_9 = t_r37_c62_5 + t_r37_c62_6;
  assign t_r37_c62_10 = t_r37_c62_7 + t_r37_c62_8;
  assign t_r37_c62_11 = t_r37_c62_9 + t_r37_c62_10;
  assign t_r37_c62_12 = t_r37_c62_11 + p_38_63;
  assign out_37_62 = t_r37_c62_12 >> 4;

  assign t_r37_c63_0 = p_36_63 << 1;
  assign t_r37_c63_1 = p_37_62 << 1;
  assign t_r37_c63_2 = p_37_63 << 2;
  assign t_r37_c63_3 = p_37_64 << 1;
  assign t_r37_c63_4 = p_38_63 << 1;
  assign t_r37_c63_5 = t_r37_c63_0 + p_36_62;
  assign t_r37_c63_6 = t_r37_c63_1 + p_36_64;
  assign t_r37_c63_7 = t_r37_c63_2 + t_r37_c63_3;
  assign t_r37_c63_8 = t_r37_c63_4 + p_38_62;
  assign t_r37_c63_9 = t_r37_c63_5 + t_r37_c63_6;
  assign t_r37_c63_10 = t_r37_c63_7 + t_r37_c63_8;
  assign t_r37_c63_11 = t_r37_c63_9 + t_r37_c63_10;
  assign t_r37_c63_12 = t_r37_c63_11 + p_38_64;
  assign out_37_63 = t_r37_c63_12 >> 4;

  assign t_r37_c64_0 = p_36_64 << 1;
  assign t_r37_c64_1 = p_37_63 << 1;
  assign t_r37_c64_2 = p_37_64 << 2;
  assign t_r37_c64_3 = p_37_65 << 1;
  assign t_r37_c64_4 = p_38_64 << 1;
  assign t_r37_c64_5 = t_r37_c64_0 + p_36_63;
  assign t_r37_c64_6 = t_r37_c64_1 + p_36_65;
  assign t_r37_c64_7 = t_r37_c64_2 + t_r37_c64_3;
  assign t_r37_c64_8 = t_r37_c64_4 + p_38_63;
  assign t_r37_c64_9 = t_r37_c64_5 + t_r37_c64_6;
  assign t_r37_c64_10 = t_r37_c64_7 + t_r37_c64_8;
  assign t_r37_c64_11 = t_r37_c64_9 + t_r37_c64_10;
  assign t_r37_c64_12 = t_r37_c64_11 + p_38_65;
  assign out_37_64 = t_r37_c64_12 >> 4;

  assign t_r38_c1_0 = p_37_1 << 1;
  assign t_r38_c1_1 = p_38_0 << 1;
  assign t_r38_c1_2 = p_38_1 << 2;
  assign t_r38_c1_3 = p_38_2 << 1;
  assign t_r38_c1_4 = p_39_1 << 1;
  assign t_r38_c1_5 = t_r38_c1_0 + p_37_0;
  assign t_r38_c1_6 = t_r38_c1_1 + p_37_2;
  assign t_r38_c1_7 = t_r38_c1_2 + t_r38_c1_3;
  assign t_r38_c1_8 = t_r38_c1_4 + p_39_0;
  assign t_r38_c1_9 = t_r38_c1_5 + t_r38_c1_6;
  assign t_r38_c1_10 = t_r38_c1_7 + t_r38_c1_8;
  assign t_r38_c1_11 = t_r38_c1_9 + t_r38_c1_10;
  assign t_r38_c1_12 = t_r38_c1_11 + p_39_2;
  assign out_38_1 = t_r38_c1_12 >> 4;

  assign t_r38_c2_0 = p_37_2 << 1;
  assign t_r38_c2_1 = p_38_1 << 1;
  assign t_r38_c2_2 = p_38_2 << 2;
  assign t_r38_c2_3 = p_38_3 << 1;
  assign t_r38_c2_4 = p_39_2 << 1;
  assign t_r38_c2_5 = t_r38_c2_0 + p_37_1;
  assign t_r38_c2_6 = t_r38_c2_1 + p_37_3;
  assign t_r38_c2_7 = t_r38_c2_2 + t_r38_c2_3;
  assign t_r38_c2_8 = t_r38_c2_4 + p_39_1;
  assign t_r38_c2_9 = t_r38_c2_5 + t_r38_c2_6;
  assign t_r38_c2_10 = t_r38_c2_7 + t_r38_c2_8;
  assign t_r38_c2_11 = t_r38_c2_9 + t_r38_c2_10;
  assign t_r38_c2_12 = t_r38_c2_11 + p_39_3;
  assign out_38_2 = t_r38_c2_12 >> 4;

  assign t_r38_c3_0 = p_37_3 << 1;
  assign t_r38_c3_1 = p_38_2 << 1;
  assign t_r38_c3_2 = p_38_3 << 2;
  assign t_r38_c3_3 = p_38_4 << 1;
  assign t_r38_c3_4 = p_39_3 << 1;
  assign t_r38_c3_5 = t_r38_c3_0 + p_37_2;
  assign t_r38_c3_6 = t_r38_c3_1 + p_37_4;
  assign t_r38_c3_7 = t_r38_c3_2 + t_r38_c3_3;
  assign t_r38_c3_8 = t_r38_c3_4 + p_39_2;
  assign t_r38_c3_9 = t_r38_c3_5 + t_r38_c3_6;
  assign t_r38_c3_10 = t_r38_c3_7 + t_r38_c3_8;
  assign t_r38_c3_11 = t_r38_c3_9 + t_r38_c3_10;
  assign t_r38_c3_12 = t_r38_c3_11 + p_39_4;
  assign out_38_3 = t_r38_c3_12 >> 4;

  assign t_r38_c4_0 = p_37_4 << 1;
  assign t_r38_c4_1 = p_38_3 << 1;
  assign t_r38_c4_2 = p_38_4 << 2;
  assign t_r38_c4_3 = p_38_5 << 1;
  assign t_r38_c4_4 = p_39_4 << 1;
  assign t_r38_c4_5 = t_r38_c4_0 + p_37_3;
  assign t_r38_c4_6 = t_r38_c4_1 + p_37_5;
  assign t_r38_c4_7 = t_r38_c4_2 + t_r38_c4_3;
  assign t_r38_c4_8 = t_r38_c4_4 + p_39_3;
  assign t_r38_c4_9 = t_r38_c4_5 + t_r38_c4_6;
  assign t_r38_c4_10 = t_r38_c4_7 + t_r38_c4_8;
  assign t_r38_c4_11 = t_r38_c4_9 + t_r38_c4_10;
  assign t_r38_c4_12 = t_r38_c4_11 + p_39_5;
  assign out_38_4 = t_r38_c4_12 >> 4;

  assign t_r38_c5_0 = p_37_5 << 1;
  assign t_r38_c5_1 = p_38_4 << 1;
  assign t_r38_c5_2 = p_38_5 << 2;
  assign t_r38_c5_3 = p_38_6 << 1;
  assign t_r38_c5_4 = p_39_5 << 1;
  assign t_r38_c5_5 = t_r38_c5_0 + p_37_4;
  assign t_r38_c5_6 = t_r38_c5_1 + p_37_6;
  assign t_r38_c5_7 = t_r38_c5_2 + t_r38_c5_3;
  assign t_r38_c5_8 = t_r38_c5_4 + p_39_4;
  assign t_r38_c5_9 = t_r38_c5_5 + t_r38_c5_6;
  assign t_r38_c5_10 = t_r38_c5_7 + t_r38_c5_8;
  assign t_r38_c5_11 = t_r38_c5_9 + t_r38_c5_10;
  assign t_r38_c5_12 = t_r38_c5_11 + p_39_6;
  assign out_38_5 = t_r38_c5_12 >> 4;

  assign t_r38_c6_0 = p_37_6 << 1;
  assign t_r38_c6_1 = p_38_5 << 1;
  assign t_r38_c6_2 = p_38_6 << 2;
  assign t_r38_c6_3 = p_38_7 << 1;
  assign t_r38_c6_4 = p_39_6 << 1;
  assign t_r38_c6_5 = t_r38_c6_0 + p_37_5;
  assign t_r38_c6_6 = t_r38_c6_1 + p_37_7;
  assign t_r38_c6_7 = t_r38_c6_2 + t_r38_c6_3;
  assign t_r38_c6_8 = t_r38_c6_4 + p_39_5;
  assign t_r38_c6_9 = t_r38_c6_5 + t_r38_c6_6;
  assign t_r38_c6_10 = t_r38_c6_7 + t_r38_c6_8;
  assign t_r38_c6_11 = t_r38_c6_9 + t_r38_c6_10;
  assign t_r38_c6_12 = t_r38_c6_11 + p_39_7;
  assign out_38_6 = t_r38_c6_12 >> 4;

  assign t_r38_c7_0 = p_37_7 << 1;
  assign t_r38_c7_1 = p_38_6 << 1;
  assign t_r38_c7_2 = p_38_7 << 2;
  assign t_r38_c7_3 = p_38_8 << 1;
  assign t_r38_c7_4 = p_39_7 << 1;
  assign t_r38_c7_5 = t_r38_c7_0 + p_37_6;
  assign t_r38_c7_6 = t_r38_c7_1 + p_37_8;
  assign t_r38_c7_7 = t_r38_c7_2 + t_r38_c7_3;
  assign t_r38_c7_8 = t_r38_c7_4 + p_39_6;
  assign t_r38_c7_9 = t_r38_c7_5 + t_r38_c7_6;
  assign t_r38_c7_10 = t_r38_c7_7 + t_r38_c7_8;
  assign t_r38_c7_11 = t_r38_c7_9 + t_r38_c7_10;
  assign t_r38_c7_12 = t_r38_c7_11 + p_39_8;
  assign out_38_7 = t_r38_c7_12 >> 4;

  assign t_r38_c8_0 = p_37_8 << 1;
  assign t_r38_c8_1 = p_38_7 << 1;
  assign t_r38_c8_2 = p_38_8 << 2;
  assign t_r38_c8_3 = p_38_9 << 1;
  assign t_r38_c8_4 = p_39_8 << 1;
  assign t_r38_c8_5 = t_r38_c8_0 + p_37_7;
  assign t_r38_c8_6 = t_r38_c8_1 + p_37_9;
  assign t_r38_c8_7 = t_r38_c8_2 + t_r38_c8_3;
  assign t_r38_c8_8 = t_r38_c8_4 + p_39_7;
  assign t_r38_c8_9 = t_r38_c8_5 + t_r38_c8_6;
  assign t_r38_c8_10 = t_r38_c8_7 + t_r38_c8_8;
  assign t_r38_c8_11 = t_r38_c8_9 + t_r38_c8_10;
  assign t_r38_c8_12 = t_r38_c8_11 + p_39_9;
  assign out_38_8 = t_r38_c8_12 >> 4;

  assign t_r38_c9_0 = p_37_9 << 1;
  assign t_r38_c9_1 = p_38_8 << 1;
  assign t_r38_c9_2 = p_38_9 << 2;
  assign t_r38_c9_3 = p_38_10 << 1;
  assign t_r38_c9_4 = p_39_9 << 1;
  assign t_r38_c9_5 = t_r38_c9_0 + p_37_8;
  assign t_r38_c9_6 = t_r38_c9_1 + p_37_10;
  assign t_r38_c9_7 = t_r38_c9_2 + t_r38_c9_3;
  assign t_r38_c9_8 = t_r38_c9_4 + p_39_8;
  assign t_r38_c9_9 = t_r38_c9_5 + t_r38_c9_6;
  assign t_r38_c9_10 = t_r38_c9_7 + t_r38_c9_8;
  assign t_r38_c9_11 = t_r38_c9_9 + t_r38_c9_10;
  assign t_r38_c9_12 = t_r38_c9_11 + p_39_10;
  assign out_38_9 = t_r38_c9_12 >> 4;

  assign t_r38_c10_0 = p_37_10 << 1;
  assign t_r38_c10_1 = p_38_9 << 1;
  assign t_r38_c10_2 = p_38_10 << 2;
  assign t_r38_c10_3 = p_38_11 << 1;
  assign t_r38_c10_4 = p_39_10 << 1;
  assign t_r38_c10_5 = t_r38_c10_0 + p_37_9;
  assign t_r38_c10_6 = t_r38_c10_1 + p_37_11;
  assign t_r38_c10_7 = t_r38_c10_2 + t_r38_c10_3;
  assign t_r38_c10_8 = t_r38_c10_4 + p_39_9;
  assign t_r38_c10_9 = t_r38_c10_5 + t_r38_c10_6;
  assign t_r38_c10_10 = t_r38_c10_7 + t_r38_c10_8;
  assign t_r38_c10_11 = t_r38_c10_9 + t_r38_c10_10;
  assign t_r38_c10_12 = t_r38_c10_11 + p_39_11;
  assign out_38_10 = t_r38_c10_12 >> 4;

  assign t_r38_c11_0 = p_37_11 << 1;
  assign t_r38_c11_1 = p_38_10 << 1;
  assign t_r38_c11_2 = p_38_11 << 2;
  assign t_r38_c11_3 = p_38_12 << 1;
  assign t_r38_c11_4 = p_39_11 << 1;
  assign t_r38_c11_5 = t_r38_c11_0 + p_37_10;
  assign t_r38_c11_6 = t_r38_c11_1 + p_37_12;
  assign t_r38_c11_7 = t_r38_c11_2 + t_r38_c11_3;
  assign t_r38_c11_8 = t_r38_c11_4 + p_39_10;
  assign t_r38_c11_9 = t_r38_c11_5 + t_r38_c11_6;
  assign t_r38_c11_10 = t_r38_c11_7 + t_r38_c11_8;
  assign t_r38_c11_11 = t_r38_c11_9 + t_r38_c11_10;
  assign t_r38_c11_12 = t_r38_c11_11 + p_39_12;
  assign out_38_11 = t_r38_c11_12 >> 4;

  assign t_r38_c12_0 = p_37_12 << 1;
  assign t_r38_c12_1 = p_38_11 << 1;
  assign t_r38_c12_2 = p_38_12 << 2;
  assign t_r38_c12_3 = p_38_13 << 1;
  assign t_r38_c12_4 = p_39_12 << 1;
  assign t_r38_c12_5 = t_r38_c12_0 + p_37_11;
  assign t_r38_c12_6 = t_r38_c12_1 + p_37_13;
  assign t_r38_c12_7 = t_r38_c12_2 + t_r38_c12_3;
  assign t_r38_c12_8 = t_r38_c12_4 + p_39_11;
  assign t_r38_c12_9 = t_r38_c12_5 + t_r38_c12_6;
  assign t_r38_c12_10 = t_r38_c12_7 + t_r38_c12_8;
  assign t_r38_c12_11 = t_r38_c12_9 + t_r38_c12_10;
  assign t_r38_c12_12 = t_r38_c12_11 + p_39_13;
  assign out_38_12 = t_r38_c12_12 >> 4;

  assign t_r38_c13_0 = p_37_13 << 1;
  assign t_r38_c13_1 = p_38_12 << 1;
  assign t_r38_c13_2 = p_38_13 << 2;
  assign t_r38_c13_3 = p_38_14 << 1;
  assign t_r38_c13_4 = p_39_13 << 1;
  assign t_r38_c13_5 = t_r38_c13_0 + p_37_12;
  assign t_r38_c13_6 = t_r38_c13_1 + p_37_14;
  assign t_r38_c13_7 = t_r38_c13_2 + t_r38_c13_3;
  assign t_r38_c13_8 = t_r38_c13_4 + p_39_12;
  assign t_r38_c13_9 = t_r38_c13_5 + t_r38_c13_6;
  assign t_r38_c13_10 = t_r38_c13_7 + t_r38_c13_8;
  assign t_r38_c13_11 = t_r38_c13_9 + t_r38_c13_10;
  assign t_r38_c13_12 = t_r38_c13_11 + p_39_14;
  assign out_38_13 = t_r38_c13_12 >> 4;

  assign t_r38_c14_0 = p_37_14 << 1;
  assign t_r38_c14_1 = p_38_13 << 1;
  assign t_r38_c14_2 = p_38_14 << 2;
  assign t_r38_c14_3 = p_38_15 << 1;
  assign t_r38_c14_4 = p_39_14 << 1;
  assign t_r38_c14_5 = t_r38_c14_0 + p_37_13;
  assign t_r38_c14_6 = t_r38_c14_1 + p_37_15;
  assign t_r38_c14_7 = t_r38_c14_2 + t_r38_c14_3;
  assign t_r38_c14_8 = t_r38_c14_4 + p_39_13;
  assign t_r38_c14_9 = t_r38_c14_5 + t_r38_c14_6;
  assign t_r38_c14_10 = t_r38_c14_7 + t_r38_c14_8;
  assign t_r38_c14_11 = t_r38_c14_9 + t_r38_c14_10;
  assign t_r38_c14_12 = t_r38_c14_11 + p_39_15;
  assign out_38_14 = t_r38_c14_12 >> 4;

  assign t_r38_c15_0 = p_37_15 << 1;
  assign t_r38_c15_1 = p_38_14 << 1;
  assign t_r38_c15_2 = p_38_15 << 2;
  assign t_r38_c15_3 = p_38_16 << 1;
  assign t_r38_c15_4 = p_39_15 << 1;
  assign t_r38_c15_5 = t_r38_c15_0 + p_37_14;
  assign t_r38_c15_6 = t_r38_c15_1 + p_37_16;
  assign t_r38_c15_7 = t_r38_c15_2 + t_r38_c15_3;
  assign t_r38_c15_8 = t_r38_c15_4 + p_39_14;
  assign t_r38_c15_9 = t_r38_c15_5 + t_r38_c15_6;
  assign t_r38_c15_10 = t_r38_c15_7 + t_r38_c15_8;
  assign t_r38_c15_11 = t_r38_c15_9 + t_r38_c15_10;
  assign t_r38_c15_12 = t_r38_c15_11 + p_39_16;
  assign out_38_15 = t_r38_c15_12 >> 4;

  assign t_r38_c16_0 = p_37_16 << 1;
  assign t_r38_c16_1 = p_38_15 << 1;
  assign t_r38_c16_2 = p_38_16 << 2;
  assign t_r38_c16_3 = p_38_17 << 1;
  assign t_r38_c16_4 = p_39_16 << 1;
  assign t_r38_c16_5 = t_r38_c16_0 + p_37_15;
  assign t_r38_c16_6 = t_r38_c16_1 + p_37_17;
  assign t_r38_c16_7 = t_r38_c16_2 + t_r38_c16_3;
  assign t_r38_c16_8 = t_r38_c16_4 + p_39_15;
  assign t_r38_c16_9 = t_r38_c16_5 + t_r38_c16_6;
  assign t_r38_c16_10 = t_r38_c16_7 + t_r38_c16_8;
  assign t_r38_c16_11 = t_r38_c16_9 + t_r38_c16_10;
  assign t_r38_c16_12 = t_r38_c16_11 + p_39_17;
  assign out_38_16 = t_r38_c16_12 >> 4;

  assign t_r38_c17_0 = p_37_17 << 1;
  assign t_r38_c17_1 = p_38_16 << 1;
  assign t_r38_c17_2 = p_38_17 << 2;
  assign t_r38_c17_3 = p_38_18 << 1;
  assign t_r38_c17_4 = p_39_17 << 1;
  assign t_r38_c17_5 = t_r38_c17_0 + p_37_16;
  assign t_r38_c17_6 = t_r38_c17_1 + p_37_18;
  assign t_r38_c17_7 = t_r38_c17_2 + t_r38_c17_3;
  assign t_r38_c17_8 = t_r38_c17_4 + p_39_16;
  assign t_r38_c17_9 = t_r38_c17_5 + t_r38_c17_6;
  assign t_r38_c17_10 = t_r38_c17_7 + t_r38_c17_8;
  assign t_r38_c17_11 = t_r38_c17_9 + t_r38_c17_10;
  assign t_r38_c17_12 = t_r38_c17_11 + p_39_18;
  assign out_38_17 = t_r38_c17_12 >> 4;

  assign t_r38_c18_0 = p_37_18 << 1;
  assign t_r38_c18_1 = p_38_17 << 1;
  assign t_r38_c18_2 = p_38_18 << 2;
  assign t_r38_c18_3 = p_38_19 << 1;
  assign t_r38_c18_4 = p_39_18 << 1;
  assign t_r38_c18_5 = t_r38_c18_0 + p_37_17;
  assign t_r38_c18_6 = t_r38_c18_1 + p_37_19;
  assign t_r38_c18_7 = t_r38_c18_2 + t_r38_c18_3;
  assign t_r38_c18_8 = t_r38_c18_4 + p_39_17;
  assign t_r38_c18_9 = t_r38_c18_5 + t_r38_c18_6;
  assign t_r38_c18_10 = t_r38_c18_7 + t_r38_c18_8;
  assign t_r38_c18_11 = t_r38_c18_9 + t_r38_c18_10;
  assign t_r38_c18_12 = t_r38_c18_11 + p_39_19;
  assign out_38_18 = t_r38_c18_12 >> 4;

  assign t_r38_c19_0 = p_37_19 << 1;
  assign t_r38_c19_1 = p_38_18 << 1;
  assign t_r38_c19_2 = p_38_19 << 2;
  assign t_r38_c19_3 = p_38_20 << 1;
  assign t_r38_c19_4 = p_39_19 << 1;
  assign t_r38_c19_5 = t_r38_c19_0 + p_37_18;
  assign t_r38_c19_6 = t_r38_c19_1 + p_37_20;
  assign t_r38_c19_7 = t_r38_c19_2 + t_r38_c19_3;
  assign t_r38_c19_8 = t_r38_c19_4 + p_39_18;
  assign t_r38_c19_9 = t_r38_c19_5 + t_r38_c19_6;
  assign t_r38_c19_10 = t_r38_c19_7 + t_r38_c19_8;
  assign t_r38_c19_11 = t_r38_c19_9 + t_r38_c19_10;
  assign t_r38_c19_12 = t_r38_c19_11 + p_39_20;
  assign out_38_19 = t_r38_c19_12 >> 4;

  assign t_r38_c20_0 = p_37_20 << 1;
  assign t_r38_c20_1 = p_38_19 << 1;
  assign t_r38_c20_2 = p_38_20 << 2;
  assign t_r38_c20_3 = p_38_21 << 1;
  assign t_r38_c20_4 = p_39_20 << 1;
  assign t_r38_c20_5 = t_r38_c20_0 + p_37_19;
  assign t_r38_c20_6 = t_r38_c20_1 + p_37_21;
  assign t_r38_c20_7 = t_r38_c20_2 + t_r38_c20_3;
  assign t_r38_c20_8 = t_r38_c20_4 + p_39_19;
  assign t_r38_c20_9 = t_r38_c20_5 + t_r38_c20_6;
  assign t_r38_c20_10 = t_r38_c20_7 + t_r38_c20_8;
  assign t_r38_c20_11 = t_r38_c20_9 + t_r38_c20_10;
  assign t_r38_c20_12 = t_r38_c20_11 + p_39_21;
  assign out_38_20 = t_r38_c20_12 >> 4;

  assign t_r38_c21_0 = p_37_21 << 1;
  assign t_r38_c21_1 = p_38_20 << 1;
  assign t_r38_c21_2 = p_38_21 << 2;
  assign t_r38_c21_3 = p_38_22 << 1;
  assign t_r38_c21_4 = p_39_21 << 1;
  assign t_r38_c21_5 = t_r38_c21_0 + p_37_20;
  assign t_r38_c21_6 = t_r38_c21_1 + p_37_22;
  assign t_r38_c21_7 = t_r38_c21_2 + t_r38_c21_3;
  assign t_r38_c21_8 = t_r38_c21_4 + p_39_20;
  assign t_r38_c21_9 = t_r38_c21_5 + t_r38_c21_6;
  assign t_r38_c21_10 = t_r38_c21_7 + t_r38_c21_8;
  assign t_r38_c21_11 = t_r38_c21_9 + t_r38_c21_10;
  assign t_r38_c21_12 = t_r38_c21_11 + p_39_22;
  assign out_38_21 = t_r38_c21_12 >> 4;

  assign t_r38_c22_0 = p_37_22 << 1;
  assign t_r38_c22_1 = p_38_21 << 1;
  assign t_r38_c22_2 = p_38_22 << 2;
  assign t_r38_c22_3 = p_38_23 << 1;
  assign t_r38_c22_4 = p_39_22 << 1;
  assign t_r38_c22_5 = t_r38_c22_0 + p_37_21;
  assign t_r38_c22_6 = t_r38_c22_1 + p_37_23;
  assign t_r38_c22_7 = t_r38_c22_2 + t_r38_c22_3;
  assign t_r38_c22_8 = t_r38_c22_4 + p_39_21;
  assign t_r38_c22_9 = t_r38_c22_5 + t_r38_c22_6;
  assign t_r38_c22_10 = t_r38_c22_7 + t_r38_c22_8;
  assign t_r38_c22_11 = t_r38_c22_9 + t_r38_c22_10;
  assign t_r38_c22_12 = t_r38_c22_11 + p_39_23;
  assign out_38_22 = t_r38_c22_12 >> 4;

  assign t_r38_c23_0 = p_37_23 << 1;
  assign t_r38_c23_1 = p_38_22 << 1;
  assign t_r38_c23_2 = p_38_23 << 2;
  assign t_r38_c23_3 = p_38_24 << 1;
  assign t_r38_c23_4 = p_39_23 << 1;
  assign t_r38_c23_5 = t_r38_c23_0 + p_37_22;
  assign t_r38_c23_6 = t_r38_c23_1 + p_37_24;
  assign t_r38_c23_7 = t_r38_c23_2 + t_r38_c23_3;
  assign t_r38_c23_8 = t_r38_c23_4 + p_39_22;
  assign t_r38_c23_9 = t_r38_c23_5 + t_r38_c23_6;
  assign t_r38_c23_10 = t_r38_c23_7 + t_r38_c23_8;
  assign t_r38_c23_11 = t_r38_c23_9 + t_r38_c23_10;
  assign t_r38_c23_12 = t_r38_c23_11 + p_39_24;
  assign out_38_23 = t_r38_c23_12 >> 4;

  assign t_r38_c24_0 = p_37_24 << 1;
  assign t_r38_c24_1 = p_38_23 << 1;
  assign t_r38_c24_2 = p_38_24 << 2;
  assign t_r38_c24_3 = p_38_25 << 1;
  assign t_r38_c24_4 = p_39_24 << 1;
  assign t_r38_c24_5 = t_r38_c24_0 + p_37_23;
  assign t_r38_c24_6 = t_r38_c24_1 + p_37_25;
  assign t_r38_c24_7 = t_r38_c24_2 + t_r38_c24_3;
  assign t_r38_c24_8 = t_r38_c24_4 + p_39_23;
  assign t_r38_c24_9 = t_r38_c24_5 + t_r38_c24_6;
  assign t_r38_c24_10 = t_r38_c24_7 + t_r38_c24_8;
  assign t_r38_c24_11 = t_r38_c24_9 + t_r38_c24_10;
  assign t_r38_c24_12 = t_r38_c24_11 + p_39_25;
  assign out_38_24 = t_r38_c24_12 >> 4;

  assign t_r38_c25_0 = p_37_25 << 1;
  assign t_r38_c25_1 = p_38_24 << 1;
  assign t_r38_c25_2 = p_38_25 << 2;
  assign t_r38_c25_3 = p_38_26 << 1;
  assign t_r38_c25_4 = p_39_25 << 1;
  assign t_r38_c25_5 = t_r38_c25_0 + p_37_24;
  assign t_r38_c25_6 = t_r38_c25_1 + p_37_26;
  assign t_r38_c25_7 = t_r38_c25_2 + t_r38_c25_3;
  assign t_r38_c25_8 = t_r38_c25_4 + p_39_24;
  assign t_r38_c25_9 = t_r38_c25_5 + t_r38_c25_6;
  assign t_r38_c25_10 = t_r38_c25_7 + t_r38_c25_8;
  assign t_r38_c25_11 = t_r38_c25_9 + t_r38_c25_10;
  assign t_r38_c25_12 = t_r38_c25_11 + p_39_26;
  assign out_38_25 = t_r38_c25_12 >> 4;

  assign t_r38_c26_0 = p_37_26 << 1;
  assign t_r38_c26_1 = p_38_25 << 1;
  assign t_r38_c26_2 = p_38_26 << 2;
  assign t_r38_c26_3 = p_38_27 << 1;
  assign t_r38_c26_4 = p_39_26 << 1;
  assign t_r38_c26_5 = t_r38_c26_0 + p_37_25;
  assign t_r38_c26_6 = t_r38_c26_1 + p_37_27;
  assign t_r38_c26_7 = t_r38_c26_2 + t_r38_c26_3;
  assign t_r38_c26_8 = t_r38_c26_4 + p_39_25;
  assign t_r38_c26_9 = t_r38_c26_5 + t_r38_c26_6;
  assign t_r38_c26_10 = t_r38_c26_7 + t_r38_c26_8;
  assign t_r38_c26_11 = t_r38_c26_9 + t_r38_c26_10;
  assign t_r38_c26_12 = t_r38_c26_11 + p_39_27;
  assign out_38_26 = t_r38_c26_12 >> 4;

  assign t_r38_c27_0 = p_37_27 << 1;
  assign t_r38_c27_1 = p_38_26 << 1;
  assign t_r38_c27_2 = p_38_27 << 2;
  assign t_r38_c27_3 = p_38_28 << 1;
  assign t_r38_c27_4 = p_39_27 << 1;
  assign t_r38_c27_5 = t_r38_c27_0 + p_37_26;
  assign t_r38_c27_6 = t_r38_c27_1 + p_37_28;
  assign t_r38_c27_7 = t_r38_c27_2 + t_r38_c27_3;
  assign t_r38_c27_8 = t_r38_c27_4 + p_39_26;
  assign t_r38_c27_9 = t_r38_c27_5 + t_r38_c27_6;
  assign t_r38_c27_10 = t_r38_c27_7 + t_r38_c27_8;
  assign t_r38_c27_11 = t_r38_c27_9 + t_r38_c27_10;
  assign t_r38_c27_12 = t_r38_c27_11 + p_39_28;
  assign out_38_27 = t_r38_c27_12 >> 4;

  assign t_r38_c28_0 = p_37_28 << 1;
  assign t_r38_c28_1 = p_38_27 << 1;
  assign t_r38_c28_2 = p_38_28 << 2;
  assign t_r38_c28_3 = p_38_29 << 1;
  assign t_r38_c28_4 = p_39_28 << 1;
  assign t_r38_c28_5 = t_r38_c28_0 + p_37_27;
  assign t_r38_c28_6 = t_r38_c28_1 + p_37_29;
  assign t_r38_c28_7 = t_r38_c28_2 + t_r38_c28_3;
  assign t_r38_c28_8 = t_r38_c28_4 + p_39_27;
  assign t_r38_c28_9 = t_r38_c28_5 + t_r38_c28_6;
  assign t_r38_c28_10 = t_r38_c28_7 + t_r38_c28_8;
  assign t_r38_c28_11 = t_r38_c28_9 + t_r38_c28_10;
  assign t_r38_c28_12 = t_r38_c28_11 + p_39_29;
  assign out_38_28 = t_r38_c28_12 >> 4;

  assign t_r38_c29_0 = p_37_29 << 1;
  assign t_r38_c29_1 = p_38_28 << 1;
  assign t_r38_c29_2 = p_38_29 << 2;
  assign t_r38_c29_3 = p_38_30 << 1;
  assign t_r38_c29_4 = p_39_29 << 1;
  assign t_r38_c29_5 = t_r38_c29_0 + p_37_28;
  assign t_r38_c29_6 = t_r38_c29_1 + p_37_30;
  assign t_r38_c29_7 = t_r38_c29_2 + t_r38_c29_3;
  assign t_r38_c29_8 = t_r38_c29_4 + p_39_28;
  assign t_r38_c29_9 = t_r38_c29_5 + t_r38_c29_6;
  assign t_r38_c29_10 = t_r38_c29_7 + t_r38_c29_8;
  assign t_r38_c29_11 = t_r38_c29_9 + t_r38_c29_10;
  assign t_r38_c29_12 = t_r38_c29_11 + p_39_30;
  assign out_38_29 = t_r38_c29_12 >> 4;

  assign t_r38_c30_0 = p_37_30 << 1;
  assign t_r38_c30_1 = p_38_29 << 1;
  assign t_r38_c30_2 = p_38_30 << 2;
  assign t_r38_c30_3 = p_38_31 << 1;
  assign t_r38_c30_4 = p_39_30 << 1;
  assign t_r38_c30_5 = t_r38_c30_0 + p_37_29;
  assign t_r38_c30_6 = t_r38_c30_1 + p_37_31;
  assign t_r38_c30_7 = t_r38_c30_2 + t_r38_c30_3;
  assign t_r38_c30_8 = t_r38_c30_4 + p_39_29;
  assign t_r38_c30_9 = t_r38_c30_5 + t_r38_c30_6;
  assign t_r38_c30_10 = t_r38_c30_7 + t_r38_c30_8;
  assign t_r38_c30_11 = t_r38_c30_9 + t_r38_c30_10;
  assign t_r38_c30_12 = t_r38_c30_11 + p_39_31;
  assign out_38_30 = t_r38_c30_12 >> 4;

  assign t_r38_c31_0 = p_37_31 << 1;
  assign t_r38_c31_1 = p_38_30 << 1;
  assign t_r38_c31_2 = p_38_31 << 2;
  assign t_r38_c31_3 = p_38_32 << 1;
  assign t_r38_c31_4 = p_39_31 << 1;
  assign t_r38_c31_5 = t_r38_c31_0 + p_37_30;
  assign t_r38_c31_6 = t_r38_c31_1 + p_37_32;
  assign t_r38_c31_7 = t_r38_c31_2 + t_r38_c31_3;
  assign t_r38_c31_8 = t_r38_c31_4 + p_39_30;
  assign t_r38_c31_9 = t_r38_c31_5 + t_r38_c31_6;
  assign t_r38_c31_10 = t_r38_c31_7 + t_r38_c31_8;
  assign t_r38_c31_11 = t_r38_c31_9 + t_r38_c31_10;
  assign t_r38_c31_12 = t_r38_c31_11 + p_39_32;
  assign out_38_31 = t_r38_c31_12 >> 4;

  assign t_r38_c32_0 = p_37_32 << 1;
  assign t_r38_c32_1 = p_38_31 << 1;
  assign t_r38_c32_2 = p_38_32 << 2;
  assign t_r38_c32_3 = p_38_33 << 1;
  assign t_r38_c32_4 = p_39_32 << 1;
  assign t_r38_c32_5 = t_r38_c32_0 + p_37_31;
  assign t_r38_c32_6 = t_r38_c32_1 + p_37_33;
  assign t_r38_c32_7 = t_r38_c32_2 + t_r38_c32_3;
  assign t_r38_c32_8 = t_r38_c32_4 + p_39_31;
  assign t_r38_c32_9 = t_r38_c32_5 + t_r38_c32_6;
  assign t_r38_c32_10 = t_r38_c32_7 + t_r38_c32_8;
  assign t_r38_c32_11 = t_r38_c32_9 + t_r38_c32_10;
  assign t_r38_c32_12 = t_r38_c32_11 + p_39_33;
  assign out_38_32 = t_r38_c32_12 >> 4;

  assign t_r38_c33_0 = p_37_33 << 1;
  assign t_r38_c33_1 = p_38_32 << 1;
  assign t_r38_c33_2 = p_38_33 << 2;
  assign t_r38_c33_3 = p_38_34 << 1;
  assign t_r38_c33_4 = p_39_33 << 1;
  assign t_r38_c33_5 = t_r38_c33_0 + p_37_32;
  assign t_r38_c33_6 = t_r38_c33_1 + p_37_34;
  assign t_r38_c33_7 = t_r38_c33_2 + t_r38_c33_3;
  assign t_r38_c33_8 = t_r38_c33_4 + p_39_32;
  assign t_r38_c33_9 = t_r38_c33_5 + t_r38_c33_6;
  assign t_r38_c33_10 = t_r38_c33_7 + t_r38_c33_8;
  assign t_r38_c33_11 = t_r38_c33_9 + t_r38_c33_10;
  assign t_r38_c33_12 = t_r38_c33_11 + p_39_34;
  assign out_38_33 = t_r38_c33_12 >> 4;

  assign t_r38_c34_0 = p_37_34 << 1;
  assign t_r38_c34_1 = p_38_33 << 1;
  assign t_r38_c34_2 = p_38_34 << 2;
  assign t_r38_c34_3 = p_38_35 << 1;
  assign t_r38_c34_4 = p_39_34 << 1;
  assign t_r38_c34_5 = t_r38_c34_0 + p_37_33;
  assign t_r38_c34_6 = t_r38_c34_1 + p_37_35;
  assign t_r38_c34_7 = t_r38_c34_2 + t_r38_c34_3;
  assign t_r38_c34_8 = t_r38_c34_4 + p_39_33;
  assign t_r38_c34_9 = t_r38_c34_5 + t_r38_c34_6;
  assign t_r38_c34_10 = t_r38_c34_7 + t_r38_c34_8;
  assign t_r38_c34_11 = t_r38_c34_9 + t_r38_c34_10;
  assign t_r38_c34_12 = t_r38_c34_11 + p_39_35;
  assign out_38_34 = t_r38_c34_12 >> 4;

  assign t_r38_c35_0 = p_37_35 << 1;
  assign t_r38_c35_1 = p_38_34 << 1;
  assign t_r38_c35_2 = p_38_35 << 2;
  assign t_r38_c35_3 = p_38_36 << 1;
  assign t_r38_c35_4 = p_39_35 << 1;
  assign t_r38_c35_5 = t_r38_c35_0 + p_37_34;
  assign t_r38_c35_6 = t_r38_c35_1 + p_37_36;
  assign t_r38_c35_7 = t_r38_c35_2 + t_r38_c35_3;
  assign t_r38_c35_8 = t_r38_c35_4 + p_39_34;
  assign t_r38_c35_9 = t_r38_c35_5 + t_r38_c35_6;
  assign t_r38_c35_10 = t_r38_c35_7 + t_r38_c35_8;
  assign t_r38_c35_11 = t_r38_c35_9 + t_r38_c35_10;
  assign t_r38_c35_12 = t_r38_c35_11 + p_39_36;
  assign out_38_35 = t_r38_c35_12 >> 4;

  assign t_r38_c36_0 = p_37_36 << 1;
  assign t_r38_c36_1 = p_38_35 << 1;
  assign t_r38_c36_2 = p_38_36 << 2;
  assign t_r38_c36_3 = p_38_37 << 1;
  assign t_r38_c36_4 = p_39_36 << 1;
  assign t_r38_c36_5 = t_r38_c36_0 + p_37_35;
  assign t_r38_c36_6 = t_r38_c36_1 + p_37_37;
  assign t_r38_c36_7 = t_r38_c36_2 + t_r38_c36_3;
  assign t_r38_c36_8 = t_r38_c36_4 + p_39_35;
  assign t_r38_c36_9 = t_r38_c36_5 + t_r38_c36_6;
  assign t_r38_c36_10 = t_r38_c36_7 + t_r38_c36_8;
  assign t_r38_c36_11 = t_r38_c36_9 + t_r38_c36_10;
  assign t_r38_c36_12 = t_r38_c36_11 + p_39_37;
  assign out_38_36 = t_r38_c36_12 >> 4;

  assign t_r38_c37_0 = p_37_37 << 1;
  assign t_r38_c37_1 = p_38_36 << 1;
  assign t_r38_c37_2 = p_38_37 << 2;
  assign t_r38_c37_3 = p_38_38 << 1;
  assign t_r38_c37_4 = p_39_37 << 1;
  assign t_r38_c37_5 = t_r38_c37_0 + p_37_36;
  assign t_r38_c37_6 = t_r38_c37_1 + p_37_38;
  assign t_r38_c37_7 = t_r38_c37_2 + t_r38_c37_3;
  assign t_r38_c37_8 = t_r38_c37_4 + p_39_36;
  assign t_r38_c37_9 = t_r38_c37_5 + t_r38_c37_6;
  assign t_r38_c37_10 = t_r38_c37_7 + t_r38_c37_8;
  assign t_r38_c37_11 = t_r38_c37_9 + t_r38_c37_10;
  assign t_r38_c37_12 = t_r38_c37_11 + p_39_38;
  assign out_38_37 = t_r38_c37_12 >> 4;

  assign t_r38_c38_0 = p_37_38 << 1;
  assign t_r38_c38_1 = p_38_37 << 1;
  assign t_r38_c38_2 = p_38_38 << 2;
  assign t_r38_c38_3 = p_38_39 << 1;
  assign t_r38_c38_4 = p_39_38 << 1;
  assign t_r38_c38_5 = t_r38_c38_0 + p_37_37;
  assign t_r38_c38_6 = t_r38_c38_1 + p_37_39;
  assign t_r38_c38_7 = t_r38_c38_2 + t_r38_c38_3;
  assign t_r38_c38_8 = t_r38_c38_4 + p_39_37;
  assign t_r38_c38_9 = t_r38_c38_5 + t_r38_c38_6;
  assign t_r38_c38_10 = t_r38_c38_7 + t_r38_c38_8;
  assign t_r38_c38_11 = t_r38_c38_9 + t_r38_c38_10;
  assign t_r38_c38_12 = t_r38_c38_11 + p_39_39;
  assign out_38_38 = t_r38_c38_12 >> 4;

  assign t_r38_c39_0 = p_37_39 << 1;
  assign t_r38_c39_1 = p_38_38 << 1;
  assign t_r38_c39_2 = p_38_39 << 2;
  assign t_r38_c39_3 = p_38_40 << 1;
  assign t_r38_c39_4 = p_39_39 << 1;
  assign t_r38_c39_5 = t_r38_c39_0 + p_37_38;
  assign t_r38_c39_6 = t_r38_c39_1 + p_37_40;
  assign t_r38_c39_7 = t_r38_c39_2 + t_r38_c39_3;
  assign t_r38_c39_8 = t_r38_c39_4 + p_39_38;
  assign t_r38_c39_9 = t_r38_c39_5 + t_r38_c39_6;
  assign t_r38_c39_10 = t_r38_c39_7 + t_r38_c39_8;
  assign t_r38_c39_11 = t_r38_c39_9 + t_r38_c39_10;
  assign t_r38_c39_12 = t_r38_c39_11 + p_39_40;
  assign out_38_39 = t_r38_c39_12 >> 4;

  assign t_r38_c40_0 = p_37_40 << 1;
  assign t_r38_c40_1 = p_38_39 << 1;
  assign t_r38_c40_2 = p_38_40 << 2;
  assign t_r38_c40_3 = p_38_41 << 1;
  assign t_r38_c40_4 = p_39_40 << 1;
  assign t_r38_c40_5 = t_r38_c40_0 + p_37_39;
  assign t_r38_c40_6 = t_r38_c40_1 + p_37_41;
  assign t_r38_c40_7 = t_r38_c40_2 + t_r38_c40_3;
  assign t_r38_c40_8 = t_r38_c40_4 + p_39_39;
  assign t_r38_c40_9 = t_r38_c40_5 + t_r38_c40_6;
  assign t_r38_c40_10 = t_r38_c40_7 + t_r38_c40_8;
  assign t_r38_c40_11 = t_r38_c40_9 + t_r38_c40_10;
  assign t_r38_c40_12 = t_r38_c40_11 + p_39_41;
  assign out_38_40 = t_r38_c40_12 >> 4;

  assign t_r38_c41_0 = p_37_41 << 1;
  assign t_r38_c41_1 = p_38_40 << 1;
  assign t_r38_c41_2 = p_38_41 << 2;
  assign t_r38_c41_3 = p_38_42 << 1;
  assign t_r38_c41_4 = p_39_41 << 1;
  assign t_r38_c41_5 = t_r38_c41_0 + p_37_40;
  assign t_r38_c41_6 = t_r38_c41_1 + p_37_42;
  assign t_r38_c41_7 = t_r38_c41_2 + t_r38_c41_3;
  assign t_r38_c41_8 = t_r38_c41_4 + p_39_40;
  assign t_r38_c41_9 = t_r38_c41_5 + t_r38_c41_6;
  assign t_r38_c41_10 = t_r38_c41_7 + t_r38_c41_8;
  assign t_r38_c41_11 = t_r38_c41_9 + t_r38_c41_10;
  assign t_r38_c41_12 = t_r38_c41_11 + p_39_42;
  assign out_38_41 = t_r38_c41_12 >> 4;

  assign t_r38_c42_0 = p_37_42 << 1;
  assign t_r38_c42_1 = p_38_41 << 1;
  assign t_r38_c42_2 = p_38_42 << 2;
  assign t_r38_c42_3 = p_38_43 << 1;
  assign t_r38_c42_4 = p_39_42 << 1;
  assign t_r38_c42_5 = t_r38_c42_0 + p_37_41;
  assign t_r38_c42_6 = t_r38_c42_1 + p_37_43;
  assign t_r38_c42_7 = t_r38_c42_2 + t_r38_c42_3;
  assign t_r38_c42_8 = t_r38_c42_4 + p_39_41;
  assign t_r38_c42_9 = t_r38_c42_5 + t_r38_c42_6;
  assign t_r38_c42_10 = t_r38_c42_7 + t_r38_c42_8;
  assign t_r38_c42_11 = t_r38_c42_9 + t_r38_c42_10;
  assign t_r38_c42_12 = t_r38_c42_11 + p_39_43;
  assign out_38_42 = t_r38_c42_12 >> 4;

  assign t_r38_c43_0 = p_37_43 << 1;
  assign t_r38_c43_1 = p_38_42 << 1;
  assign t_r38_c43_2 = p_38_43 << 2;
  assign t_r38_c43_3 = p_38_44 << 1;
  assign t_r38_c43_4 = p_39_43 << 1;
  assign t_r38_c43_5 = t_r38_c43_0 + p_37_42;
  assign t_r38_c43_6 = t_r38_c43_1 + p_37_44;
  assign t_r38_c43_7 = t_r38_c43_2 + t_r38_c43_3;
  assign t_r38_c43_8 = t_r38_c43_4 + p_39_42;
  assign t_r38_c43_9 = t_r38_c43_5 + t_r38_c43_6;
  assign t_r38_c43_10 = t_r38_c43_7 + t_r38_c43_8;
  assign t_r38_c43_11 = t_r38_c43_9 + t_r38_c43_10;
  assign t_r38_c43_12 = t_r38_c43_11 + p_39_44;
  assign out_38_43 = t_r38_c43_12 >> 4;

  assign t_r38_c44_0 = p_37_44 << 1;
  assign t_r38_c44_1 = p_38_43 << 1;
  assign t_r38_c44_2 = p_38_44 << 2;
  assign t_r38_c44_3 = p_38_45 << 1;
  assign t_r38_c44_4 = p_39_44 << 1;
  assign t_r38_c44_5 = t_r38_c44_0 + p_37_43;
  assign t_r38_c44_6 = t_r38_c44_1 + p_37_45;
  assign t_r38_c44_7 = t_r38_c44_2 + t_r38_c44_3;
  assign t_r38_c44_8 = t_r38_c44_4 + p_39_43;
  assign t_r38_c44_9 = t_r38_c44_5 + t_r38_c44_6;
  assign t_r38_c44_10 = t_r38_c44_7 + t_r38_c44_8;
  assign t_r38_c44_11 = t_r38_c44_9 + t_r38_c44_10;
  assign t_r38_c44_12 = t_r38_c44_11 + p_39_45;
  assign out_38_44 = t_r38_c44_12 >> 4;

  assign t_r38_c45_0 = p_37_45 << 1;
  assign t_r38_c45_1 = p_38_44 << 1;
  assign t_r38_c45_2 = p_38_45 << 2;
  assign t_r38_c45_3 = p_38_46 << 1;
  assign t_r38_c45_4 = p_39_45 << 1;
  assign t_r38_c45_5 = t_r38_c45_0 + p_37_44;
  assign t_r38_c45_6 = t_r38_c45_1 + p_37_46;
  assign t_r38_c45_7 = t_r38_c45_2 + t_r38_c45_3;
  assign t_r38_c45_8 = t_r38_c45_4 + p_39_44;
  assign t_r38_c45_9 = t_r38_c45_5 + t_r38_c45_6;
  assign t_r38_c45_10 = t_r38_c45_7 + t_r38_c45_8;
  assign t_r38_c45_11 = t_r38_c45_9 + t_r38_c45_10;
  assign t_r38_c45_12 = t_r38_c45_11 + p_39_46;
  assign out_38_45 = t_r38_c45_12 >> 4;

  assign t_r38_c46_0 = p_37_46 << 1;
  assign t_r38_c46_1 = p_38_45 << 1;
  assign t_r38_c46_2 = p_38_46 << 2;
  assign t_r38_c46_3 = p_38_47 << 1;
  assign t_r38_c46_4 = p_39_46 << 1;
  assign t_r38_c46_5 = t_r38_c46_0 + p_37_45;
  assign t_r38_c46_6 = t_r38_c46_1 + p_37_47;
  assign t_r38_c46_7 = t_r38_c46_2 + t_r38_c46_3;
  assign t_r38_c46_8 = t_r38_c46_4 + p_39_45;
  assign t_r38_c46_9 = t_r38_c46_5 + t_r38_c46_6;
  assign t_r38_c46_10 = t_r38_c46_7 + t_r38_c46_8;
  assign t_r38_c46_11 = t_r38_c46_9 + t_r38_c46_10;
  assign t_r38_c46_12 = t_r38_c46_11 + p_39_47;
  assign out_38_46 = t_r38_c46_12 >> 4;

  assign t_r38_c47_0 = p_37_47 << 1;
  assign t_r38_c47_1 = p_38_46 << 1;
  assign t_r38_c47_2 = p_38_47 << 2;
  assign t_r38_c47_3 = p_38_48 << 1;
  assign t_r38_c47_4 = p_39_47 << 1;
  assign t_r38_c47_5 = t_r38_c47_0 + p_37_46;
  assign t_r38_c47_6 = t_r38_c47_1 + p_37_48;
  assign t_r38_c47_7 = t_r38_c47_2 + t_r38_c47_3;
  assign t_r38_c47_8 = t_r38_c47_4 + p_39_46;
  assign t_r38_c47_9 = t_r38_c47_5 + t_r38_c47_6;
  assign t_r38_c47_10 = t_r38_c47_7 + t_r38_c47_8;
  assign t_r38_c47_11 = t_r38_c47_9 + t_r38_c47_10;
  assign t_r38_c47_12 = t_r38_c47_11 + p_39_48;
  assign out_38_47 = t_r38_c47_12 >> 4;

  assign t_r38_c48_0 = p_37_48 << 1;
  assign t_r38_c48_1 = p_38_47 << 1;
  assign t_r38_c48_2 = p_38_48 << 2;
  assign t_r38_c48_3 = p_38_49 << 1;
  assign t_r38_c48_4 = p_39_48 << 1;
  assign t_r38_c48_5 = t_r38_c48_0 + p_37_47;
  assign t_r38_c48_6 = t_r38_c48_1 + p_37_49;
  assign t_r38_c48_7 = t_r38_c48_2 + t_r38_c48_3;
  assign t_r38_c48_8 = t_r38_c48_4 + p_39_47;
  assign t_r38_c48_9 = t_r38_c48_5 + t_r38_c48_6;
  assign t_r38_c48_10 = t_r38_c48_7 + t_r38_c48_8;
  assign t_r38_c48_11 = t_r38_c48_9 + t_r38_c48_10;
  assign t_r38_c48_12 = t_r38_c48_11 + p_39_49;
  assign out_38_48 = t_r38_c48_12 >> 4;

  assign t_r38_c49_0 = p_37_49 << 1;
  assign t_r38_c49_1 = p_38_48 << 1;
  assign t_r38_c49_2 = p_38_49 << 2;
  assign t_r38_c49_3 = p_38_50 << 1;
  assign t_r38_c49_4 = p_39_49 << 1;
  assign t_r38_c49_5 = t_r38_c49_0 + p_37_48;
  assign t_r38_c49_6 = t_r38_c49_1 + p_37_50;
  assign t_r38_c49_7 = t_r38_c49_2 + t_r38_c49_3;
  assign t_r38_c49_8 = t_r38_c49_4 + p_39_48;
  assign t_r38_c49_9 = t_r38_c49_5 + t_r38_c49_6;
  assign t_r38_c49_10 = t_r38_c49_7 + t_r38_c49_8;
  assign t_r38_c49_11 = t_r38_c49_9 + t_r38_c49_10;
  assign t_r38_c49_12 = t_r38_c49_11 + p_39_50;
  assign out_38_49 = t_r38_c49_12 >> 4;

  assign t_r38_c50_0 = p_37_50 << 1;
  assign t_r38_c50_1 = p_38_49 << 1;
  assign t_r38_c50_2 = p_38_50 << 2;
  assign t_r38_c50_3 = p_38_51 << 1;
  assign t_r38_c50_4 = p_39_50 << 1;
  assign t_r38_c50_5 = t_r38_c50_0 + p_37_49;
  assign t_r38_c50_6 = t_r38_c50_1 + p_37_51;
  assign t_r38_c50_7 = t_r38_c50_2 + t_r38_c50_3;
  assign t_r38_c50_8 = t_r38_c50_4 + p_39_49;
  assign t_r38_c50_9 = t_r38_c50_5 + t_r38_c50_6;
  assign t_r38_c50_10 = t_r38_c50_7 + t_r38_c50_8;
  assign t_r38_c50_11 = t_r38_c50_9 + t_r38_c50_10;
  assign t_r38_c50_12 = t_r38_c50_11 + p_39_51;
  assign out_38_50 = t_r38_c50_12 >> 4;

  assign t_r38_c51_0 = p_37_51 << 1;
  assign t_r38_c51_1 = p_38_50 << 1;
  assign t_r38_c51_2 = p_38_51 << 2;
  assign t_r38_c51_3 = p_38_52 << 1;
  assign t_r38_c51_4 = p_39_51 << 1;
  assign t_r38_c51_5 = t_r38_c51_0 + p_37_50;
  assign t_r38_c51_6 = t_r38_c51_1 + p_37_52;
  assign t_r38_c51_7 = t_r38_c51_2 + t_r38_c51_3;
  assign t_r38_c51_8 = t_r38_c51_4 + p_39_50;
  assign t_r38_c51_9 = t_r38_c51_5 + t_r38_c51_6;
  assign t_r38_c51_10 = t_r38_c51_7 + t_r38_c51_8;
  assign t_r38_c51_11 = t_r38_c51_9 + t_r38_c51_10;
  assign t_r38_c51_12 = t_r38_c51_11 + p_39_52;
  assign out_38_51 = t_r38_c51_12 >> 4;

  assign t_r38_c52_0 = p_37_52 << 1;
  assign t_r38_c52_1 = p_38_51 << 1;
  assign t_r38_c52_2 = p_38_52 << 2;
  assign t_r38_c52_3 = p_38_53 << 1;
  assign t_r38_c52_4 = p_39_52 << 1;
  assign t_r38_c52_5 = t_r38_c52_0 + p_37_51;
  assign t_r38_c52_6 = t_r38_c52_1 + p_37_53;
  assign t_r38_c52_7 = t_r38_c52_2 + t_r38_c52_3;
  assign t_r38_c52_8 = t_r38_c52_4 + p_39_51;
  assign t_r38_c52_9 = t_r38_c52_5 + t_r38_c52_6;
  assign t_r38_c52_10 = t_r38_c52_7 + t_r38_c52_8;
  assign t_r38_c52_11 = t_r38_c52_9 + t_r38_c52_10;
  assign t_r38_c52_12 = t_r38_c52_11 + p_39_53;
  assign out_38_52 = t_r38_c52_12 >> 4;

  assign t_r38_c53_0 = p_37_53 << 1;
  assign t_r38_c53_1 = p_38_52 << 1;
  assign t_r38_c53_2 = p_38_53 << 2;
  assign t_r38_c53_3 = p_38_54 << 1;
  assign t_r38_c53_4 = p_39_53 << 1;
  assign t_r38_c53_5 = t_r38_c53_0 + p_37_52;
  assign t_r38_c53_6 = t_r38_c53_1 + p_37_54;
  assign t_r38_c53_7 = t_r38_c53_2 + t_r38_c53_3;
  assign t_r38_c53_8 = t_r38_c53_4 + p_39_52;
  assign t_r38_c53_9 = t_r38_c53_5 + t_r38_c53_6;
  assign t_r38_c53_10 = t_r38_c53_7 + t_r38_c53_8;
  assign t_r38_c53_11 = t_r38_c53_9 + t_r38_c53_10;
  assign t_r38_c53_12 = t_r38_c53_11 + p_39_54;
  assign out_38_53 = t_r38_c53_12 >> 4;

  assign t_r38_c54_0 = p_37_54 << 1;
  assign t_r38_c54_1 = p_38_53 << 1;
  assign t_r38_c54_2 = p_38_54 << 2;
  assign t_r38_c54_3 = p_38_55 << 1;
  assign t_r38_c54_4 = p_39_54 << 1;
  assign t_r38_c54_5 = t_r38_c54_0 + p_37_53;
  assign t_r38_c54_6 = t_r38_c54_1 + p_37_55;
  assign t_r38_c54_7 = t_r38_c54_2 + t_r38_c54_3;
  assign t_r38_c54_8 = t_r38_c54_4 + p_39_53;
  assign t_r38_c54_9 = t_r38_c54_5 + t_r38_c54_6;
  assign t_r38_c54_10 = t_r38_c54_7 + t_r38_c54_8;
  assign t_r38_c54_11 = t_r38_c54_9 + t_r38_c54_10;
  assign t_r38_c54_12 = t_r38_c54_11 + p_39_55;
  assign out_38_54 = t_r38_c54_12 >> 4;

  assign t_r38_c55_0 = p_37_55 << 1;
  assign t_r38_c55_1 = p_38_54 << 1;
  assign t_r38_c55_2 = p_38_55 << 2;
  assign t_r38_c55_3 = p_38_56 << 1;
  assign t_r38_c55_4 = p_39_55 << 1;
  assign t_r38_c55_5 = t_r38_c55_0 + p_37_54;
  assign t_r38_c55_6 = t_r38_c55_1 + p_37_56;
  assign t_r38_c55_7 = t_r38_c55_2 + t_r38_c55_3;
  assign t_r38_c55_8 = t_r38_c55_4 + p_39_54;
  assign t_r38_c55_9 = t_r38_c55_5 + t_r38_c55_6;
  assign t_r38_c55_10 = t_r38_c55_7 + t_r38_c55_8;
  assign t_r38_c55_11 = t_r38_c55_9 + t_r38_c55_10;
  assign t_r38_c55_12 = t_r38_c55_11 + p_39_56;
  assign out_38_55 = t_r38_c55_12 >> 4;

  assign t_r38_c56_0 = p_37_56 << 1;
  assign t_r38_c56_1 = p_38_55 << 1;
  assign t_r38_c56_2 = p_38_56 << 2;
  assign t_r38_c56_3 = p_38_57 << 1;
  assign t_r38_c56_4 = p_39_56 << 1;
  assign t_r38_c56_5 = t_r38_c56_0 + p_37_55;
  assign t_r38_c56_6 = t_r38_c56_1 + p_37_57;
  assign t_r38_c56_7 = t_r38_c56_2 + t_r38_c56_3;
  assign t_r38_c56_8 = t_r38_c56_4 + p_39_55;
  assign t_r38_c56_9 = t_r38_c56_5 + t_r38_c56_6;
  assign t_r38_c56_10 = t_r38_c56_7 + t_r38_c56_8;
  assign t_r38_c56_11 = t_r38_c56_9 + t_r38_c56_10;
  assign t_r38_c56_12 = t_r38_c56_11 + p_39_57;
  assign out_38_56 = t_r38_c56_12 >> 4;

  assign t_r38_c57_0 = p_37_57 << 1;
  assign t_r38_c57_1 = p_38_56 << 1;
  assign t_r38_c57_2 = p_38_57 << 2;
  assign t_r38_c57_3 = p_38_58 << 1;
  assign t_r38_c57_4 = p_39_57 << 1;
  assign t_r38_c57_5 = t_r38_c57_0 + p_37_56;
  assign t_r38_c57_6 = t_r38_c57_1 + p_37_58;
  assign t_r38_c57_7 = t_r38_c57_2 + t_r38_c57_3;
  assign t_r38_c57_8 = t_r38_c57_4 + p_39_56;
  assign t_r38_c57_9 = t_r38_c57_5 + t_r38_c57_6;
  assign t_r38_c57_10 = t_r38_c57_7 + t_r38_c57_8;
  assign t_r38_c57_11 = t_r38_c57_9 + t_r38_c57_10;
  assign t_r38_c57_12 = t_r38_c57_11 + p_39_58;
  assign out_38_57 = t_r38_c57_12 >> 4;

  assign t_r38_c58_0 = p_37_58 << 1;
  assign t_r38_c58_1 = p_38_57 << 1;
  assign t_r38_c58_2 = p_38_58 << 2;
  assign t_r38_c58_3 = p_38_59 << 1;
  assign t_r38_c58_4 = p_39_58 << 1;
  assign t_r38_c58_5 = t_r38_c58_0 + p_37_57;
  assign t_r38_c58_6 = t_r38_c58_1 + p_37_59;
  assign t_r38_c58_7 = t_r38_c58_2 + t_r38_c58_3;
  assign t_r38_c58_8 = t_r38_c58_4 + p_39_57;
  assign t_r38_c58_9 = t_r38_c58_5 + t_r38_c58_6;
  assign t_r38_c58_10 = t_r38_c58_7 + t_r38_c58_8;
  assign t_r38_c58_11 = t_r38_c58_9 + t_r38_c58_10;
  assign t_r38_c58_12 = t_r38_c58_11 + p_39_59;
  assign out_38_58 = t_r38_c58_12 >> 4;

  assign t_r38_c59_0 = p_37_59 << 1;
  assign t_r38_c59_1 = p_38_58 << 1;
  assign t_r38_c59_2 = p_38_59 << 2;
  assign t_r38_c59_3 = p_38_60 << 1;
  assign t_r38_c59_4 = p_39_59 << 1;
  assign t_r38_c59_5 = t_r38_c59_0 + p_37_58;
  assign t_r38_c59_6 = t_r38_c59_1 + p_37_60;
  assign t_r38_c59_7 = t_r38_c59_2 + t_r38_c59_3;
  assign t_r38_c59_8 = t_r38_c59_4 + p_39_58;
  assign t_r38_c59_9 = t_r38_c59_5 + t_r38_c59_6;
  assign t_r38_c59_10 = t_r38_c59_7 + t_r38_c59_8;
  assign t_r38_c59_11 = t_r38_c59_9 + t_r38_c59_10;
  assign t_r38_c59_12 = t_r38_c59_11 + p_39_60;
  assign out_38_59 = t_r38_c59_12 >> 4;

  assign t_r38_c60_0 = p_37_60 << 1;
  assign t_r38_c60_1 = p_38_59 << 1;
  assign t_r38_c60_2 = p_38_60 << 2;
  assign t_r38_c60_3 = p_38_61 << 1;
  assign t_r38_c60_4 = p_39_60 << 1;
  assign t_r38_c60_5 = t_r38_c60_0 + p_37_59;
  assign t_r38_c60_6 = t_r38_c60_1 + p_37_61;
  assign t_r38_c60_7 = t_r38_c60_2 + t_r38_c60_3;
  assign t_r38_c60_8 = t_r38_c60_4 + p_39_59;
  assign t_r38_c60_9 = t_r38_c60_5 + t_r38_c60_6;
  assign t_r38_c60_10 = t_r38_c60_7 + t_r38_c60_8;
  assign t_r38_c60_11 = t_r38_c60_9 + t_r38_c60_10;
  assign t_r38_c60_12 = t_r38_c60_11 + p_39_61;
  assign out_38_60 = t_r38_c60_12 >> 4;

  assign t_r38_c61_0 = p_37_61 << 1;
  assign t_r38_c61_1 = p_38_60 << 1;
  assign t_r38_c61_2 = p_38_61 << 2;
  assign t_r38_c61_3 = p_38_62 << 1;
  assign t_r38_c61_4 = p_39_61 << 1;
  assign t_r38_c61_5 = t_r38_c61_0 + p_37_60;
  assign t_r38_c61_6 = t_r38_c61_1 + p_37_62;
  assign t_r38_c61_7 = t_r38_c61_2 + t_r38_c61_3;
  assign t_r38_c61_8 = t_r38_c61_4 + p_39_60;
  assign t_r38_c61_9 = t_r38_c61_5 + t_r38_c61_6;
  assign t_r38_c61_10 = t_r38_c61_7 + t_r38_c61_8;
  assign t_r38_c61_11 = t_r38_c61_9 + t_r38_c61_10;
  assign t_r38_c61_12 = t_r38_c61_11 + p_39_62;
  assign out_38_61 = t_r38_c61_12 >> 4;

  assign t_r38_c62_0 = p_37_62 << 1;
  assign t_r38_c62_1 = p_38_61 << 1;
  assign t_r38_c62_2 = p_38_62 << 2;
  assign t_r38_c62_3 = p_38_63 << 1;
  assign t_r38_c62_4 = p_39_62 << 1;
  assign t_r38_c62_5 = t_r38_c62_0 + p_37_61;
  assign t_r38_c62_6 = t_r38_c62_1 + p_37_63;
  assign t_r38_c62_7 = t_r38_c62_2 + t_r38_c62_3;
  assign t_r38_c62_8 = t_r38_c62_4 + p_39_61;
  assign t_r38_c62_9 = t_r38_c62_5 + t_r38_c62_6;
  assign t_r38_c62_10 = t_r38_c62_7 + t_r38_c62_8;
  assign t_r38_c62_11 = t_r38_c62_9 + t_r38_c62_10;
  assign t_r38_c62_12 = t_r38_c62_11 + p_39_63;
  assign out_38_62 = t_r38_c62_12 >> 4;

  assign t_r38_c63_0 = p_37_63 << 1;
  assign t_r38_c63_1 = p_38_62 << 1;
  assign t_r38_c63_2 = p_38_63 << 2;
  assign t_r38_c63_3 = p_38_64 << 1;
  assign t_r38_c63_4 = p_39_63 << 1;
  assign t_r38_c63_5 = t_r38_c63_0 + p_37_62;
  assign t_r38_c63_6 = t_r38_c63_1 + p_37_64;
  assign t_r38_c63_7 = t_r38_c63_2 + t_r38_c63_3;
  assign t_r38_c63_8 = t_r38_c63_4 + p_39_62;
  assign t_r38_c63_9 = t_r38_c63_5 + t_r38_c63_6;
  assign t_r38_c63_10 = t_r38_c63_7 + t_r38_c63_8;
  assign t_r38_c63_11 = t_r38_c63_9 + t_r38_c63_10;
  assign t_r38_c63_12 = t_r38_c63_11 + p_39_64;
  assign out_38_63 = t_r38_c63_12 >> 4;

  assign t_r38_c64_0 = p_37_64 << 1;
  assign t_r38_c64_1 = p_38_63 << 1;
  assign t_r38_c64_2 = p_38_64 << 2;
  assign t_r38_c64_3 = p_38_65 << 1;
  assign t_r38_c64_4 = p_39_64 << 1;
  assign t_r38_c64_5 = t_r38_c64_0 + p_37_63;
  assign t_r38_c64_6 = t_r38_c64_1 + p_37_65;
  assign t_r38_c64_7 = t_r38_c64_2 + t_r38_c64_3;
  assign t_r38_c64_8 = t_r38_c64_4 + p_39_63;
  assign t_r38_c64_9 = t_r38_c64_5 + t_r38_c64_6;
  assign t_r38_c64_10 = t_r38_c64_7 + t_r38_c64_8;
  assign t_r38_c64_11 = t_r38_c64_9 + t_r38_c64_10;
  assign t_r38_c64_12 = t_r38_c64_11 + p_39_65;
  assign out_38_64 = t_r38_c64_12 >> 4;

  assign t_r39_c1_0 = p_38_1 << 1;
  assign t_r39_c1_1 = p_39_0 << 1;
  assign t_r39_c1_2 = p_39_1 << 2;
  assign t_r39_c1_3 = p_39_2 << 1;
  assign t_r39_c1_4 = p_40_1 << 1;
  assign t_r39_c1_5 = t_r39_c1_0 + p_38_0;
  assign t_r39_c1_6 = t_r39_c1_1 + p_38_2;
  assign t_r39_c1_7 = t_r39_c1_2 + t_r39_c1_3;
  assign t_r39_c1_8 = t_r39_c1_4 + p_40_0;
  assign t_r39_c1_9 = t_r39_c1_5 + t_r39_c1_6;
  assign t_r39_c1_10 = t_r39_c1_7 + t_r39_c1_8;
  assign t_r39_c1_11 = t_r39_c1_9 + t_r39_c1_10;
  assign t_r39_c1_12 = t_r39_c1_11 + p_40_2;
  assign out_39_1 = t_r39_c1_12 >> 4;

  assign t_r39_c2_0 = p_38_2 << 1;
  assign t_r39_c2_1 = p_39_1 << 1;
  assign t_r39_c2_2 = p_39_2 << 2;
  assign t_r39_c2_3 = p_39_3 << 1;
  assign t_r39_c2_4 = p_40_2 << 1;
  assign t_r39_c2_5 = t_r39_c2_0 + p_38_1;
  assign t_r39_c2_6 = t_r39_c2_1 + p_38_3;
  assign t_r39_c2_7 = t_r39_c2_2 + t_r39_c2_3;
  assign t_r39_c2_8 = t_r39_c2_4 + p_40_1;
  assign t_r39_c2_9 = t_r39_c2_5 + t_r39_c2_6;
  assign t_r39_c2_10 = t_r39_c2_7 + t_r39_c2_8;
  assign t_r39_c2_11 = t_r39_c2_9 + t_r39_c2_10;
  assign t_r39_c2_12 = t_r39_c2_11 + p_40_3;
  assign out_39_2 = t_r39_c2_12 >> 4;

  assign t_r39_c3_0 = p_38_3 << 1;
  assign t_r39_c3_1 = p_39_2 << 1;
  assign t_r39_c3_2 = p_39_3 << 2;
  assign t_r39_c3_3 = p_39_4 << 1;
  assign t_r39_c3_4 = p_40_3 << 1;
  assign t_r39_c3_5 = t_r39_c3_0 + p_38_2;
  assign t_r39_c3_6 = t_r39_c3_1 + p_38_4;
  assign t_r39_c3_7 = t_r39_c3_2 + t_r39_c3_3;
  assign t_r39_c3_8 = t_r39_c3_4 + p_40_2;
  assign t_r39_c3_9 = t_r39_c3_5 + t_r39_c3_6;
  assign t_r39_c3_10 = t_r39_c3_7 + t_r39_c3_8;
  assign t_r39_c3_11 = t_r39_c3_9 + t_r39_c3_10;
  assign t_r39_c3_12 = t_r39_c3_11 + p_40_4;
  assign out_39_3 = t_r39_c3_12 >> 4;

  assign t_r39_c4_0 = p_38_4 << 1;
  assign t_r39_c4_1 = p_39_3 << 1;
  assign t_r39_c4_2 = p_39_4 << 2;
  assign t_r39_c4_3 = p_39_5 << 1;
  assign t_r39_c4_4 = p_40_4 << 1;
  assign t_r39_c4_5 = t_r39_c4_0 + p_38_3;
  assign t_r39_c4_6 = t_r39_c4_1 + p_38_5;
  assign t_r39_c4_7 = t_r39_c4_2 + t_r39_c4_3;
  assign t_r39_c4_8 = t_r39_c4_4 + p_40_3;
  assign t_r39_c4_9 = t_r39_c4_5 + t_r39_c4_6;
  assign t_r39_c4_10 = t_r39_c4_7 + t_r39_c4_8;
  assign t_r39_c4_11 = t_r39_c4_9 + t_r39_c4_10;
  assign t_r39_c4_12 = t_r39_c4_11 + p_40_5;
  assign out_39_4 = t_r39_c4_12 >> 4;

  assign t_r39_c5_0 = p_38_5 << 1;
  assign t_r39_c5_1 = p_39_4 << 1;
  assign t_r39_c5_2 = p_39_5 << 2;
  assign t_r39_c5_3 = p_39_6 << 1;
  assign t_r39_c5_4 = p_40_5 << 1;
  assign t_r39_c5_5 = t_r39_c5_0 + p_38_4;
  assign t_r39_c5_6 = t_r39_c5_1 + p_38_6;
  assign t_r39_c5_7 = t_r39_c5_2 + t_r39_c5_3;
  assign t_r39_c5_8 = t_r39_c5_4 + p_40_4;
  assign t_r39_c5_9 = t_r39_c5_5 + t_r39_c5_6;
  assign t_r39_c5_10 = t_r39_c5_7 + t_r39_c5_8;
  assign t_r39_c5_11 = t_r39_c5_9 + t_r39_c5_10;
  assign t_r39_c5_12 = t_r39_c5_11 + p_40_6;
  assign out_39_5 = t_r39_c5_12 >> 4;

  assign t_r39_c6_0 = p_38_6 << 1;
  assign t_r39_c6_1 = p_39_5 << 1;
  assign t_r39_c6_2 = p_39_6 << 2;
  assign t_r39_c6_3 = p_39_7 << 1;
  assign t_r39_c6_4 = p_40_6 << 1;
  assign t_r39_c6_5 = t_r39_c6_0 + p_38_5;
  assign t_r39_c6_6 = t_r39_c6_1 + p_38_7;
  assign t_r39_c6_7 = t_r39_c6_2 + t_r39_c6_3;
  assign t_r39_c6_8 = t_r39_c6_4 + p_40_5;
  assign t_r39_c6_9 = t_r39_c6_5 + t_r39_c6_6;
  assign t_r39_c6_10 = t_r39_c6_7 + t_r39_c6_8;
  assign t_r39_c6_11 = t_r39_c6_9 + t_r39_c6_10;
  assign t_r39_c6_12 = t_r39_c6_11 + p_40_7;
  assign out_39_6 = t_r39_c6_12 >> 4;

  assign t_r39_c7_0 = p_38_7 << 1;
  assign t_r39_c7_1 = p_39_6 << 1;
  assign t_r39_c7_2 = p_39_7 << 2;
  assign t_r39_c7_3 = p_39_8 << 1;
  assign t_r39_c7_4 = p_40_7 << 1;
  assign t_r39_c7_5 = t_r39_c7_0 + p_38_6;
  assign t_r39_c7_6 = t_r39_c7_1 + p_38_8;
  assign t_r39_c7_7 = t_r39_c7_2 + t_r39_c7_3;
  assign t_r39_c7_8 = t_r39_c7_4 + p_40_6;
  assign t_r39_c7_9 = t_r39_c7_5 + t_r39_c7_6;
  assign t_r39_c7_10 = t_r39_c7_7 + t_r39_c7_8;
  assign t_r39_c7_11 = t_r39_c7_9 + t_r39_c7_10;
  assign t_r39_c7_12 = t_r39_c7_11 + p_40_8;
  assign out_39_7 = t_r39_c7_12 >> 4;

  assign t_r39_c8_0 = p_38_8 << 1;
  assign t_r39_c8_1 = p_39_7 << 1;
  assign t_r39_c8_2 = p_39_8 << 2;
  assign t_r39_c8_3 = p_39_9 << 1;
  assign t_r39_c8_4 = p_40_8 << 1;
  assign t_r39_c8_5 = t_r39_c8_0 + p_38_7;
  assign t_r39_c8_6 = t_r39_c8_1 + p_38_9;
  assign t_r39_c8_7 = t_r39_c8_2 + t_r39_c8_3;
  assign t_r39_c8_8 = t_r39_c8_4 + p_40_7;
  assign t_r39_c8_9 = t_r39_c8_5 + t_r39_c8_6;
  assign t_r39_c8_10 = t_r39_c8_7 + t_r39_c8_8;
  assign t_r39_c8_11 = t_r39_c8_9 + t_r39_c8_10;
  assign t_r39_c8_12 = t_r39_c8_11 + p_40_9;
  assign out_39_8 = t_r39_c8_12 >> 4;

  assign t_r39_c9_0 = p_38_9 << 1;
  assign t_r39_c9_1 = p_39_8 << 1;
  assign t_r39_c9_2 = p_39_9 << 2;
  assign t_r39_c9_3 = p_39_10 << 1;
  assign t_r39_c9_4 = p_40_9 << 1;
  assign t_r39_c9_5 = t_r39_c9_0 + p_38_8;
  assign t_r39_c9_6 = t_r39_c9_1 + p_38_10;
  assign t_r39_c9_7 = t_r39_c9_2 + t_r39_c9_3;
  assign t_r39_c9_8 = t_r39_c9_4 + p_40_8;
  assign t_r39_c9_9 = t_r39_c9_5 + t_r39_c9_6;
  assign t_r39_c9_10 = t_r39_c9_7 + t_r39_c9_8;
  assign t_r39_c9_11 = t_r39_c9_9 + t_r39_c9_10;
  assign t_r39_c9_12 = t_r39_c9_11 + p_40_10;
  assign out_39_9 = t_r39_c9_12 >> 4;

  assign t_r39_c10_0 = p_38_10 << 1;
  assign t_r39_c10_1 = p_39_9 << 1;
  assign t_r39_c10_2 = p_39_10 << 2;
  assign t_r39_c10_3 = p_39_11 << 1;
  assign t_r39_c10_4 = p_40_10 << 1;
  assign t_r39_c10_5 = t_r39_c10_0 + p_38_9;
  assign t_r39_c10_6 = t_r39_c10_1 + p_38_11;
  assign t_r39_c10_7 = t_r39_c10_2 + t_r39_c10_3;
  assign t_r39_c10_8 = t_r39_c10_4 + p_40_9;
  assign t_r39_c10_9 = t_r39_c10_5 + t_r39_c10_6;
  assign t_r39_c10_10 = t_r39_c10_7 + t_r39_c10_8;
  assign t_r39_c10_11 = t_r39_c10_9 + t_r39_c10_10;
  assign t_r39_c10_12 = t_r39_c10_11 + p_40_11;
  assign out_39_10 = t_r39_c10_12 >> 4;

  assign t_r39_c11_0 = p_38_11 << 1;
  assign t_r39_c11_1 = p_39_10 << 1;
  assign t_r39_c11_2 = p_39_11 << 2;
  assign t_r39_c11_3 = p_39_12 << 1;
  assign t_r39_c11_4 = p_40_11 << 1;
  assign t_r39_c11_5 = t_r39_c11_0 + p_38_10;
  assign t_r39_c11_6 = t_r39_c11_1 + p_38_12;
  assign t_r39_c11_7 = t_r39_c11_2 + t_r39_c11_3;
  assign t_r39_c11_8 = t_r39_c11_4 + p_40_10;
  assign t_r39_c11_9 = t_r39_c11_5 + t_r39_c11_6;
  assign t_r39_c11_10 = t_r39_c11_7 + t_r39_c11_8;
  assign t_r39_c11_11 = t_r39_c11_9 + t_r39_c11_10;
  assign t_r39_c11_12 = t_r39_c11_11 + p_40_12;
  assign out_39_11 = t_r39_c11_12 >> 4;

  assign t_r39_c12_0 = p_38_12 << 1;
  assign t_r39_c12_1 = p_39_11 << 1;
  assign t_r39_c12_2 = p_39_12 << 2;
  assign t_r39_c12_3 = p_39_13 << 1;
  assign t_r39_c12_4 = p_40_12 << 1;
  assign t_r39_c12_5 = t_r39_c12_0 + p_38_11;
  assign t_r39_c12_6 = t_r39_c12_1 + p_38_13;
  assign t_r39_c12_7 = t_r39_c12_2 + t_r39_c12_3;
  assign t_r39_c12_8 = t_r39_c12_4 + p_40_11;
  assign t_r39_c12_9 = t_r39_c12_5 + t_r39_c12_6;
  assign t_r39_c12_10 = t_r39_c12_7 + t_r39_c12_8;
  assign t_r39_c12_11 = t_r39_c12_9 + t_r39_c12_10;
  assign t_r39_c12_12 = t_r39_c12_11 + p_40_13;
  assign out_39_12 = t_r39_c12_12 >> 4;

  assign t_r39_c13_0 = p_38_13 << 1;
  assign t_r39_c13_1 = p_39_12 << 1;
  assign t_r39_c13_2 = p_39_13 << 2;
  assign t_r39_c13_3 = p_39_14 << 1;
  assign t_r39_c13_4 = p_40_13 << 1;
  assign t_r39_c13_5 = t_r39_c13_0 + p_38_12;
  assign t_r39_c13_6 = t_r39_c13_1 + p_38_14;
  assign t_r39_c13_7 = t_r39_c13_2 + t_r39_c13_3;
  assign t_r39_c13_8 = t_r39_c13_4 + p_40_12;
  assign t_r39_c13_9 = t_r39_c13_5 + t_r39_c13_6;
  assign t_r39_c13_10 = t_r39_c13_7 + t_r39_c13_8;
  assign t_r39_c13_11 = t_r39_c13_9 + t_r39_c13_10;
  assign t_r39_c13_12 = t_r39_c13_11 + p_40_14;
  assign out_39_13 = t_r39_c13_12 >> 4;

  assign t_r39_c14_0 = p_38_14 << 1;
  assign t_r39_c14_1 = p_39_13 << 1;
  assign t_r39_c14_2 = p_39_14 << 2;
  assign t_r39_c14_3 = p_39_15 << 1;
  assign t_r39_c14_4 = p_40_14 << 1;
  assign t_r39_c14_5 = t_r39_c14_0 + p_38_13;
  assign t_r39_c14_6 = t_r39_c14_1 + p_38_15;
  assign t_r39_c14_7 = t_r39_c14_2 + t_r39_c14_3;
  assign t_r39_c14_8 = t_r39_c14_4 + p_40_13;
  assign t_r39_c14_9 = t_r39_c14_5 + t_r39_c14_6;
  assign t_r39_c14_10 = t_r39_c14_7 + t_r39_c14_8;
  assign t_r39_c14_11 = t_r39_c14_9 + t_r39_c14_10;
  assign t_r39_c14_12 = t_r39_c14_11 + p_40_15;
  assign out_39_14 = t_r39_c14_12 >> 4;

  assign t_r39_c15_0 = p_38_15 << 1;
  assign t_r39_c15_1 = p_39_14 << 1;
  assign t_r39_c15_2 = p_39_15 << 2;
  assign t_r39_c15_3 = p_39_16 << 1;
  assign t_r39_c15_4 = p_40_15 << 1;
  assign t_r39_c15_5 = t_r39_c15_0 + p_38_14;
  assign t_r39_c15_6 = t_r39_c15_1 + p_38_16;
  assign t_r39_c15_7 = t_r39_c15_2 + t_r39_c15_3;
  assign t_r39_c15_8 = t_r39_c15_4 + p_40_14;
  assign t_r39_c15_9 = t_r39_c15_5 + t_r39_c15_6;
  assign t_r39_c15_10 = t_r39_c15_7 + t_r39_c15_8;
  assign t_r39_c15_11 = t_r39_c15_9 + t_r39_c15_10;
  assign t_r39_c15_12 = t_r39_c15_11 + p_40_16;
  assign out_39_15 = t_r39_c15_12 >> 4;

  assign t_r39_c16_0 = p_38_16 << 1;
  assign t_r39_c16_1 = p_39_15 << 1;
  assign t_r39_c16_2 = p_39_16 << 2;
  assign t_r39_c16_3 = p_39_17 << 1;
  assign t_r39_c16_4 = p_40_16 << 1;
  assign t_r39_c16_5 = t_r39_c16_0 + p_38_15;
  assign t_r39_c16_6 = t_r39_c16_1 + p_38_17;
  assign t_r39_c16_7 = t_r39_c16_2 + t_r39_c16_3;
  assign t_r39_c16_8 = t_r39_c16_4 + p_40_15;
  assign t_r39_c16_9 = t_r39_c16_5 + t_r39_c16_6;
  assign t_r39_c16_10 = t_r39_c16_7 + t_r39_c16_8;
  assign t_r39_c16_11 = t_r39_c16_9 + t_r39_c16_10;
  assign t_r39_c16_12 = t_r39_c16_11 + p_40_17;
  assign out_39_16 = t_r39_c16_12 >> 4;

  assign t_r39_c17_0 = p_38_17 << 1;
  assign t_r39_c17_1 = p_39_16 << 1;
  assign t_r39_c17_2 = p_39_17 << 2;
  assign t_r39_c17_3 = p_39_18 << 1;
  assign t_r39_c17_4 = p_40_17 << 1;
  assign t_r39_c17_5 = t_r39_c17_0 + p_38_16;
  assign t_r39_c17_6 = t_r39_c17_1 + p_38_18;
  assign t_r39_c17_7 = t_r39_c17_2 + t_r39_c17_3;
  assign t_r39_c17_8 = t_r39_c17_4 + p_40_16;
  assign t_r39_c17_9 = t_r39_c17_5 + t_r39_c17_6;
  assign t_r39_c17_10 = t_r39_c17_7 + t_r39_c17_8;
  assign t_r39_c17_11 = t_r39_c17_9 + t_r39_c17_10;
  assign t_r39_c17_12 = t_r39_c17_11 + p_40_18;
  assign out_39_17 = t_r39_c17_12 >> 4;

  assign t_r39_c18_0 = p_38_18 << 1;
  assign t_r39_c18_1 = p_39_17 << 1;
  assign t_r39_c18_2 = p_39_18 << 2;
  assign t_r39_c18_3 = p_39_19 << 1;
  assign t_r39_c18_4 = p_40_18 << 1;
  assign t_r39_c18_5 = t_r39_c18_0 + p_38_17;
  assign t_r39_c18_6 = t_r39_c18_1 + p_38_19;
  assign t_r39_c18_7 = t_r39_c18_2 + t_r39_c18_3;
  assign t_r39_c18_8 = t_r39_c18_4 + p_40_17;
  assign t_r39_c18_9 = t_r39_c18_5 + t_r39_c18_6;
  assign t_r39_c18_10 = t_r39_c18_7 + t_r39_c18_8;
  assign t_r39_c18_11 = t_r39_c18_9 + t_r39_c18_10;
  assign t_r39_c18_12 = t_r39_c18_11 + p_40_19;
  assign out_39_18 = t_r39_c18_12 >> 4;

  assign t_r39_c19_0 = p_38_19 << 1;
  assign t_r39_c19_1 = p_39_18 << 1;
  assign t_r39_c19_2 = p_39_19 << 2;
  assign t_r39_c19_3 = p_39_20 << 1;
  assign t_r39_c19_4 = p_40_19 << 1;
  assign t_r39_c19_5 = t_r39_c19_0 + p_38_18;
  assign t_r39_c19_6 = t_r39_c19_1 + p_38_20;
  assign t_r39_c19_7 = t_r39_c19_2 + t_r39_c19_3;
  assign t_r39_c19_8 = t_r39_c19_4 + p_40_18;
  assign t_r39_c19_9 = t_r39_c19_5 + t_r39_c19_6;
  assign t_r39_c19_10 = t_r39_c19_7 + t_r39_c19_8;
  assign t_r39_c19_11 = t_r39_c19_9 + t_r39_c19_10;
  assign t_r39_c19_12 = t_r39_c19_11 + p_40_20;
  assign out_39_19 = t_r39_c19_12 >> 4;

  assign t_r39_c20_0 = p_38_20 << 1;
  assign t_r39_c20_1 = p_39_19 << 1;
  assign t_r39_c20_2 = p_39_20 << 2;
  assign t_r39_c20_3 = p_39_21 << 1;
  assign t_r39_c20_4 = p_40_20 << 1;
  assign t_r39_c20_5 = t_r39_c20_0 + p_38_19;
  assign t_r39_c20_6 = t_r39_c20_1 + p_38_21;
  assign t_r39_c20_7 = t_r39_c20_2 + t_r39_c20_3;
  assign t_r39_c20_8 = t_r39_c20_4 + p_40_19;
  assign t_r39_c20_9 = t_r39_c20_5 + t_r39_c20_6;
  assign t_r39_c20_10 = t_r39_c20_7 + t_r39_c20_8;
  assign t_r39_c20_11 = t_r39_c20_9 + t_r39_c20_10;
  assign t_r39_c20_12 = t_r39_c20_11 + p_40_21;
  assign out_39_20 = t_r39_c20_12 >> 4;

  assign t_r39_c21_0 = p_38_21 << 1;
  assign t_r39_c21_1 = p_39_20 << 1;
  assign t_r39_c21_2 = p_39_21 << 2;
  assign t_r39_c21_3 = p_39_22 << 1;
  assign t_r39_c21_4 = p_40_21 << 1;
  assign t_r39_c21_5 = t_r39_c21_0 + p_38_20;
  assign t_r39_c21_6 = t_r39_c21_1 + p_38_22;
  assign t_r39_c21_7 = t_r39_c21_2 + t_r39_c21_3;
  assign t_r39_c21_8 = t_r39_c21_4 + p_40_20;
  assign t_r39_c21_9 = t_r39_c21_5 + t_r39_c21_6;
  assign t_r39_c21_10 = t_r39_c21_7 + t_r39_c21_8;
  assign t_r39_c21_11 = t_r39_c21_9 + t_r39_c21_10;
  assign t_r39_c21_12 = t_r39_c21_11 + p_40_22;
  assign out_39_21 = t_r39_c21_12 >> 4;

  assign t_r39_c22_0 = p_38_22 << 1;
  assign t_r39_c22_1 = p_39_21 << 1;
  assign t_r39_c22_2 = p_39_22 << 2;
  assign t_r39_c22_3 = p_39_23 << 1;
  assign t_r39_c22_4 = p_40_22 << 1;
  assign t_r39_c22_5 = t_r39_c22_0 + p_38_21;
  assign t_r39_c22_6 = t_r39_c22_1 + p_38_23;
  assign t_r39_c22_7 = t_r39_c22_2 + t_r39_c22_3;
  assign t_r39_c22_8 = t_r39_c22_4 + p_40_21;
  assign t_r39_c22_9 = t_r39_c22_5 + t_r39_c22_6;
  assign t_r39_c22_10 = t_r39_c22_7 + t_r39_c22_8;
  assign t_r39_c22_11 = t_r39_c22_9 + t_r39_c22_10;
  assign t_r39_c22_12 = t_r39_c22_11 + p_40_23;
  assign out_39_22 = t_r39_c22_12 >> 4;

  assign t_r39_c23_0 = p_38_23 << 1;
  assign t_r39_c23_1 = p_39_22 << 1;
  assign t_r39_c23_2 = p_39_23 << 2;
  assign t_r39_c23_3 = p_39_24 << 1;
  assign t_r39_c23_4 = p_40_23 << 1;
  assign t_r39_c23_5 = t_r39_c23_0 + p_38_22;
  assign t_r39_c23_6 = t_r39_c23_1 + p_38_24;
  assign t_r39_c23_7 = t_r39_c23_2 + t_r39_c23_3;
  assign t_r39_c23_8 = t_r39_c23_4 + p_40_22;
  assign t_r39_c23_9 = t_r39_c23_5 + t_r39_c23_6;
  assign t_r39_c23_10 = t_r39_c23_7 + t_r39_c23_8;
  assign t_r39_c23_11 = t_r39_c23_9 + t_r39_c23_10;
  assign t_r39_c23_12 = t_r39_c23_11 + p_40_24;
  assign out_39_23 = t_r39_c23_12 >> 4;

  assign t_r39_c24_0 = p_38_24 << 1;
  assign t_r39_c24_1 = p_39_23 << 1;
  assign t_r39_c24_2 = p_39_24 << 2;
  assign t_r39_c24_3 = p_39_25 << 1;
  assign t_r39_c24_4 = p_40_24 << 1;
  assign t_r39_c24_5 = t_r39_c24_0 + p_38_23;
  assign t_r39_c24_6 = t_r39_c24_1 + p_38_25;
  assign t_r39_c24_7 = t_r39_c24_2 + t_r39_c24_3;
  assign t_r39_c24_8 = t_r39_c24_4 + p_40_23;
  assign t_r39_c24_9 = t_r39_c24_5 + t_r39_c24_6;
  assign t_r39_c24_10 = t_r39_c24_7 + t_r39_c24_8;
  assign t_r39_c24_11 = t_r39_c24_9 + t_r39_c24_10;
  assign t_r39_c24_12 = t_r39_c24_11 + p_40_25;
  assign out_39_24 = t_r39_c24_12 >> 4;

  assign t_r39_c25_0 = p_38_25 << 1;
  assign t_r39_c25_1 = p_39_24 << 1;
  assign t_r39_c25_2 = p_39_25 << 2;
  assign t_r39_c25_3 = p_39_26 << 1;
  assign t_r39_c25_4 = p_40_25 << 1;
  assign t_r39_c25_5 = t_r39_c25_0 + p_38_24;
  assign t_r39_c25_6 = t_r39_c25_1 + p_38_26;
  assign t_r39_c25_7 = t_r39_c25_2 + t_r39_c25_3;
  assign t_r39_c25_8 = t_r39_c25_4 + p_40_24;
  assign t_r39_c25_9 = t_r39_c25_5 + t_r39_c25_6;
  assign t_r39_c25_10 = t_r39_c25_7 + t_r39_c25_8;
  assign t_r39_c25_11 = t_r39_c25_9 + t_r39_c25_10;
  assign t_r39_c25_12 = t_r39_c25_11 + p_40_26;
  assign out_39_25 = t_r39_c25_12 >> 4;

  assign t_r39_c26_0 = p_38_26 << 1;
  assign t_r39_c26_1 = p_39_25 << 1;
  assign t_r39_c26_2 = p_39_26 << 2;
  assign t_r39_c26_3 = p_39_27 << 1;
  assign t_r39_c26_4 = p_40_26 << 1;
  assign t_r39_c26_5 = t_r39_c26_0 + p_38_25;
  assign t_r39_c26_6 = t_r39_c26_1 + p_38_27;
  assign t_r39_c26_7 = t_r39_c26_2 + t_r39_c26_3;
  assign t_r39_c26_8 = t_r39_c26_4 + p_40_25;
  assign t_r39_c26_9 = t_r39_c26_5 + t_r39_c26_6;
  assign t_r39_c26_10 = t_r39_c26_7 + t_r39_c26_8;
  assign t_r39_c26_11 = t_r39_c26_9 + t_r39_c26_10;
  assign t_r39_c26_12 = t_r39_c26_11 + p_40_27;
  assign out_39_26 = t_r39_c26_12 >> 4;

  assign t_r39_c27_0 = p_38_27 << 1;
  assign t_r39_c27_1 = p_39_26 << 1;
  assign t_r39_c27_2 = p_39_27 << 2;
  assign t_r39_c27_3 = p_39_28 << 1;
  assign t_r39_c27_4 = p_40_27 << 1;
  assign t_r39_c27_5 = t_r39_c27_0 + p_38_26;
  assign t_r39_c27_6 = t_r39_c27_1 + p_38_28;
  assign t_r39_c27_7 = t_r39_c27_2 + t_r39_c27_3;
  assign t_r39_c27_8 = t_r39_c27_4 + p_40_26;
  assign t_r39_c27_9 = t_r39_c27_5 + t_r39_c27_6;
  assign t_r39_c27_10 = t_r39_c27_7 + t_r39_c27_8;
  assign t_r39_c27_11 = t_r39_c27_9 + t_r39_c27_10;
  assign t_r39_c27_12 = t_r39_c27_11 + p_40_28;
  assign out_39_27 = t_r39_c27_12 >> 4;

  assign t_r39_c28_0 = p_38_28 << 1;
  assign t_r39_c28_1 = p_39_27 << 1;
  assign t_r39_c28_2 = p_39_28 << 2;
  assign t_r39_c28_3 = p_39_29 << 1;
  assign t_r39_c28_4 = p_40_28 << 1;
  assign t_r39_c28_5 = t_r39_c28_0 + p_38_27;
  assign t_r39_c28_6 = t_r39_c28_1 + p_38_29;
  assign t_r39_c28_7 = t_r39_c28_2 + t_r39_c28_3;
  assign t_r39_c28_8 = t_r39_c28_4 + p_40_27;
  assign t_r39_c28_9 = t_r39_c28_5 + t_r39_c28_6;
  assign t_r39_c28_10 = t_r39_c28_7 + t_r39_c28_8;
  assign t_r39_c28_11 = t_r39_c28_9 + t_r39_c28_10;
  assign t_r39_c28_12 = t_r39_c28_11 + p_40_29;
  assign out_39_28 = t_r39_c28_12 >> 4;

  assign t_r39_c29_0 = p_38_29 << 1;
  assign t_r39_c29_1 = p_39_28 << 1;
  assign t_r39_c29_2 = p_39_29 << 2;
  assign t_r39_c29_3 = p_39_30 << 1;
  assign t_r39_c29_4 = p_40_29 << 1;
  assign t_r39_c29_5 = t_r39_c29_0 + p_38_28;
  assign t_r39_c29_6 = t_r39_c29_1 + p_38_30;
  assign t_r39_c29_7 = t_r39_c29_2 + t_r39_c29_3;
  assign t_r39_c29_8 = t_r39_c29_4 + p_40_28;
  assign t_r39_c29_9 = t_r39_c29_5 + t_r39_c29_6;
  assign t_r39_c29_10 = t_r39_c29_7 + t_r39_c29_8;
  assign t_r39_c29_11 = t_r39_c29_9 + t_r39_c29_10;
  assign t_r39_c29_12 = t_r39_c29_11 + p_40_30;
  assign out_39_29 = t_r39_c29_12 >> 4;

  assign t_r39_c30_0 = p_38_30 << 1;
  assign t_r39_c30_1 = p_39_29 << 1;
  assign t_r39_c30_2 = p_39_30 << 2;
  assign t_r39_c30_3 = p_39_31 << 1;
  assign t_r39_c30_4 = p_40_30 << 1;
  assign t_r39_c30_5 = t_r39_c30_0 + p_38_29;
  assign t_r39_c30_6 = t_r39_c30_1 + p_38_31;
  assign t_r39_c30_7 = t_r39_c30_2 + t_r39_c30_3;
  assign t_r39_c30_8 = t_r39_c30_4 + p_40_29;
  assign t_r39_c30_9 = t_r39_c30_5 + t_r39_c30_6;
  assign t_r39_c30_10 = t_r39_c30_7 + t_r39_c30_8;
  assign t_r39_c30_11 = t_r39_c30_9 + t_r39_c30_10;
  assign t_r39_c30_12 = t_r39_c30_11 + p_40_31;
  assign out_39_30 = t_r39_c30_12 >> 4;

  assign t_r39_c31_0 = p_38_31 << 1;
  assign t_r39_c31_1 = p_39_30 << 1;
  assign t_r39_c31_2 = p_39_31 << 2;
  assign t_r39_c31_3 = p_39_32 << 1;
  assign t_r39_c31_4 = p_40_31 << 1;
  assign t_r39_c31_5 = t_r39_c31_0 + p_38_30;
  assign t_r39_c31_6 = t_r39_c31_1 + p_38_32;
  assign t_r39_c31_7 = t_r39_c31_2 + t_r39_c31_3;
  assign t_r39_c31_8 = t_r39_c31_4 + p_40_30;
  assign t_r39_c31_9 = t_r39_c31_5 + t_r39_c31_6;
  assign t_r39_c31_10 = t_r39_c31_7 + t_r39_c31_8;
  assign t_r39_c31_11 = t_r39_c31_9 + t_r39_c31_10;
  assign t_r39_c31_12 = t_r39_c31_11 + p_40_32;
  assign out_39_31 = t_r39_c31_12 >> 4;

  assign t_r39_c32_0 = p_38_32 << 1;
  assign t_r39_c32_1 = p_39_31 << 1;
  assign t_r39_c32_2 = p_39_32 << 2;
  assign t_r39_c32_3 = p_39_33 << 1;
  assign t_r39_c32_4 = p_40_32 << 1;
  assign t_r39_c32_5 = t_r39_c32_0 + p_38_31;
  assign t_r39_c32_6 = t_r39_c32_1 + p_38_33;
  assign t_r39_c32_7 = t_r39_c32_2 + t_r39_c32_3;
  assign t_r39_c32_8 = t_r39_c32_4 + p_40_31;
  assign t_r39_c32_9 = t_r39_c32_5 + t_r39_c32_6;
  assign t_r39_c32_10 = t_r39_c32_7 + t_r39_c32_8;
  assign t_r39_c32_11 = t_r39_c32_9 + t_r39_c32_10;
  assign t_r39_c32_12 = t_r39_c32_11 + p_40_33;
  assign out_39_32 = t_r39_c32_12 >> 4;

  assign t_r39_c33_0 = p_38_33 << 1;
  assign t_r39_c33_1 = p_39_32 << 1;
  assign t_r39_c33_2 = p_39_33 << 2;
  assign t_r39_c33_3 = p_39_34 << 1;
  assign t_r39_c33_4 = p_40_33 << 1;
  assign t_r39_c33_5 = t_r39_c33_0 + p_38_32;
  assign t_r39_c33_6 = t_r39_c33_1 + p_38_34;
  assign t_r39_c33_7 = t_r39_c33_2 + t_r39_c33_3;
  assign t_r39_c33_8 = t_r39_c33_4 + p_40_32;
  assign t_r39_c33_9 = t_r39_c33_5 + t_r39_c33_6;
  assign t_r39_c33_10 = t_r39_c33_7 + t_r39_c33_8;
  assign t_r39_c33_11 = t_r39_c33_9 + t_r39_c33_10;
  assign t_r39_c33_12 = t_r39_c33_11 + p_40_34;
  assign out_39_33 = t_r39_c33_12 >> 4;

  assign t_r39_c34_0 = p_38_34 << 1;
  assign t_r39_c34_1 = p_39_33 << 1;
  assign t_r39_c34_2 = p_39_34 << 2;
  assign t_r39_c34_3 = p_39_35 << 1;
  assign t_r39_c34_4 = p_40_34 << 1;
  assign t_r39_c34_5 = t_r39_c34_0 + p_38_33;
  assign t_r39_c34_6 = t_r39_c34_1 + p_38_35;
  assign t_r39_c34_7 = t_r39_c34_2 + t_r39_c34_3;
  assign t_r39_c34_8 = t_r39_c34_4 + p_40_33;
  assign t_r39_c34_9 = t_r39_c34_5 + t_r39_c34_6;
  assign t_r39_c34_10 = t_r39_c34_7 + t_r39_c34_8;
  assign t_r39_c34_11 = t_r39_c34_9 + t_r39_c34_10;
  assign t_r39_c34_12 = t_r39_c34_11 + p_40_35;
  assign out_39_34 = t_r39_c34_12 >> 4;

  assign t_r39_c35_0 = p_38_35 << 1;
  assign t_r39_c35_1 = p_39_34 << 1;
  assign t_r39_c35_2 = p_39_35 << 2;
  assign t_r39_c35_3 = p_39_36 << 1;
  assign t_r39_c35_4 = p_40_35 << 1;
  assign t_r39_c35_5 = t_r39_c35_0 + p_38_34;
  assign t_r39_c35_6 = t_r39_c35_1 + p_38_36;
  assign t_r39_c35_7 = t_r39_c35_2 + t_r39_c35_3;
  assign t_r39_c35_8 = t_r39_c35_4 + p_40_34;
  assign t_r39_c35_9 = t_r39_c35_5 + t_r39_c35_6;
  assign t_r39_c35_10 = t_r39_c35_7 + t_r39_c35_8;
  assign t_r39_c35_11 = t_r39_c35_9 + t_r39_c35_10;
  assign t_r39_c35_12 = t_r39_c35_11 + p_40_36;
  assign out_39_35 = t_r39_c35_12 >> 4;

  assign t_r39_c36_0 = p_38_36 << 1;
  assign t_r39_c36_1 = p_39_35 << 1;
  assign t_r39_c36_2 = p_39_36 << 2;
  assign t_r39_c36_3 = p_39_37 << 1;
  assign t_r39_c36_4 = p_40_36 << 1;
  assign t_r39_c36_5 = t_r39_c36_0 + p_38_35;
  assign t_r39_c36_6 = t_r39_c36_1 + p_38_37;
  assign t_r39_c36_7 = t_r39_c36_2 + t_r39_c36_3;
  assign t_r39_c36_8 = t_r39_c36_4 + p_40_35;
  assign t_r39_c36_9 = t_r39_c36_5 + t_r39_c36_6;
  assign t_r39_c36_10 = t_r39_c36_7 + t_r39_c36_8;
  assign t_r39_c36_11 = t_r39_c36_9 + t_r39_c36_10;
  assign t_r39_c36_12 = t_r39_c36_11 + p_40_37;
  assign out_39_36 = t_r39_c36_12 >> 4;

  assign t_r39_c37_0 = p_38_37 << 1;
  assign t_r39_c37_1 = p_39_36 << 1;
  assign t_r39_c37_2 = p_39_37 << 2;
  assign t_r39_c37_3 = p_39_38 << 1;
  assign t_r39_c37_4 = p_40_37 << 1;
  assign t_r39_c37_5 = t_r39_c37_0 + p_38_36;
  assign t_r39_c37_6 = t_r39_c37_1 + p_38_38;
  assign t_r39_c37_7 = t_r39_c37_2 + t_r39_c37_3;
  assign t_r39_c37_8 = t_r39_c37_4 + p_40_36;
  assign t_r39_c37_9 = t_r39_c37_5 + t_r39_c37_6;
  assign t_r39_c37_10 = t_r39_c37_7 + t_r39_c37_8;
  assign t_r39_c37_11 = t_r39_c37_9 + t_r39_c37_10;
  assign t_r39_c37_12 = t_r39_c37_11 + p_40_38;
  assign out_39_37 = t_r39_c37_12 >> 4;

  assign t_r39_c38_0 = p_38_38 << 1;
  assign t_r39_c38_1 = p_39_37 << 1;
  assign t_r39_c38_2 = p_39_38 << 2;
  assign t_r39_c38_3 = p_39_39 << 1;
  assign t_r39_c38_4 = p_40_38 << 1;
  assign t_r39_c38_5 = t_r39_c38_0 + p_38_37;
  assign t_r39_c38_6 = t_r39_c38_1 + p_38_39;
  assign t_r39_c38_7 = t_r39_c38_2 + t_r39_c38_3;
  assign t_r39_c38_8 = t_r39_c38_4 + p_40_37;
  assign t_r39_c38_9 = t_r39_c38_5 + t_r39_c38_6;
  assign t_r39_c38_10 = t_r39_c38_7 + t_r39_c38_8;
  assign t_r39_c38_11 = t_r39_c38_9 + t_r39_c38_10;
  assign t_r39_c38_12 = t_r39_c38_11 + p_40_39;
  assign out_39_38 = t_r39_c38_12 >> 4;

  assign t_r39_c39_0 = p_38_39 << 1;
  assign t_r39_c39_1 = p_39_38 << 1;
  assign t_r39_c39_2 = p_39_39 << 2;
  assign t_r39_c39_3 = p_39_40 << 1;
  assign t_r39_c39_4 = p_40_39 << 1;
  assign t_r39_c39_5 = t_r39_c39_0 + p_38_38;
  assign t_r39_c39_6 = t_r39_c39_1 + p_38_40;
  assign t_r39_c39_7 = t_r39_c39_2 + t_r39_c39_3;
  assign t_r39_c39_8 = t_r39_c39_4 + p_40_38;
  assign t_r39_c39_9 = t_r39_c39_5 + t_r39_c39_6;
  assign t_r39_c39_10 = t_r39_c39_7 + t_r39_c39_8;
  assign t_r39_c39_11 = t_r39_c39_9 + t_r39_c39_10;
  assign t_r39_c39_12 = t_r39_c39_11 + p_40_40;
  assign out_39_39 = t_r39_c39_12 >> 4;

  assign t_r39_c40_0 = p_38_40 << 1;
  assign t_r39_c40_1 = p_39_39 << 1;
  assign t_r39_c40_2 = p_39_40 << 2;
  assign t_r39_c40_3 = p_39_41 << 1;
  assign t_r39_c40_4 = p_40_40 << 1;
  assign t_r39_c40_5 = t_r39_c40_0 + p_38_39;
  assign t_r39_c40_6 = t_r39_c40_1 + p_38_41;
  assign t_r39_c40_7 = t_r39_c40_2 + t_r39_c40_3;
  assign t_r39_c40_8 = t_r39_c40_4 + p_40_39;
  assign t_r39_c40_9 = t_r39_c40_5 + t_r39_c40_6;
  assign t_r39_c40_10 = t_r39_c40_7 + t_r39_c40_8;
  assign t_r39_c40_11 = t_r39_c40_9 + t_r39_c40_10;
  assign t_r39_c40_12 = t_r39_c40_11 + p_40_41;
  assign out_39_40 = t_r39_c40_12 >> 4;

  assign t_r39_c41_0 = p_38_41 << 1;
  assign t_r39_c41_1 = p_39_40 << 1;
  assign t_r39_c41_2 = p_39_41 << 2;
  assign t_r39_c41_3 = p_39_42 << 1;
  assign t_r39_c41_4 = p_40_41 << 1;
  assign t_r39_c41_5 = t_r39_c41_0 + p_38_40;
  assign t_r39_c41_6 = t_r39_c41_1 + p_38_42;
  assign t_r39_c41_7 = t_r39_c41_2 + t_r39_c41_3;
  assign t_r39_c41_8 = t_r39_c41_4 + p_40_40;
  assign t_r39_c41_9 = t_r39_c41_5 + t_r39_c41_6;
  assign t_r39_c41_10 = t_r39_c41_7 + t_r39_c41_8;
  assign t_r39_c41_11 = t_r39_c41_9 + t_r39_c41_10;
  assign t_r39_c41_12 = t_r39_c41_11 + p_40_42;
  assign out_39_41 = t_r39_c41_12 >> 4;

  assign t_r39_c42_0 = p_38_42 << 1;
  assign t_r39_c42_1 = p_39_41 << 1;
  assign t_r39_c42_2 = p_39_42 << 2;
  assign t_r39_c42_3 = p_39_43 << 1;
  assign t_r39_c42_4 = p_40_42 << 1;
  assign t_r39_c42_5 = t_r39_c42_0 + p_38_41;
  assign t_r39_c42_6 = t_r39_c42_1 + p_38_43;
  assign t_r39_c42_7 = t_r39_c42_2 + t_r39_c42_3;
  assign t_r39_c42_8 = t_r39_c42_4 + p_40_41;
  assign t_r39_c42_9 = t_r39_c42_5 + t_r39_c42_6;
  assign t_r39_c42_10 = t_r39_c42_7 + t_r39_c42_8;
  assign t_r39_c42_11 = t_r39_c42_9 + t_r39_c42_10;
  assign t_r39_c42_12 = t_r39_c42_11 + p_40_43;
  assign out_39_42 = t_r39_c42_12 >> 4;

  assign t_r39_c43_0 = p_38_43 << 1;
  assign t_r39_c43_1 = p_39_42 << 1;
  assign t_r39_c43_2 = p_39_43 << 2;
  assign t_r39_c43_3 = p_39_44 << 1;
  assign t_r39_c43_4 = p_40_43 << 1;
  assign t_r39_c43_5 = t_r39_c43_0 + p_38_42;
  assign t_r39_c43_6 = t_r39_c43_1 + p_38_44;
  assign t_r39_c43_7 = t_r39_c43_2 + t_r39_c43_3;
  assign t_r39_c43_8 = t_r39_c43_4 + p_40_42;
  assign t_r39_c43_9 = t_r39_c43_5 + t_r39_c43_6;
  assign t_r39_c43_10 = t_r39_c43_7 + t_r39_c43_8;
  assign t_r39_c43_11 = t_r39_c43_9 + t_r39_c43_10;
  assign t_r39_c43_12 = t_r39_c43_11 + p_40_44;
  assign out_39_43 = t_r39_c43_12 >> 4;

  assign t_r39_c44_0 = p_38_44 << 1;
  assign t_r39_c44_1 = p_39_43 << 1;
  assign t_r39_c44_2 = p_39_44 << 2;
  assign t_r39_c44_3 = p_39_45 << 1;
  assign t_r39_c44_4 = p_40_44 << 1;
  assign t_r39_c44_5 = t_r39_c44_0 + p_38_43;
  assign t_r39_c44_6 = t_r39_c44_1 + p_38_45;
  assign t_r39_c44_7 = t_r39_c44_2 + t_r39_c44_3;
  assign t_r39_c44_8 = t_r39_c44_4 + p_40_43;
  assign t_r39_c44_9 = t_r39_c44_5 + t_r39_c44_6;
  assign t_r39_c44_10 = t_r39_c44_7 + t_r39_c44_8;
  assign t_r39_c44_11 = t_r39_c44_9 + t_r39_c44_10;
  assign t_r39_c44_12 = t_r39_c44_11 + p_40_45;
  assign out_39_44 = t_r39_c44_12 >> 4;

  assign t_r39_c45_0 = p_38_45 << 1;
  assign t_r39_c45_1 = p_39_44 << 1;
  assign t_r39_c45_2 = p_39_45 << 2;
  assign t_r39_c45_3 = p_39_46 << 1;
  assign t_r39_c45_4 = p_40_45 << 1;
  assign t_r39_c45_5 = t_r39_c45_0 + p_38_44;
  assign t_r39_c45_6 = t_r39_c45_1 + p_38_46;
  assign t_r39_c45_7 = t_r39_c45_2 + t_r39_c45_3;
  assign t_r39_c45_8 = t_r39_c45_4 + p_40_44;
  assign t_r39_c45_9 = t_r39_c45_5 + t_r39_c45_6;
  assign t_r39_c45_10 = t_r39_c45_7 + t_r39_c45_8;
  assign t_r39_c45_11 = t_r39_c45_9 + t_r39_c45_10;
  assign t_r39_c45_12 = t_r39_c45_11 + p_40_46;
  assign out_39_45 = t_r39_c45_12 >> 4;

  assign t_r39_c46_0 = p_38_46 << 1;
  assign t_r39_c46_1 = p_39_45 << 1;
  assign t_r39_c46_2 = p_39_46 << 2;
  assign t_r39_c46_3 = p_39_47 << 1;
  assign t_r39_c46_4 = p_40_46 << 1;
  assign t_r39_c46_5 = t_r39_c46_0 + p_38_45;
  assign t_r39_c46_6 = t_r39_c46_1 + p_38_47;
  assign t_r39_c46_7 = t_r39_c46_2 + t_r39_c46_3;
  assign t_r39_c46_8 = t_r39_c46_4 + p_40_45;
  assign t_r39_c46_9 = t_r39_c46_5 + t_r39_c46_6;
  assign t_r39_c46_10 = t_r39_c46_7 + t_r39_c46_8;
  assign t_r39_c46_11 = t_r39_c46_9 + t_r39_c46_10;
  assign t_r39_c46_12 = t_r39_c46_11 + p_40_47;
  assign out_39_46 = t_r39_c46_12 >> 4;

  assign t_r39_c47_0 = p_38_47 << 1;
  assign t_r39_c47_1 = p_39_46 << 1;
  assign t_r39_c47_2 = p_39_47 << 2;
  assign t_r39_c47_3 = p_39_48 << 1;
  assign t_r39_c47_4 = p_40_47 << 1;
  assign t_r39_c47_5 = t_r39_c47_0 + p_38_46;
  assign t_r39_c47_6 = t_r39_c47_1 + p_38_48;
  assign t_r39_c47_7 = t_r39_c47_2 + t_r39_c47_3;
  assign t_r39_c47_8 = t_r39_c47_4 + p_40_46;
  assign t_r39_c47_9 = t_r39_c47_5 + t_r39_c47_6;
  assign t_r39_c47_10 = t_r39_c47_7 + t_r39_c47_8;
  assign t_r39_c47_11 = t_r39_c47_9 + t_r39_c47_10;
  assign t_r39_c47_12 = t_r39_c47_11 + p_40_48;
  assign out_39_47 = t_r39_c47_12 >> 4;

  assign t_r39_c48_0 = p_38_48 << 1;
  assign t_r39_c48_1 = p_39_47 << 1;
  assign t_r39_c48_2 = p_39_48 << 2;
  assign t_r39_c48_3 = p_39_49 << 1;
  assign t_r39_c48_4 = p_40_48 << 1;
  assign t_r39_c48_5 = t_r39_c48_0 + p_38_47;
  assign t_r39_c48_6 = t_r39_c48_1 + p_38_49;
  assign t_r39_c48_7 = t_r39_c48_2 + t_r39_c48_3;
  assign t_r39_c48_8 = t_r39_c48_4 + p_40_47;
  assign t_r39_c48_9 = t_r39_c48_5 + t_r39_c48_6;
  assign t_r39_c48_10 = t_r39_c48_7 + t_r39_c48_8;
  assign t_r39_c48_11 = t_r39_c48_9 + t_r39_c48_10;
  assign t_r39_c48_12 = t_r39_c48_11 + p_40_49;
  assign out_39_48 = t_r39_c48_12 >> 4;

  assign t_r39_c49_0 = p_38_49 << 1;
  assign t_r39_c49_1 = p_39_48 << 1;
  assign t_r39_c49_2 = p_39_49 << 2;
  assign t_r39_c49_3 = p_39_50 << 1;
  assign t_r39_c49_4 = p_40_49 << 1;
  assign t_r39_c49_5 = t_r39_c49_0 + p_38_48;
  assign t_r39_c49_6 = t_r39_c49_1 + p_38_50;
  assign t_r39_c49_7 = t_r39_c49_2 + t_r39_c49_3;
  assign t_r39_c49_8 = t_r39_c49_4 + p_40_48;
  assign t_r39_c49_9 = t_r39_c49_5 + t_r39_c49_6;
  assign t_r39_c49_10 = t_r39_c49_7 + t_r39_c49_8;
  assign t_r39_c49_11 = t_r39_c49_9 + t_r39_c49_10;
  assign t_r39_c49_12 = t_r39_c49_11 + p_40_50;
  assign out_39_49 = t_r39_c49_12 >> 4;

  assign t_r39_c50_0 = p_38_50 << 1;
  assign t_r39_c50_1 = p_39_49 << 1;
  assign t_r39_c50_2 = p_39_50 << 2;
  assign t_r39_c50_3 = p_39_51 << 1;
  assign t_r39_c50_4 = p_40_50 << 1;
  assign t_r39_c50_5 = t_r39_c50_0 + p_38_49;
  assign t_r39_c50_6 = t_r39_c50_1 + p_38_51;
  assign t_r39_c50_7 = t_r39_c50_2 + t_r39_c50_3;
  assign t_r39_c50_8 = t_r39_c50_4 + p_40_49;
  assign t_r39_c50_9 = t_r39_c50_5 + t_r39_c50_6;
  assign t_r39_c50_10 = t_r39_c50_7 + t_r39_c50_8;
  assign t_r39_c50_11 = t_r39_c50_9 + t_r39_c50_10;
  assign t_r39_c50_12 = t_r39_c50_11 + p_40_51;
  assign out_39_50 = t_r39_c50_12 >> 4;

  assign t_r39_c51_0 = p_38_51 << 1;
  assign t_r39_c51_1 = p_39_50 << 1;
  assign t_r39_c51_2 = p_39_51 << 2;
  assign t_r39_c51_3 = p_39_52 << 1;
  assign t_r39_c51_4 = p_40_51 << 1;
  assign t_r39_c51_5 = t_r39_c51_0 + p_38_50;
  assign t_r39_c51_6 = t_r39_c51_1 + p_38_52;
  assign t_r39_c51_7 = t_r39_c51_2 + t_r39_c51_3;
  assign t_r39_c51_8 = t_r39_c51_4 + p_40_50;
  assign t_r39_c51_9 = t_r39_c51_5 + t_r39_c51_6;
  assign t_r39_c51_10 = t_r39_c51_7 + t_r39_c51_8;
  assign t_r39_c51_11 = t_r39_c51_9 + t_r39_c51_10;
  assign t_r39_c51_12 = t_r39_c51_11 + p_40_52;
  assign out_39_51 = t_r39_c51_12 >> 4;

  assign t_r39_c52_0 = p_38_52 << 1;
  assign t_r39_c52_1 = p_39_51 << 1;
  assign t_r39_c52_2 = p_39_52 << 2;
  assign t_r39_c52_3 = p_39_53 << 1;
  assign t_r39_c52_4 = p_40_52 << 1;
  assign t_r39_c52_5 = t_r39_c52_0 + p_38_51;
  assign t_r39_c52_6 = t_r39_c52_1 + p_38_53;
  assign t_r39_c52_7 = t_r39_c52_2 + t_r39_c52_3;
  assign t_r39_c52_8 = t_r39_c52_4 + p_40_51;
  assign t_r39_c52_9 = t_r39_c52_5 + t_r39_c52_6;
  assign t_r39_c52_10 = t_r39_c52_7 + t_r39_c52_8;
  assign t_r39_c52_11 = t_r39_c52_9 + t_r39_c52_10;
  assign t_r39_c52_12 = t_r39_c52_11 + p_40_53;
  assign out_39_52 = t_r39_c52_12 >> 4;

  assign t_r39_c53_0 = p_38_53 << 1;
  assign t_r39_c53_1 = p_39_52 << 1;
  assign t_r39_c53_2 = p_39_53 << 2;
  assign t_r39_c53_3 = p_39_54 << 1;
  assign t_r39_c53_4 = p_40_53 << 1;
  assign t_r39_c53_5 = t_r39_c53_0 + p_38_52;
  assign t_r39_c53_6 = t_r39_c53_1 + p_38_54;
  assign t_r39_c53_7 = t_r39_c53_2 + t_r39_c53_3;
  assign t_r39_c53_8 = t_r39_c53_4 + p_40_52;
  assign t_r39_c53_9 = t_r39_c53_5 + t_r39_c53_6;
  assign t_r39_c53_10 = t_r39_c53_7 + t_r39_c53_8;
  assign t_r39_c53_11 = t_r39_c53_9 + t_r39_c53_10;
  assign t_r39_c53_12 = t_r39_c53_11 + p_40_54;
  assign out_39_53 = t_r39_c53_12 >> 4;

  assign t_r39_c54_0 = p_38_54 << 1;
  assign t_r39_c54_1 = p_39_53 << 1;
  assign t_r39_c54_2 = p_39_54 << 2;
  assign t_r39_c54_3 = p_39_55 << 1;
  assign t_r39_c54_4 = p_40_54 << 1;
  assign t_r39_c54_5 = t_r39_c54_0 + p_38_53;
  assign t_r39_c54_6 = t_r39_c54_1 + p_38_55;
  assign t_r39_c54_7 = t_r39_c54_2 + t_r39_c54_3;
  assign t_r39_c54_8 = t_r39_c54_4 + p_40_53;
  assign t_r39_c54_9 = t_r39_c54_5 + t_r39_c54_6;
  assign t_r39_c54_10 = t_r39_c54_7 + t_r39_c54_8;
  assign t_r39_c54_11 = t_r39_c54_9 + t_r39_c54_10;
  assign t_r39_c54_12 = t_r39_c54_11 + p_40_55;
  assign out_39_54 = t_r39_c54_12 >> 4;

  assign t_r39_c55_0 = p_38_55 << 1;
  assign t_r39_c55_1 = p_39_54 << 1;
  assign t_r39_c55_2 = p_39_55 << 2;
  assign t_r39_c55_3 = p_39_56 << 1;
  assign t_r39_c55_4 = p_40_55 << 1;
  assign t_r39_c55_5 = t_r39_c55_0 + p_38_54;
  assign t_r39_c55_6 = t_r39_c55_1 + p_38_56;
  assign t_r39_c55_7 = t_r39_c55_2 + t_r39_c55_3;
  assign t_r39_c55_8 = t_r39_c55_4 + p_40_54;
  assign t_r39_c55_9 = t_r39_c55_5 + t_r39_c55_6;
  assign t_r39_c55_10 = t_r39_c55_7 + t_r39_c55_8;
  assign t_r39_c55_11 = t_r39_c55_9 + t_r39_c55_10;
  assign t_r39_c55_12 = t_r39_c55_11 + p_40_56;
  assign out_39_55 = t_r39_c55_12 >> 4;

  assign t_r39_c56_0 = p_38_56 << 1;
  assign t_r39_c56_1 = p_39_55 << 1;
  assign t_r39_c56_2 = p_39_56 << 2;
  assign t_r39_c56_3 = p_39_57 << 1;
  assign t_r39_c56_4 = p_40_56 << 1;
  assign t_r39_c56_5 = t_r39_c56_0 + p_38_55;
  assign t_r39_c56_6 = t_r39_c56_1 + p_38_57;
  assign t_r39_c56_7 = t_r39_c56_2 + t_r39_c56_3;
  assign t_r39_c56_8 = t_r39_c56_4 + p_40_55;
  assign t_r39_c56_9 = t_r39_c56_5 + t_r39_c56_6;
  assign t_r39_c56_10 = t_r39_c56_7 + t_r39_c56_8;
  assign t_r39_c56_11 = t_r39_c56_9 + t_r39_c56_10;
  assign t_r39_c56_12 = t_r39_c56_11 + p_40_57;
  assign out_39_56 = t_r39_c56_12 >> 4;

  assign t_r39_c57_0 = p_38_57 << 1;
  assign t_r39_c57_1 = p_39_56 << 1;
  assign t_r39_c57_2 = p_39_57 << 2;
  assign t_r39_c57_3 = p_39_58 << 1;
  assign t_r39_c57_4 = p_40_57 << 1;
  assign t_r39_c57_5 = t_r39_c57_0 + p_38_56;
  assign t_r39_c57_6 = t_r39_c57_1 + p_38_58;
  assign t_r39_c57_7 = t_r39_c57_2 + t_r39_c57_3;
  assign t_r39_c57_8 = t_r39_c57_4 + p_40_56;
  assign t_r39_c57_9 = t_r39_c57_5 + t_r39_c57_6;
  assign t_r39_c57_10 = t_r39_c57_7 + t_r39_c57_8;
  assign t_r39_c57_11 = t_r39_c57_9 + t_r39_c57_10;
  assign t_r39_c57_12 = t_r39_c57_11 + p_40_58;
  assign out_39_57 = t_r39_c57_12 >> 4;

  assign t_r39_c58_0 = p_38_58 << 1;
  assign t_r39_c58_1 = p_39_57 << 1;
  assign t_r39_c58_2 = p_39_58 << 2;
  assign t_r39_c58_3 = p_39_59 << 1;
  assign t_r39_c58_4 = p_40_58 << 1;
  assign t_r39_c58_5 = t_r39_c58_0 + p_38_57;
  assign t_r39_c58_6 = t_r39_c58_1 + p_38_59;
  assign t_r39_c58_7 = t_r39_c58_2 + t_r39_c58_3;
  assign t_r39_c58_8 = t_r39_c58_4 + p_40_57;
  assign t_r39_c58_9 = t_r39_c58_5 + t_r39_c58_6;
  assign t_r39_c58_10 = t_r39_c58_7 + t_r39_c58_8;
  assign t_r39_c58_11 = t_r39_c58_9 + t_r39_c58_10;
  assign t_r39_c58_12 = t_r39_c58_11 + p_40_59;
  assign out_39_58 = t_r39_c58_12 >> 4;

  assign t_r39_c59_0 = p_38_59 << 1;
  assign t_r39_c59_1 = p_39_58 << 1;
  assign t_r39_c59_2 = p_39_59 << 2;
  assign t_r39_c59_3 = p_39_60 << 1;
  assign t_r39_c59_4 = p_40_59 << 1;
  assign t_r39_c59_5 = t_r39_c59_0 + p_38_58;
  assign t_r39_c59_6 = t_r39_c59_1 + p_38_60;
  assign t_r39_c59_7 = t_r39_c59_2 + t_r39_c59_3;
  assign t_r39_c59_8 = t_r39_c59_4 + p_40_58;
  assign t_r39_c59_9 = t_r39_c59_5 + t_r39_c59_6;
  assign t_r39_c59_10 = t_r39_c59_7 + t_r39_c59_8;
  assign t_r39_c59_11 = t_r39_c59_9 + t_r39_c59_10;
  assign t_r39_c59_12 = t_r39_c59_11 + p_40_60;
  assign out_39_59 = t_r39_c59_12 >> 4;

  assign t_r39_c60_0 = p_38_60 << 1;
  assign t_r39_c60_1 = p_39_59 << 1;
  assign t_r39_c60_2 = p_39_60 << 2;
  assign t_r39_c60_3 = p_39_61 << 1;
  assign t_r39_c60_4 = p_40_60 << 1;
  assign t_r39_c60_5 = t_r39_c60_0 + p_38_59;
  assign t_r39_c60_6 = t_r39_c60_1 + p_38_61;
  assign t_r39_c60_7 = t_r39_c60_2 + t_r39_c60_3;
  assign t_r39_c60_8 = t_r39_c60_4 + p_40_59;
  assign t_r39_c60_9 = t_r39_c60_5 + t_r39_c60_6;
  assign t_r39_c60_10 = t_r39_c60_7 + t_r39_c60_8;
  assign t_r39_c60_11 = t_r39_c60_9 + t_r39_c60_10;
  assign t_r39_c60_12 = t_r39_c60_11 + p_40_61;
  assign out_39_60 = t_r39_c60_12 >> 4;

  assign t_r39_c61_0 = p_38_61 << 1;
  assign t_r39_c61_1 = p_39_60 << 1;
  assign t_r39_c61_2 = p_39_61 << 2;
  assign t_r39_c61_3 = p_39_62 << 1;
  assign t_r39_c61_4 = p_40_61 << 1;
  assign t_r39_c61_5 = t_r39_c61_0 + p_38_60;
  assign t_r39_c61_6 = t_r39_c61_1 + p_38_62;
  assign t_r39_c61_7 = t_r39_c61_2 + t_r39_c61_3;
  assign t_r39_c61_8 = t_r39_c61_4 + p_40_60;
  assign t_r39_c61_9 = t_r39_c61_5 + t_r39_c61_6;
  assign t_r39_c61_10 = t_r39_c61_7 + t_r39_c61_8;
  assign t_r39_c61_11 = t_r39_c61_9 + t_r39_c61_10;
  assign t_r39_c61_12 = t_r39_c61_11 + p_40_62;
  assign out_39_61 = t_r39_c61_12 >> 4;

  assign t_r39_c62_0 = p_38_62 << 1;
  assign t_r39_c62_1 = p_39_61 << 1;
  assign t_r39_c62_2 = p_39_62 << 2;
  assign t_r39_c62_3 = p_39_63 << 1;
  assign t_r39_c62_4 = p_40_62 << 1;
  assign t_r39_c62_5 = t_r39_c62_0 + p_38_61;
  assign t_r39_c62_6 = t_r39_c62_1 + p_38_63;
  assign t_r39_c62_7 = t_r39_c62_2 + t_r39_c62_3;
  assign t_r39_c62_8 = t_r39_c62_4 + p_40_61;
  assign t_r39_c62_9 = t_r39_c62_5 + t_r39_c62_6;
  assign t_r39_c62_10 = t_r39_c62_7 + t_r39_c62_8;
  assign t_r39_c62_11 = t_r39_c62_9 + t_r39_c62_10;
  assign t_r39_c62_12 = t_r39_c62_11 + p_40_63;
  assign out_39_62 = t_r39_c62_12 >> 4;

  assign t_r39_c63_0 = p_38_63 << 1;
  assign t_r39_c63_1 = p_39_62 << 1;
  assign t_r39_c63_2 = p_39_63 << 2;
  assign t_r39_c63_3 = p_39_64 << 1;
  assign t_r39_c63_4 = p_40_63 << 1;
  assign t_r39_c63_5 = t_r39_c63_0 + p_38_62;
  assign t_r39_c63_6 = t_r39_c63_1 + p_38_64;
  assign t_r39_c63_7 = t_r39_c63_2 + t_r39_c63_3;
  assign t_r39_c63_8 = t_r39_c63_4 + p_40_62;
  assign t_r39_c63_9 = t_r39_c63_5 + t_r39_c63_6;
  assign t_r39_c63_10 = t_r39_c63_7 + t_r39_c63_8;
  assign t_r39_c63_11 = t_r39_c63_9 + t_r39_c63_10;
  assign t_r39_c63_12 = t_r39_c63_11 + p_40_64;
  assign out_39_63 = t_r39_c63_12 >> 4;

  assign t_r39_c64_0 = p_38_64 << 1;
  assign t_r39_c64_1 = p_39_63 << 1;
  assign t_r39_c64_2 = p_39_64 << 2;
  assign t_r39_c64_3 = p_39_65 << 1;
  assign t_r39_c64_4 = p_40_64 << 1;
  assign t_r39_c64_5 = t_r39_c64_0 + p_38_63;
  assign t_r39_c64_6 = t_r39_c64_1 + p_38_65;
  assign t_r39_c64_7 = t_r39_c64_2 + t_r39_c64_3;
  assign t_r39_c64_8 = t_r39_c64_4 + p_40_63;
  assign t_r39_c64_9 = t_r39_c64_5 + t_r39_c64_6;
  assign t_r39_c64_10 = t_r39_c64_7 + t_r39_c64_8;
  assign t_r39_c64_11 = t_r39_c64_9 + t_r39_c64_10;
  assign t_r39_c64_12 = t_r39_c64_11 + p_40_65;
  assign out_39_64 = t_r39_c64_12 >> 4;

  assign t_r40_c1_0 = p_39_1 << 1;
  assign t_r40_c1_1 = p_40_0 << 1;
  assign t_r40_c1_2 = p_40_1 << 2;
  assign t_r40_c1_3 = p_40_2 << 1;
  assign t_r40_c1_4 = p_41_1 << 1;
  assign t_r40_c1_5 = t_r40_c1_0 + p_39_0;
  assign t_r40_c1_6 = t_r40_c1_1 + p_39_2;
  assign t_r40_c1_7 = t_r40_c1_2 + t_r40_c1_3;
  assign t_r40_c1_8 = t_r40_c1_4 + p_41_0;
  assign t_r40_c1_9 = t_r40_c1_5 + t_r40_c1_6;
  assign t_r40_c1_10 = t_r40_c1_7 + t_r40_c1_8;
  assign t_r40_c1_11 = t_r40_c1_9 + t_r40_c1_10;
  assign t_r40_c1_12 = t_r40_c1_11 + p_41_2;
  assign out_40_1 = t_r40_c1_12 >> 4;

  assign t_r40_c2_0 = p_39_2 << 1;
  assign t_r40_c2_1 = p_40_1 << 1;
  assign t_r40_c2_2 = p_40_2 << 2;
  assign t_r40_c2_3 = p_40_3 << 1;
  assign t_r40_c2_4 = p_41_2 << 1;
  assign t_r40_c2_5 = t_r40_c2_0 + p_39_1;
  assign t_r40_c2_6 = t_r40_c2_1 + p_39_3;
  assign t_r40_c2_7 = t_r40_c2_2 + t_r40_c2_3;
  assign t_r40_c2_8 = t_r40_c2_4 + p_41_1;
  assign t_r40_c2_9 = t_r40_c2_5 + t_r40_c2_6;
  assign t_r40_c2_10 = t_r40_c2_7 + t_r40_c2_8;
  assign t_r40_c2_11 = t_r40_c2_9 + t_r40_c2_10;
  assign t_r40_c2_12 = t_r40_c2_11 + p_41_3;
  assign out_40_2 = t_r40_c2_12 >> 4;

  assign t_r40_c3_0 = p_39_3 << 1;
  assign t_r40_c3_1 = p_40_2 << 1;
  assign t_r40_c3_2 = p_40_3 << 2;
  assign t_r40_c3_3 = p_40_4 << 1;
  assign t_r40_c3_4 = p_41_3 << 1;
  assign t_r40_c3_5 = t_r40_c3_0 + p_39_2;
  assign t_r40_c3_6 = t_r40_c3_1 + p_39_4;
  assign t_r40_c3_7 = t_r40_c3_2 + t_r40_c3_3;
  assign t_r40_c3_8 = t_r40_c3_4 + p_41_2;
  assign t_r40_c3_9 = t_r40_c3_5 + t_r40_c3_6;
  assign t_r40_c3_10 = t_r40_c3_7 + t_r40_c3_8;
  assign t_r40_c3_11 = t_r40_c3_9 + t_r40_c3_10;
  assign t_r40_c3_12 = t_r40_c3_11 + p_41_4;
  assign out_40_3 = t_r40_c3_12 >> 4;

  assign t_r40_c4_0 = p_39_4 << 1;
  assign t_r40_c4_1 = p_40_3 << 1;
  assign t_r40_c4_2 = p_40_4 << 2;
  assign t_r40_c4_3 = p_40_5 << 1;
  assign t_r40_c4_4 = p_41_4 << 1;
  assign t_r40_c4_5 = t_r40_c4_0 + p_39_3;
  assign t_r40_c4_6 = t_r40_c4_1 + p_39_5;
  assign t_r40_c4_7 = t_r40_c4_2 + t_r40_c4_3;
  assign t_r40_c4_8 = t_r40_c4_4 + p_41_3;
  assign t_r40_c4_9 = t_r40_c4_5 + t_r40_c4_6;
  assign t_r40_c4_10 = t_r40_c4_7 + t_r40_c4_8;
  assign t_r40_c4_11 = t_r40_c4_9 + t_r40_c4_10;
  assign t_r40_c4_12 = t_r40_c4_11 + p_41_5;
  assign out_40_4 = t_r40_c4_12 >> 4;

  assign t_r40_c5_0 = p_39_5 << 1;
  assign t_r40_c5_1 = p_40_4 << 1;
  assign t_r40_c5_2 = p_40_5 << 2;
  assign t_r40_c5_3 = p_40_6 << 1;
  assign t_r40_c5_4 = p_41_5 << 1;
  assign t_r40_c5_5 = t_r40_c5_0 + p_39_4;
  assign t_r40_c5_6 = t_r40_c5_1 + p_39_6;
  assign t_r40_c5_7 = t_r40_c5_2 + t_r40_c5_3;
  assign t_r40_c5_8 = t_r40_c5_4 + p_41_4;
  assign t_r40_c5_9 = t_r40_c5_5 + t_r40_c5_6;
  assign t_r40_c5_10 = t_r40_c5_7 + t_r40_c5_8;
  assign t_r40_c5_11 = t_r40_c5_9 + t_r40_c5_10;
  assign t_r40_c5_12 = t_r40_c5_11 + p_41_6;
  assign out_40_5 = t_r40_c5_12 >> 4;

  assign t_r40_c6_0 = p_39_6 << 1;
  assign t_r40_c6_1 = p_40_5 << 1;
  assign t_r40_c6_2 = p_40_6 << 2;
  assign t_r40_c6_3 = p_40_7 << 1;
  assign t_r40_c6_4 = p_41_6 << 1;
  assign t_r40_c6_5 = t_r40_c6_0 + p_39_5;
  assign t_r40_c6_6 = t_r40_c6_1 + p_39_7;
  assign t_r40_c6_7 = t_r40_c6_2 + t_r40_c6_3;
  assign t_r40_c6_8 = t_r40_c6_4 + p_41_5;
  assign t_r40_c6_9 = t_r40_c6_5 + t_r40_c6_6;
  assign t_r40_c6_10 = t_r40_c6_7 + t_r40_c6_8;
  assign t_r40_c6_11 = t_r40_c6_9 + t_r40_c6_10;
  assign t_r40_c6_12 = t_r40_c6_11 + p_41_7;
  assign out_40_6 = t_r40_c6_12 >> 4;

  assign t_r40_c7_0 = p_39_7 << 1;
  assign t_r40_c7_1 = p_40_6 << 1;
  assign t_r40_c7_2 = p_40_7 << 2;
  assign t_r40_c7_3 = p_40_8 << 1;
  assign t_r40_c7_4 = p_41_7 << 1;
  assign t_r40_c7_5 = t_r40_c7_0 + p_39_6;
  assign t_r40_c7_6 = t_r40_c7_1 + p_39_8;
  assign t_r40_c7_7 = t_r40_c7_2 + t_r40_c7_3;
  assign t_r40_c7_8 = t_r40_c7_4 + p_41_6;
  assign t_r40_c7_9 = t_r40_c7_5 + t_r40_c7_6;
  assign t_r40_c7_10 = t_r40_c7_7 + t_r40_c7_8;
  assign t_r40_c7_11 = t_r40_c7_9 + t_r40_c7_10;
  assign t_r40_c7_12 = t_r40_c7_11 + p_41_8;
  assign out_40_7 = t_r40_c7_12 >> 4;

  assign t_r40_c8_0 = p_39_8 << 1;
  assign t_r40_c8_1 = p_40_7 << 1;
  assign t_r40_c8_2 = p_40_8 << 2;
  assign t_r40_c8_3 = p_40_9 << 1;
  assign t_r40_c8_4 = p_41_8 << 1;
  assign t_r40_c8_5 = t_r40_c8_0 + p_39_7;
  assign t_r40_c8_6 = t_r40_c8_1 + p_39_9;
  assign t_r40_c8_7 = t_r40_c8_2 + t_r40_c8_3;
  assign t_r40_c8_8 = t_r40_c8_4 + p_41_7;
  assign t_r40_c8_9 = t_r40_c8_5 + t_r40_c8_6;
  assign t_r40_c8_10 = t_r40_c8_7 + t_r40_c8_8;
  assign t_r40_c8_11 = t_r40_c8_9 + t_r40_c8_10;
  assign t_r40_c8_12 = t_r40_c8_11 + p_41_9;
  assign out_40_8 = t_r40_c8_12 >> 4;

  assign t_r40_c9_0 = p_39_9 << 1;
  assign t_r40_c9_1 = p_40_8 << 1;
  assign t_r40_c9_2 = p_40_9 << 2;
  assign t_r40_c9_3 = p_40_10 << 1;
  assign t_r40_c9_4 = p_41_9 << 1;
  assign t_r40_c9_5 = t_r40_c9_0 + p_39_8;
  assign t_r40_c9_6 = t_r40_c9_1 + p_39_10;
  assign t_r40_c9_7 = t_r40_c9_2 + t_r40_c9_3;
  assign t_r40_c9_8 = t_r40_c9_4 + p_41_8;
  assign t_r40_c9_9 = t_r40_c9_5 + t_r40_c9_6;
  assign t_r40_c9_10 = t_r40_c9_7 + t_r40_c9_8;
  assign t_r40_c9_11 = t_r40_c9_9 + t_r40_c9_10;
  assign t_r40_c9_12 = t_r40_c9_11 + p_41_10;
  assign out_40_9 = t_r40_c9_12 >> 4;

  assign t_r40_c10_0 = p_39_10 << 1;
  assign t_r40_c10_1 = p_40_9 << 1;
  assign t_r40_c10_2 = p_40_10 << 2;
  assign t_r40_c10_3 = p_40_11 << 1;
  assign t_r40_c10_4 = p_41_10 << 1;
  assign t_r40_c10_5 = t_r40_c10_0 + p_39_9;
  assign t_r40_c10_6 = t_r40_c10_1 + p_39_11;
  assign t_r40_c10_7 = t_r40_c10_2 + t_r40_c10_3;
  assign t_r40_c10_8 = t_r40_c10_4 + p_41_9;
  assign t_r40_c10_9 = t_r40_c10_5 + t_r40_c10_6;
  assign t_r40_c10_10 = t_r40_c10_7 + t_r40_c10_8;
  assign t_r40_c10_11 = t_r40_c10_9 + t_r40_c10_10;
  assign t_r40_c10_12 = t_r40_c10_11 + p_41_11;
  assign out_40_10 = t_r40_c10_12 >> 4;

  assign t_r40_c11_0 = p_39_11 << 1;
  assign t_r40_c11_1 = p_40_10 << 1;
  assign t_r40_c11_2 = p_40_11 << 2;
  assign t_r40_c11_3 = p_40_12 << 1;
  assign t_r40_c11_4 = p_41_11 << 1;
  assign t_r40_c11_5 = t_r40_c11_0 + p_39_10;
  assign t_r40_c11_6 = t_r40_c11_1 + p_39_12;
  assign t_r40_c11_7 = t_r40_c11_2 + t_r40_c11_3;
  assign t_r40_c11_8 = t_r40_c11_4 + p_41_10;
  assign t_r40_c11_9 = t_r40_c11_5 + t_r40_c11_6;
  assign t_r40_c11_10 = t_r40_c11_7 + t_r40_c11_8;
  assign t_r40_c11_11 = t_r40_c11_9 + t_r40_c11_10;
  assign t_r40_c11_12 = t_r40_c11_11 + p_41_12;
  assign out_40_11 = t_r40_c11_12 >> 4;

  assign t_r40_c12_0 = p_39_12 << 1;
  assign t_r40_c12_1 = p_40_11 << 1;
  assign t_r40_c12_2 = p_40_12 << 2;
  assign t_r40_c12_3 = p_40_13 << 1;
  assign t_r40_c12_4 = p_41_12 << 1;
  assign t_r40_c12_5 = t_r40_c12_0 + p_39_11;
  assign t_r40_c12_6 = t_r40_c12_1 + p_39_13;
  assign t_r40_c12_7 = t_r40_c12_2 + t_r40_c12_3;
  assign t_r40_c12_8 = t_r40_c12_4 + p_41_11;
  assign t_r40_c12_9 = t_r40_c12_5 + t_r40_c12_6;
  assign t_r40_c12_10 = t_r40_c12_7 + t_r40_c12_8;
  assign t_r40_c12_11 = t_r40_c12_9 + t_r40_c12_10;
  assign t_r40_c12_12 = t_r40_c12_11 + p_41_13;
  assign out_40_12 = t_r40_c12_12 >> 4;

  assign t_r40_c13_0 = p_39_13 << 1;
  assign t_r40_c13_1 = p_40_12 << 1;
  assign t_r40_c13_2 = p_40_13 << 2;
  assign t_r40_c13_3 = p_40_14 << 1;
  assign t_r40_c13_4 = p_41_13 << 1;
  assign t_r40_c13_5 = t_r40_c13_0 + p_39_12;
  assign t_r40_c13_6 = t_r40_c13_1 + p_39_14;
  assign t_r40_c13_7 = t_r40_c13_2 + t_r40_c13_3;
  assign t_r40_c13_8 = t_r40_c13_4 + p_41_12;
  assign t_r40_c13_9 = t_r40_c13_5 + t_r40_c13_6;
  assign t_r40_c13_10 = t_r40_c13_7 + t_r40_c13_8;
  assign t_r40_c13_11 = t_r40_c13_9 + t_r40_c13_10;
  assign t_r40_c13_12 = t_r40_c13_11 + p_41_14;
  assign out_40_13 = t_r40_c13_12 >> 4;

  assign t_r40_c14_0 = p_39_14 << 1;
  assign t_r40_c14_1 = p_40_13 << 1;
  assign t_r40_c14_2 = p_40_14 << 2;
  assign t_r40_c14_3 = p_40_15 << 1;
  assign t_r40_c14_4 = p_41_14 << 1;
  assign t_r40_c14_5 = t_r40_c14_0 + p_39_13;
  assign t_r40_c14_6 = t_r40_c14_1 + p_39_15;
  assign t_r40_c14_7 = t_r40_c14_2 + t_r40_c14_3;
  assign t_r40_c14_8 = t_r40_c14_4 + p_41_13;
  assign t_r40_c14_9 = t_r40_c14_5 + t_r40_c14_6;
  assign t_r40_c14_10 = t_r40_c14_7 + t_r40_c14_8;
  assign t_r40_c14_11 = t_r40_c14_9 + t_r40_c14_10;
  assign t_r40_c14_12 = t_r40_c14_11 + p_41_15;
  assign out_40_14 = t_r40_c14_12 >> 4;

  assign t_r40_c15_0 = p_39_15 << 1;
  assign t_r40_c15_1 = p_40_14 << 1;
  assign t_r40_c15_2 = p_40_15 << 2;
  assign t_r40_c15_3 = p_40_16 << 1;
  assign t_r40_c15_4 = p_41_15 << 1;
  assign t_r40_c15_5 = t_r40_c15_0 + p_39_14;
  assign t_r40_c15_6 = t_r40_c15_1 + p_39_16;
  assign t_r40_c15_7 = t_r40_c15_2 + t_r40_c15_3;
  assign t_r40_c15_8 = t_r40_c15_4 + p_41_14;
  assign t_r40_c15_9 = t_r40_c15_5 + t_r40_c15_6;
  assign t_r40_c15_10 = t_r40_c15_7 + t_r40_c15_8;
  assign t_r40_c15_11 = t_r40_c15_9 + t_r40_c15_10;
  assign t_r40_c15_12 = t_r40_c15_11 + p_41_16;
  assign out_40_15 = t_r40_c15_12 >> 4;

  assign t_r40_c16_0 = p_39_16 << 1;
  assign t_r40_c16_1 = p_40_15 << 1;
  assign t_r40_c16_2 = p_40_16 << 2;
  assign t_r40_c16_3 = p_40_17 << 1;
  assign t_r40_c16_4 = p_41_16 << 1;
  assign t_r40_c16_5 = t_r40_c16_0 + p_39_15;
  assign t_r40_c16_6 = t_r40_c16_1 + p_39_17;
  assign t_r40_c16_7 = t_r40_c16_2 + t_r40_c16_3;
  assign t_r40_c16_8 = t_r40_c16_4 + p_41_15;
  assign t_r40_c16_9 = t_r40_c16_5 + t_r40_c16_6;
  assign t_r40_c16_10 = t_r40_c16_7 + t_r40_c16_8;
  assign t_r40_c16_11 = t_r40_c16_9 + t_r40_c16_10;
  assign t_r40_c16_12 = t_r40_c16_11 + p_41_17;
  assign out_40_16 = t_r40_c16_12 >> 4;

  assign t_r40_c17_0 = p_39_17 << 1;
  assign t_r40_c17_1 = p_40_16 << 1;
  assign t_r40_c17_2 = p_40_17 << 2;
  assign t_r40_c17_3 = p_40_18 << 1;
  assign t_r40_c17_4 = p_41_17 << 1;
  assign t_r40_c17_5 = t_r40_c17_0 + p_39_16;
  assign t_r40_c17_6 = t_r40_c17_1 + p_39_18;
  assign t_r40_c17_7 = t_r40_c17_2 + t_r40_c17_3;
  assign t_r40_c17_8 = t_r40_c17_4 + p_41_16;
  assign t_r40_c17_9 = t_r40_c17_5 + t_r40_c17_6;
  assign t_r40_c17_10 = t_r40_c17_7 + t_r40_c17_8;
  assign t_r40_c17_11 = t_r40_c17_9 + t_r40_c17_10;
  assign t_r40_c17_12 = t_r40_c17_11 + p_41_18;
  assign out_40_17 = t_r40_c17_12 >> 4;

  assign t_r40_c18_0 = p_39_18 << 1;
  assign t_r40_c18_1 = p_40_17 << 1;
  assign t_r40_c18_2 = p_40_18 << 2;
  assign t_r40_c18_3 = p_40_19 << 1;
  assign t_r40_c18_4 = p_41_18 << 1;
  assign t_r40_c18_5 = t_r40_c18_0 + p_39_17;
  assign t_r40_c18_6 = t_r40_c18_1 + p_39_19;
  assign t_r40_c18_7 = t_r40_c18_2 + t_r40_c18_3;
  assign t_r40_c18_8 = t_r40_c18_4 + p_41_17;
  assign t_r40_c18_9 = t_r40_c18_5 + t_r40_c18_6;
  assign t_r40_c18_10 = t_r40_c18_7 + t_r40_c18_8;
  assign t_r40_c18_11 = t_r40_c18_9 + t_r40_c18_10;
  assign t_r40_c18_12 = t_r40_c18_11 + p_41_19;
  assign out_40_18 = t_r40_c18_12 >> 4;

  assign t_r40_c19_0 = p_39_19 << 1;
  assign t_r40_c19_1 = p_40_18 << 1;
  assign t_r40_c19_2 = p_40_19 << 2;
  assign t_r40_c19_3 = p_40_20 << 1;
  assign t_r40_c19_4 = p_41_19 << 1;
  assign t_r40_c19_5 = t_r40_c19_0 + p_39_18;
  assign t_r40_c19_6 = t_r40_c19_1 + p_39_20;
  assign t_r40_c19_7 = t_r40_c19_2 + t_r40_c19_3;
  assign t_r40_c19_8 = t_r40_c19_4 + p_41_18;
  assign t_r40_c19_9 = t_r40_c19_5 + t_r40_c19_6;
  assign t_r40_c19_10 = t_r40_c19_7 + t_r40_c19_8;
  assign t_r40_c19_11 = t_r40_c19_9 + t_r40_c19_10;
  assign t_r40_c19_12 = t_r40_c19_11 + p_41_20;
  assign out_40_19 = t_r40_c19_12 >> 4;

  assign t_r40_c20_0 = p_39_20 << 1;
  assign t_r40_c20_1 = p_40_19 << 1;
  assign t_r40_c20_2 = p_40_20 << 2;
  assign t_r40_c20_3 = p_40_21 << 1;
  assign t_r40_c20_4 = p_41_20 << 1;
  assign t_r40_c20_5 = t_r40_c20_0 + p_39_19;
  assign t_r40_c20_6 = t_r40_c20_1 + p_39_21;
  assign t_r40_c20_7 = t_r40_c20_2 + t_r40_c20_3;
  assign t_r40_c20_8 = t_r40_c20_4 + p_41_19;
  assign t_r40_c20_9 = t_r40_c20_5 + t_r40_c20_6;
  assign t_r40_c20_10 = t_r40_c20_7 + t_r40_c20_8;
  assign t_r40_c20_11 = t_r40_c20_9 + t_r40_c20_10;
  assign t_r40_c20_12 = t_r40_c20_11 + p_41_21;
  assign out_40_20 = t_r40_c20_12 >> 4;

  assign t_r40_c21_0 = p_39_21 << 1;
  assign t_r40_c21_1 = p_40_20 << 1;
  assign t_r40_c21_2 = p_40_21 << 2;
  assign t_r40_c21_3 = p_40_22 << 1;
  assign t_r40_c21_4 = p_41_21 << 1;
  assign t_r40_c21_5 = t_r40_c21_0 + p_39_20;
  assign t_r40_c21_6 = t_r40_c21_1 + p_39_22;
  assign t_r40_c21_7 = t_r40_c21_2 + t_r40_c21_3;
  assign t_r40_c21_8 = t_r40_c21_4 + p_41_20;
  assign t_r40_c21_9 = t_r40_c21_5 + t_r40_c21_6;
  assign t_r40_c21_10 = t_r40_c21_7 + t_r40_c21_8;
  assign t_r40_c21_11 = t_r40_c21_9 + t_r40_c21_10;
  assign t_r40_c21_12 = t_r40_c21_11 + p_41_22;
  assign out_40_21 = t_r40_c21_12 >> 4;

  assign t_r40_c22_0 = p_39_22 << 1;
  assign t_r40_c22_1 = p_40_21 << 1;
  assign t_r40_c22_2 = p_40_22 << 2;
  assign t_r40_c22_3 = p_40_23 << 1;
  assign t_r40_c22_4 = p_41_22 << 1;
  assign t_r40_c22_5 = t_r40_c22_0 + p_39_21;
  assign t_r40_c22_6 = t_r40_c22_1 + p_39_23;
  assign t_r40_c22_7 = t_r40_c22_2 + t_r40_c22_3;
  assign t_r40_c22_8 = t_r40_c22_4 + p_41_21;
  assign t_r40_c22_9 = t_r40_c22_5 + t_r40_c22_6;
  assign t_r40_c22_10 = t_r40_c22_7 + t_r40_c22_8;
  assign t_r40_c22_11 = t_r40_c22_9 + t_r40_c22_10;
  assign t_r40_c22_12 = t_r40_c22_11 + p_41_23;
  assign out_40_22 = t_r40_c22_12 >> 4;

  assign t_r40_c23_0 = p_39_23 << 1;
  assign t_r40_c23_1 = p_40_22 << 1;
  assign t_r40_c23_2 = p_40_23 << 2;
  assign t_r40_c23_3 = p_40_24 << 1;
  assign t_r40_c23_4 = p_41_23 << 1;
  assign t_r40_c23_5 = t_r40_c23_0 + p_39_22;
  assign t_r40_c23_6 = t_r40_c23_1 + p_39_24;
  assign t_r40_c23_7 = t_r40_c23_2 + t_r40_c23_3;
  assign t_r40_c23_8 = t_r40_c23_4 + p_41_22;
  assign t_r40_c23_9 = t_r40_c23_5 + t_r40_c23_6;
  assign t_r40_c23_10 = t_r40_c23_7 + t_r40_c23_8;
  assign t_r40_c23_11 = t_r40_c23_9 + t_r40_c23_10;
  assign t_r40_c23_12 = t_r40_c23_11 + p_41_24;
  assign out_40_23 = t_r40_c23_12 >> 4;

  assign t_r40_c24_0 = p_39_24 << 1;
  assign t_r40_c24_1 = p_40_23 << 1;
  assign t_r40_c24_2 = p_40_24 << 2;
  assign t_r40_c24_3 = p_40_25 << 1;
  assign t_r40_c24_4 = p_41_24 << 1;
  assign t_r40_c24_5 = t_r40_c24_0 + p_39_23;
  assign t_r40_c24_6 = t_r40_c24_1 + p_39_25;
  assign t_r40_c24_7 = t_r40_c24_2 + t_r40_c24_3;
  assign t_r40_c24_8 = t_r40_c24_4 + p_41_23;
  assign t_r40_c24_9 = t_r40_c24_5 + t_r40_c24_6;
  assign t_r40_c24_10 = t_r40_c24_7 + t_r40_c24_8;
  assign t_r40_c24_11 = t_r40_c24_9 + t_r40_c24_10;
  assign t_r40_c24_12 = t_r40_c24_11 + p_41_25;
  assign out_40_24 = t_r40_c24_12 >> 4;

  assign t_r40_c25_0 = p_39_25 << 1;
  assign t_r40_c25_1 = p_40_24 << 1;
  assign t_r40_c25_2 = p_40_25 << 2;
  assign t_r40_c25_3 = p_40_26 << 1;
  assign t_r40_c25_4 = p_41_25 << 1;
  assign t_r40_c25_5 = t_r40_c25_0 + p_39_24;
  assign t_r40_c25_6 = t_r40_c25_1 + p_39_26;
  assign t_r40_c25_7 = t_r40_c25_2 + t_r40_c25_3;
  assign t_r40_c25_8 = t_r40_c25_4 + p_41_24;
  assign t_r40_c25_9 = t_r40_c25_5 + t_r40_c25_6;
  assign t_r40_c25_10 = t_r40_c25_7 + t_r40_c25_8;
  assign t_r40_c25_11 = t_r40_c25_9 + t_r40_c25_10;
  assign t_r40_c25_12 = t_r40_c25_11 + p_41_26;
  assign out_40_25 = t_r40_c25_12 >> 4;

  assign t_r40_c26_0 = p_39_26 << 1;
  assign t_r40_c26_1 = p_40_25 << 1;
  assign t_r40_c26_2 = p_40_26 << 2;
  assign t_r40_c26_3 = p_40_27 << 1;
  assign t_r40_c26_4 = p_41_26 << 1;
  assign t_r40_c26_5 = t_r40_c26_0 + p_39_25;
  assign t_r40_c26_6 = t_r40_c26_1 + p_39_27;
  assign t_r40_c26_7 = t_r40_c26_2 + t_r40_c26_3;
  assign t_r40_c26_8 = t_r40_c26_4 + p_41_25;
  assign t_r40_c26_9 = t_r40_c26_5 + t_r40_c26_6;
  assign t_r40_c26_10 = t_r40_c26_7 + t_r40_c26_8;
  assign t_r40_c26_11 = t_r40_c26_9 + t_r40_c26_10;
  assign t_r40_c26_12 = t_r40_c26_11 + p_41_27;
  assign out_40_26 = t_r40_c26_12 >> 4;

  assign t_r40_c27_0 = p_39_27 << 1;
  assign t_r40_c27_1 = p_40_26 << 1;
  assign t_r40_c27_2 = p_40_27 << 2;
  assign t_r40_c27_3 = p_40_28 << 1;
  assign t_r40_c27_4 = p_41_27 << 1;
  assign t_r40_c27_5 = t_r40_c27_0 + p_39_26;
  assign t_r40_c27_6 = t_r40_c27_1 + p_39_28;
  assign t_r40_c27_7 = t_r40_c27_2 + t_r40_c27_3;
  assign t_r40_c27_8 = t_r40_c27_4 + p_41_26;
  assign t_r40_c27_9 = t_r40_c27_5 + t_r40_c27_6;
  assign t_r40_c27_10 = t_r40_c27_7 + t_r40_c27_8;
  assign t_r40_c27_11 = t_r40_c27_9 + t_r40_c27_10;
  assign t_r40_c27_12 = t_r40_c27_11 + p_41_28;
  assign out_40_27 = t_r40_c27_12 >> 4;

  assign t_r40_c28_0 = p_39_28 << 1;
  assign t_r40_c28_1 = p_40_27 << 1;
  assign t_r40_c28_2 = p_40_28 << 2;
  assign t_r40_c28_3 = p_40_29 << 1;
  assign t_r40_c28_4 = p_41_28 << 1;
  assign t_r40_c28_5 = t_r40_c28_0 + p_39_27;
  assign t_r40_c28_6 = t_r40_c28_1 + p_39_29;
  assign t_r40_c28_7 = t_r40_c28_2 + t_r40_c28_3;
  assign t_r40_c28_8 = t_r40_c28_4 + p_41_27;
  assign t_r40_c28_9 = t_r40_c28_5 + t_r40_c28_6;
  assign t_r40_c28_10 = t_r40_c28_7 + t_r40_c28_8;
  assign t_r40_c28_11 = t_r40_c28_9 + t_r40_c28_10;
  assign t_r40_c28_12 = t_r40_c28_11 + p_41_29;
  assign out_40_28 = t_r40_c28_12 >> 4;

  assign t_r40_c29_0 = p_39_29 << 1;
  assign t_r40_c29_1 = p_40_28 << 1;
  assign t_r40_c29_2 = p_40_29 << 2;
  assign t_r40_c29_3 = p_40_30 << 1;
  assign t_r40_c29_4 = p_41_29 << 1;
  assign t_r40_c29_5 = t_r40_c29_0 + p_39_28;
  assign t_r40_c29_6 = t_r40_c29_1 + p_39_30;
  assign t_r40_c29_7 = t_r40_c29_2 + t_r40_c29_3;
  assign t_r40_c29_8 = t_r40_c29_4 + p_41_28;
  assign t_r40_c29_9 = t_r40_c29_5 + t_r40_c29_6;
  assign t_r40_c29_10 = t_r40_c29_7 + t_r40_c29_8;
  assign t_r40_c29_11 = t_r40_c29_9 + t_r40_c29_10;
  assign t_r40_c29_12 = t_r40_c29_11 + p_41_30;
  assign out_40_29 = t_r40_c29_12 >> 4;

  assign t_r40_c30_0 = p_39_30 << 1;
  assign t_r40_c30_1 = p_40_29 << 1;
  assign t_r40_c30_2 = p_40_30 << 2;
  assign t_r40_c30_3 = p_40_31 << 1;
  assign t_r40_c30_4 = p_41_30 << 1;
  assign t_r40_c30_5 = t_r40_c30_0 + p_39_29;
  assign t_r40_c30_6 = t_r40_c30_1 + p_39_31;
  assign t_r40_c30_7 = t_r40_c30_2 + t_r40_c30_3;
  assign t_r40_c30_8 = t_r40_c30_4 + p_41_29;
  assign t_r40_c30_9 = t_r40_c30_5 + t_r40_c30_6;
  assign t_r40_c30_10 = t_r40_c30_7 + t_r40_c30_8;
  assign t_r40_c30_11 = t_r40_c30_9 + t_r40_c30_10;
  assign t_r40_c30_12 = t_r40_c30_11 + p_41_31;
  assign out_40_30 = t_r40_c30_12 >> 4;

  assign t_r40_c31_0 = p_39_31 << 1;
  assign t_r40_c31_1 = p_40_30 << 1;
  assign t_r40_c31_2 = p_40_31 << 2;
  assign t_r40_c31_3 = p_40_32 << 1;
  assign t_r40_c31_4 = p_41_31 << 1;
  assign t_r40_c31_5 = t_r40_c31_0 + p_39_30;
  assign t_r40_c31_6 = t_r40_c31_1 + p_39_32;
  assign t_r40_c31_7 = t_r40_c31_2 + t_r40_c31_3;
  assign t_r40_c31_8 = t_r40_c31_4 + p_41_30;
  assign t_r40_c31_9 = t_r40_c31_5 + t_r40_c31_6;
  assign t_r40_c31_10 = t_r40_c31_7 + t_r40_c31_8;
  assign t_r40_c31_11 = t_r40_c31_9 + t_r40_c31_10;
  assign t_r40_c31_12 = t_r40_c31_11 + p_41_32;
  assign out_40_31 = t_r40_c31_12 >> 4;

  assign t_r40_c32_0 = p_39_32 << 1;
  assign t_r40_c32_1 = p_40_31 << 1;
  assign t_r40_c32_2 = p_40_32 << 2;
  assign t_r40_c32_3 = p_40_33 << 1;
  assign t_r40_c32_4 = p_41_32 << 1;
  assign t_r40_c32_5 = t_r40_c32_0 + p_39_31;
  assign t_r40_c32_6 = t_r40_c32_1 + p_39_33;
  assign t_r40_c32_7 = t_r40_c32_2 + t_r40_c32_3;
  assign t_r40_c32_8 = t_r40_c32_4 + p_41_31;
  assign t_r40_c32_9 = t_r40_c32_5 + t_r40_c32_6;
  assign t_r40_c32_10 = t_r40_c32_7 + t_r40_c32_8;
  assign t_r40_c32_11 = t_r40_c32_9 + t_r40_c32_10;
  assign t_r40_c32_12 = t_r40_c32_11 + p_41_33;
  assign out_40_32 = t_r40_c32_12 >> 4;

  assign t_r40_c33_0 = p_39_33 << 1;
  assign t_r40_c33_1 = p_40_32 << 1;
  assign t_r40_c33_2 = p_40_33 << 2;
  assign t_r40_c33_3 = p_40_34 << 1;
  assign t_r40_c33_4 = p_41_33 << 1;
  assign t_r40_c33_5 = t_r40_c33_0 + p_39_32;
  assign t_r40_c33_6 = t_r40_c33_1 + p_39_34;
  assign t_r40_c33_7 = t_r40_c33_2 + t_r40_c33_3;
  assign t_r40_c33_8 = t_r40_c33_4 + p_41_32;
  assign t_r40_c33_9 = t_r40_c33_5 + t_r40_c33_6;
  assign t_r40_c33_10 = t_r40_c33_7 + t_r40_c33_8;
  assign t_r40_c33_11 = t_r40_c33_9 + t_r40_c33_10;
  assign t_r40_c33_12 = t_r40_c33_11 + p_41_34;
  assign out_40_33 = t_r40_c33_12 >> 4;

  assign t_r40_c34_0 = p_39_34 << 1;
  assign t_r40_c34_1 = p_40_33 << 1;
  assign t_r40_c34_2 = p_40_34 << 2;
  assign t_r40_c34_3 = p_40_35 << 1;
  assign t_r40_c34_4 = p_41_34 << 1;
  assign t_r40_c34_5 = t_r40_c34_0 + p_39_33;
  assign t_r40_c34_6 = t_r40_c34_1 + p_39_35;
  assign t_r40_c34_7 = t_r40_c34_2 + t_r40_c34_3;
  assign t_r40_c34_8 = t_r40_c34_4 + p_41_33;
  assign t_r40_c34_9 = t_r40_c34_5 + t_r40_c34_6;
  assign t_r40_c34_10 = t_r40_c34_7 + t_r40_c34_8;
  assign t_r40_c34_11 = t_r40_c34_9 + t_r40_c34_10;
  assign t_r40_c34_12 = t_r40_c34_11 + p_41_35;
  assign out_40_34 = t_r40_c34_12 >> 4;

  assign t_r40_c35_0 = p_39_35 << 1;
  assign t_r40_c35_1 = p_40_34 << 1;
  assign t_r40_c35_2 = p_40_35 << 2;
  assign t_r40_c35_3 = p_40_36 << 1;
  assign t_r40_c35_4 = p_41_35 << 1;
  assign t_r40_c35_5 = t_r40_c35_0 + p_39_34;
  assign t_r40_c35_6 = t_r40_c35_1 + p_39_36;
  assign t_r40_c35_7 = t_r40_c35_2 + t_r40_c35_3;
  assign t_r40_c35_8 = t_r40_c35_4 + p_41_34;
  assign t_r40_c35_9 = t_r40_c35_5 + t_r40_c35_6;
  assign t_r40_c35_10 = t_r40_c35_7 + t_r40_c35_8;
  assign t_r40_c35_11 = t_r40_c35_9 + t_r40_c35_10;
  assign t_r40_c35_12 = t_r40_c35_11 + p_41_36;
  assign out_40_35 = t_r40_c35_12 >> 4;

  assign t_r40_c36_0 = p_39_36 << 1;
  assign t_r40_c36_1 = p_40_35 << 1;
  assign t_r40_c36_2 = p_40_36 << 2;
  assign t_r40_c36_3 = p_40_37 << 1;
  assign t_r40_c36_4 = p_41_36 << 1;
  assign t_r40_c36_5 = t_r40_c36_0 + p_39_35;
  assign t_r40_c36_6 = t_r40_c36_1 + p_39_37;
  assign t_r40_c36_7 = t_r40_c36_2 + t_r40_c36_3;
  assign t_r40_c36_8 = t_r40_c36_4 + p_41_35;
  assign t_r40_c36_9 = t_r40_c36_5 + t_r40_c36_6;
  assign t_r40_c36_10 = t_r40_c36_7 + t_r40_c36_8;
  assign t_r40_c36_11 = t_r40_c36_9 + t_r40_c36_10;
  assign t_r40_c36_12 = t_r40_c36_11 + p_41_37;
  assign out_40_36 = t_r40_c36_12 >> 4;

  assign t_r40_c37_0 = p_39_37 << 1;
  assign t_r40_c37_1 = p_40_36 << 1;
  assign t_r40_c37_2 = p_40_37 << 2;
  assign t_r40_c37_3 = p_40_38 << 1;
  assign t_r40_c37_4 = p_41_37 << 1;
  assign t_r40_c37_5 = t_r40_c37_0 + p_39_36;
  assign t_r40_c37_6 = t_r40_c37_1 + p_39_38;
  assign t_r40_c37_7 = t_r40_c37_2 + t_r40_c37_3;
  assign t_r40_c37_8 = t_r40_c37_4 + p_41_36;
  assign t_r40_c37_9 = t_r40_c37_5 + t_r40_c37_6;
  assign t_r40_c37_10 = t_r40_c37_7 + t_r40_c37_8;
  assign t_r40_c37_11 = t_r40_c37_9 + t_r40_c37_10;
  assign t_r40_c37_12 = t_r40_c37_11 + p_41_38;
  assign out_40_37 = t_r40_c37_12 >> 4;

  assign t_r40_c38_0 = p_39_38 << 1;
  assign t_r40_c38_1 = p_40_37 << 1;
  assign t_r40_c38_2 = p_40_38 << 2;
  assign t_r40_c38_3 = p_40_39 << 1;
  assign t_r40_c38_4 = p_41_38 << 1;
  assign t_r40_c38_5 = t_r40_c38_0 + p_39_37;
  assign t_r40_c38_6 = t_r40_c38_1 + p_39_39;
  assign t_r40_c38_7 = t_r40_c38_2 + t_r40_c38_3;
  assign t_r40_c38_8 = t_r40_c38_4 + p_41_37;
  assign t_r40_c38_9 = t_r40_c38_5 + t_r40_c38_6;
  assign t_r40_c38_10 = t_r40_c38_7 + t_r40_c38_8;
  assign t_r40_c38_11 = t_r40_c38_9 + t_r40_c38_10;
  assign t_r40_c38_12 = t_r40_c38_11 + p_41_39;
  assign out_40_38 = t_r40_c38_12 >> 4;

  assign t_r40_c39_0 = p_39_39 << 1;
  assign t_r40_c39_1 = p_40_38 << 1;
  assign t_r40_c39_2 = p_40_39 << 2;
  assign t_r40_c39_3 = p_40_40 << 1;
  assign t_r40_c39_4 = p_41_39 << 1;
  assign t_r40_c39_5 = t_r40_c39_0 + p_39_38;
  assign t_r40_c39_6 = t_r40_c39_1 + p_39_40;
  assign t_r40_c39_7 = t_r40_c39_2 + t_r40_c39_3;
  assign t_r40_c39_8 = t_r40_c39_4 + p_41_38;
  assign t_r40_c39_9 = t_r40_c39_5 + t_r40_c39_6;
  assign t_r40_c39_10 = t_r40_c39_7 + t_r40_c39_8;
  assign t_r40_c39_11 = t_r40_c39_9 + t_r40_c39_10;
  assign t_r40_c39_12 = t_r40_c39_11 + p_41_40;
  assign out_40_39 = t_r40_c39_12 >> 4;

  assign t_r40_c40_0 = p_39_40 << 1;
  assign t_r40_c40_1 = p_40_39 << 1;
  assign t_r40_c40_2 = p_40_40 << 2;
  assign t_r40_c40_3 = p_40_41 << 1;
  assign t_r40_c40_4 = p_41_40 << 1;
  assign t_r40_c40_5 = t_r40_c40_0 + p_39_39;
  assign t_r40_c40_6 = t_r40_c40_1 + p_39_41;
  assign t_r40_c40_7 = t_r40_c40_2 + t_r40_c40_3;
  assign t_r40_c40_8 = t_r40_c40_4 + p_41_39;
  assign t_r40_c40_9 = t_r40_c40_5 + t_r40_c40_6;
  assign t_r40_c40_10 = t_r40_c40_7 + t_r40_c40_8;
  assign t_r40_c40_11 = t_r40_c40_9 + t_r40_c40_10;
  assign t_r40_c40_12 = t_r40_c40_11 + p_41_41;
  assign out_40_40 = t_r40_c40_12 >> 4;

  assign t_r40_c41_0 = p_39_41 << 1;
  assign t_r40_c41_1 = p_40_40 << 1;
  assign t_r40_c41_2 = p_40_41 << 2;
  assign t_r40_c41_3 = p_40_42 << 1;
  assign t_r40_c41_4 = p_41_41 << 1;
  assign t_r40_c41_5 = t_r40_c41_0 + p_39_40;
  assign t_r40_c41_6 = t_r40_c41_1 + p_39_42;
  assign t_r40_c41_7 = t_r40_c41_2 + t_r40_c41_3;
  assign t_r40_c41_8 = t_r40_c41_4 + p_41_40;
  assign t_r40_c41_9 = t_r40_c41_5 + t_r40_c41_6;
  assign t_r40_c41_10 = t_r40_c41_7 + t_r40_c41_8;
  assign t_r40_c41_11 = t_r40_c41_9 + t_r40_c41_10;
  assign t_r40_c41_12 = t_r40_c41_11 + p_41_42;
  assign out_40_41 = t_r40_c41_12 >> 4;

  assign t_r40_c42_0 = p_39_42 << 1;
  assign t_r40_c42_1 = p_40_41 << 1;
  assign t_r40_c42_2 = p_40_42 << 2;
  assign t_r40_c42_3 = p_40_43 << 1;
  assign t_r40_c42_4 = p_41_42 << 1;
  assign t_r40_c42_5 = t_r40_c42_0 + p_39_41;
  assign t_r40_c42_6 = t_r40_c42_1 + p_39_43;
  assign t_r40_c42_7 = t_r40_c42_2 + t_r40_c42_3;
  assign t_r40_c42_8 = t_r40_c42_4 + p_41_41;
  assign t_r40_c42_9 = t_r40_c42_5 + t_r40_c42_6;
  assign t_r40_c42_10 = t_r40_c42_7 + t_r40_c42_8;
  assign t_r40_c42_11 = t_r40_c42_9 + t_r40_c42_10;
  assign t_r40_c42_12 = t_r40_c42_11 + p_41_43;
  assign out_40_42 = t_r40_c42_12 >> 4;

  assign t_r40_c43_0 = p_39_43 << 1;
  assign t_r40_c43_1 = p_40_42 << 1;
  assign t_r40_c43_2 = p_40_43 << 2;
  assign t_r40_c43_3 = p_40_44 << 1;
  assign t_r40_c43_4 = p_41_43 << 1;
  assign t_r40_c43_5 = t_r40_c43_0 + p_39_42;
  assign t_r40_c43_6 = t_r40_c43_1 + p_39_44;
  assign t_r40_c43_7 = t_r40_c43_2 + t_r40_c43_3;
  assign t_r40_c43_8 = t_r40_c43_4 + p_41_42;
  assign t_r40_c43_9 = t_r40_c43_5 + t_r40_c43_6;
  assign t_r40_c43_10 = t_r40_c43_7 + t_r40_c43_8;
  assign t_r40_c43_11 = t_r40_c43_9 + t_r40_c43_10;
  assign t_r40_c43_12 = t_r40_c43_11 + p_41_44;
  assign out_40_43 = t_r40_c43_12 >> 4;

  assign t_r40_c44_0 = p_39_44 << 1;
  assign t_r40_c44_1 = p_40_43 << 1;
  assign t_r40_c44_2 = p_40_44 << 2;
  assign t_r40_c44_3 = p_40_45 << 1;
  assign t_r40_c44_4 = p_41_44 << 1;
  assign t_r40_c44_5 = t_r40_c44_0 + p_39_43;
  assign t_r40_c44_6 = t_r40_c44_1 + p_39_45;
  assign t_r40_c44_7 = t_r40_c44_2 + t_r40_c44_3;
  assign t_r40_c44_8 = t_r40_c44_4 + p_41_43;
  assign t_r40_c44_9 = t_r40_c44_5 + t_r40_c44_6;
  assign t_r40_c44_10 = t_r40_c44_7 + t_r40_c44_8;
  assign t_r40_c44_11 = t_r40_c44_9 + t_r40_c44_10;
  assign t_r40_c44_12 = t_r40_c44_11 + p_41_45;
  assign out_40_44 = t_r40_c44_12 >> 4;

  assign t_r40_c45_0 = p_39_45 << 1;
  assign t_r40_c45_1 = p_40_44 << 1;
  assign t_r40_c45_2 = p_40_45 << 2;
  assign t_r40_c45_3 = p_40_46 << 1;
  assign t_r40_c45_4 = p_41_45 << 1;
  assign t_r40_c45_5 = t_r40_c45_0 + p_39_44;
  assign t_r40_c45_6 = t_r40_c45_1 + p_39_46;
  assign t_r40_c45_7 = t_r40_c45_2 + t_r40_c45_3;
  assign t_r40_c45_8 = t_r40_c45_4 + p_41_44;
  assign t_r40_c45_9 = t_r40_c45_5 + t_r40_c45_6;
  assign t_r40_c45_10 = t_r40_c45_7 + t_r40_c45_8;
  assign t_r40_c45_11 = t_r40_c45_9 + t_r40_c45_10;
  assign t_r40_c45_12 = t_r40_c45_11 + p_41_46;
  assign out_40_45 = t_r40_c45_12 >> 4;

  assign t_r40_c46_0 = p_39_46 << 1;
  assign t_r40_c46_1 = p_40_45 << 1;
  assign t_r40_c46_2 = p_40_46 << 2;
  assign t_r40_c46_3 = p_40_47 << 1;
  assign t_r40_c46_4 = p_41_46 << 1;
  assign t_r40_c46_5 = t_r40_c46_0 + p_39_45;
  assign t_r40_c46_6 = t_r40_c46_1 + p_39_47;
  assign t_r40_c46_7 = t_r40_c46_2 + t_r40_c46_3;
  assign t_r40_c46_8 = t_r40_c46_4 + p_41_45;
  assign t_r40_c46_9 = t_r40_c46_5 + t_r40_c46_6;
  assign t_r40_c46_10 = t_r40_c46_7 + t_r40_c46_8;
  assign t_r40_c46_11 = t_r40_c46_9 + t_r40_c46_10;
  assign t_r40_c46_12 = t_r40_c46_11 + p_41_47;
  assign out_40_46 = t_r40_c46_12 >> 4;

  assign t_r40_c47_0 = p_39_47 << 1;
  assign t_r40_c47_1 = p_40_46 << 1;
  assign t_r40_c47_2 = p_40_47 << 2;
  assign t_r40_c47_3 = p_40_48 << 1;
  assign t_r40_c47_4 = p_41_47 << 1;
  assign t_r40_c47_5 = t_r40_c47_0 + p_39_46;
  assign t_r40_c47_6 = t_r40_c47_1 + p_39_48;
  assign t_r40_c47_7 = t_r40_c47_2 + t_r40_c47_3;
  assign t_r40_c47_8 = t_r40_c47_4 + p_41_46;
  assign t_r40_c47_9 = t_r40_c47_5 + t_r40_c47_6;
  assign t_r40_c47_10 = t_r40_c47_7 + t_r40_c47_8;
  assign t_r40_c47_11 = t_r40_c47_9 + t_r40_c47_10;
  assign t_r40_c47_12 = t_r40_c47_11 + p_41_48;
  assign out_40_47 = t_r40_c47_12 >> 4;

  assign t_r40_c48_0 = p_39_48 << 1;
  assign t_r40_c48_1 = p_40_47 << 1;
  assign t_r40_c48_2 = p_40_48 << 2;
  assign t_r40_c48_3 = p_40_49 << 1;
  assign t_r40_c48_4 = p_41_48 << 1;
  assign t_r40_c48_5 = t_r40_c48_0 + p_39_47;
  assign t_r40_c48_6 = t_r40_c48_1 + p_39_49;
  assign t_r40_c48_7 = t_r40_c48_2 + t_r40_c48_3;
  assign t_r40_c48_8 = t_r40_c48_4 + p_41_47;
  assign t_r40_c48_9 = t_r40_c48_5 + t_r40_c48_6;
  assign t_r40_c48_10 = t_r40_c48_7 + t_r40_c48_8;
  assign t_r40_c48_11 = t_r40_c48_9 + t_r40_c48_10;
  assign t_r40_c48_12 = t_r40_c48_11 + p_41_49;
  assign out_40_48 = t_r40_c48_12 >> 4;

  assign t_r40_c49_0 = p_39_49 << 1;
  assign t_r40_c49_1 = p_40_48 << 1;
  assign t_r40_c49_2 = p_40_49 << 2;
  assign t_r40_c49_3 = p_40_50 << 1;
  assign t_r40_c49_4 = p_41_49 << 1;
  assign t_r40_c49_5 = t_r40_c49_0 + p_39_48;
  assign t_r40_c49_6 = t_r40_c49_1 + p_39_50;
  assign t_r40_c49_7 = t_r40_c49_2 + t_r40_c49_3;
  assign t_r40_c49_8 = t_r40_c49_4 + p_41_48;
  assign t_r40_c49_9 = t_r40_c49_5 + t_r40_c49_6;
  assign t_r40_c49_10 = t_r40_c49_7 + t_r40_c49_8;
  assign t_r40_c49_11 = t_r40_c49_9 + t_r40_c49_10;
  assign t_r40_c49_12 = t_r40_c49_11 + p_41_50;
  assign out_40_49 = t_r40_c49_12 >> 4;

  assign t_r40_c50_0 = p_39_50 << 1;
  assign t_r40_c50_1 = p_40_49 << 1;
  assign t_r40_c50_2 = p_40_50 << 2;
  assign t_r40_c50_3 = p_40_51 << 1;
  assign t_r40_c50_4 = p_41_50 << 1;
  assign t_r40_c50_5 = t_r40_c50_0 + p_39_49;
  assign t_r40_c50_6 = t_r40_c50_1 + p_39_51;
  assign t_r40_c50_7 = t_r40_c50_2 + t_r40_c50_3;
  assign t_r40_c50_8 = t_r40_c50_4 + p_41_49;
  assign t_r40_c50_9 = t_r40_c50_5 + t_r40_c50_6;
  assign t_r40_c50_10 = t_r40_c50_7 + t_r40_c50_8;
  assign t_r40_c50_11 = t_r40_c50_9 + t_r40_c50_10;
  assign t_r40_c50_12 = t_r40_c50_11 + p_41_51;
  assign out_40_50 = t_r40_c50_12 >> 4;

  assign t_r40_c51_0 = p_39_51 << 1;
  assign t_r40_c51_1 = p_40_50 << 1;
  assign t_r40_c51_2 = p_40_51 << 2;
  assign t_r40_c51_3 = p_40_52 << 1;
  assign t_r40_c51_4 = p_41_51 << 1;
  assign t_r40_c51_5 = t_r40_c51_0 + p_39_50;
  assign t_r40_c51_6 = t_r40_c51_1 + p_39_52;
  assign t_r40_c51_7 = t_r40_c51_2 + t_r40_c51_3;
  assign t_r40_c51_8 = t_r40_c51_4 + p_41_50;
  assign t_r40_c51_9 = t_r40_c51_5 + t_r40_c51_6;
  assign t_r40_c51_10 = t_r40_c51_7 + t_r40_c51_8;
  assign t_r40_c51_11 = t_r40_c51_9 + t_r40_c51_10;
  assign t_r40_c51_12 = t_r40_c51_11 + p_41_52;
  assign out_40_51 = t_r40_c51_12 >> 4;

  assign t_r40_c52_0 = p_39_52 << 1;
  assign t_r40_c52_1 = p_40_51 << 1;
  assign t_r40_c52_2 = p_40_52 << 2;
  assign t_r40_c52_3 = p_40_53 << 1;
  assign t_r40_c52_4 = p_41_52 << 1;
  assign t_r40_c52_5 = t_r40_c52_0 + p_39_51;
  assign t_r40_c52_6 = t_r40_c52_1 + p_39_53;
  assign t_r40_c52_7 = t_r40_c52_2 + t_r40_c52_3;
  assign t_r40_c52_8 = t_r40_c52_4 + p_41_51;
  assign t_r40_c52_9 = t_r40_c52_5 + t_r40_c52_6;
  assign t_r40_c52_10 = t_r40_c52_7 + t_r40_c52_8;
  assign t_r40_c52_11 = t_r40_c52_9 + t_r40_c52_10;
  assign t_r40_c52_12 = t_r40_c52_11 + p_41_53;
  assign out_40_52 = t_r40_c52_12 >> 4;

  assign t_r40_c53_0 = p_39_53 << 1;
  assign t_r40_c53_1 = p_40_52 << 1;
  assign t_r40_c53_2 = p_40_53 << 2;
  assign t_r40_c53_3 = p_40_54 << 1;
  assign t_r40_c53_4 = p_41_53 << 1;
  assign t_r40_c53_5 = t_r40_c53_0 + p_39_52;
  assign t_r40_c53_6 = t_r40_c53_1 + p_39_54;
  assign t_r40_c53_7 = t_r40_c53_2 + t_r40_c53_3;
  assign t_r40_c53_8 = t_r40_c53_4 + p_41_52;
  assign t_r40_c53_9 = t_r40_c53_5 + t_r40_c53_6;
  assign t_r40_c53_10 = t_r40_c53_7 + t_r40_c53_8;
  assign t_r40_c53_11 = t_r40_c53_9 + t_r40_c53_10;
  assign t_r40_c53_12 = t_r40_c53_11 + p_41_54;
  assign out_40_53 = t_r40_c53_12 >> 4;

  assign t_r40_c54_0 = p_39_54 << 1;
  assign t_r40_c54_1 = p_40_53 << 1;
  assign t_r40_c54_2 = p_40_54 << 2;
  assign t_r40_c54_3 = p_40_55 << 1;
  assign t_r40_c54_4 = p_41_54 << 1;
  assign t_r40_c54_5 = t_r40_c54_0 + p_39_53;
  assign t_r40_c54_6 = t_r40_c54_1 + p_39_55;
  assign t_r40_c54_7 = t_r40_c54_2 + t_r40_c54_3;
  assign t_r40_c54_8 = t_r40_c54_4 + p_41_53;
  assign t_r40_c54_9 = t_r40_c54_5 + t_r40_c54_6;
  assign t_r40_c54_10 = t_r40_c54_7 + t_r40_c54_8;
  assign t_r40_c54_11 = t_r40_c54_9 + t_r40_c54_10;
  assign t_r40_c54_12 = t_r40_c54_11 + p_41_55;
  assign out_40_54 = t_r40_c54_12 >> 4;

  assign t_r40_c55_0 = p_39_55 << 1;
  assign t_r40_c55_1 = p_40_54 << 1;
  assign t_r40_c55_2 = p_40_55 << 2;
  assign t_r40_c55_3 = p_40_56 << 1;
  assign t_r40_c55_4 = p_41_55 << 1;
  assign t_r40_c55_5 = t_r40_c55_0 + p_39_54;
  assign t_r40_c55_6 = t_r40_c55_1 + p_39_56;
  assign t_r40_c55_7 = t_r40_c55_2 + t_r40_c55_3;
  assign t_r40_c55_8 = t_r40_c55_4 + p_41_54;
  assign t_r40_c55_9 = t_r40_c55_5 + t_r40_c55_6;
  assign t_r40_c55_10 = t_r40_c55_7 + t_r40_c55_8;
  assign t_r40_c55_11 = t_r40_c55_9 + t_r40_c55_10;
  assign t_r40_c55_12 = t_r40_c55_11 + p_41_56;
  assign out_40_55 = t_r40_c55_12 >> 4;

  assign t_r40_c56_0 = p_39_56 << 1;
  assign t_r40_c56_1 = p_40_55 << 1;
  assign t_r40_c56_2 = p_40_56 << 2;
  assign t_r40_c56_3 = p_40_57 << 1;
  assign t_r40_c56_4 = p_41_56 << 1;
  assign t_r40_c56_5 = t_r40_c56_0 + p_39_55;
  assign t_r40_c56_6 = t_r40_c56_1 + p_39_57;
  assign t_r40_c56_7 = t_r40_c56_2 + t_r40_c56_3;
  assign t_r40_c56_8 = t_r40_c56_4 + p_41_55;
  assign t_r40_c56_9 = t_r40_c56_5 + t_r40_c56_6;
  assign t_r40_c56_10 = t_r40_c56_7 + t_r40_c56_8;
  assign t_r40_c56_11 = t_r40_c56_9 + t_r40_c56_10;
  assign t_r40_c56_12 = t_r40_c56_11 + p_41_57;
  assign out_40_56 = t_r40_c56_12 >> 4;

  assign t_r40_c57_0 = p_39_57 << 1;
  assign t_r40_c57_1 = p_40_56 << 1;
  assign t_r40_c57_2 = p_40_57 << 2;
  assign t_r40_c57_3 = p_40_58 << 1;
  assign t_r40_c57_4 = p_41_57 << 1;
  assign t_r40_c57_5 = t_r40_c57_0 + p_39_56;
  assign t_r40_c57_6 = t_r40_c57_1 + p_39_58;
  assign t_r40_c57_7 = t_r40_c57_2 + t_r40_c57_3;
  assign t_r40_c57_8 = t_r40_c57_4 + p_41_56;
  assign t_r40_c57_9 = t_r40_c57_5 + t_r40_c57_6;
  assign t_r40_c57_10 = t_r40_c57_7 + t_r40_c57_8;
  assign t_r40_c57_11 = t_r40_c57_9 + t_r40_c57_10;
  assign t_r40_c57_12 = t_r40_c57_11 + p_41_58;
  assign out_40_57 = t_r40_c57_12 >> 4;

  assign t_r40_c58_0 = p_39_58 << 1;
  assign t_r40_c58_1 = p_40_57 << 1;
  assign t_r40_c58_2 = p_40_58 << 2;
  assign t_r40_c58_3 = p_40_59 << 1;
  assign t_r40_c58_4 = p_41_58 << 1;
  assign t_r40_c58_5 = t_r40_c58_0 + p_39_57;
  assign t_r40_c58_6 = t_r40_c58_1 + p_39_59;
  assign t_r40_c58_7 = t_r40_c58_2 + t_r40_c58_3;
  assign t_r40_c58_8 = t_r40_c58_4 + p_41_57;
  assign t_r40_c58_9 = t_r40_c58_5 + t_r40_c58_6;
  assign t_r40_c58_10 = t_r40_c58_7 + t_r40_c58_8;
  assign t_r40_c58_11 = t_r40_c58_9 + t_r40_c58_10;
  assign t_r40_c58_12 = t_r40_c58_11 + p_41_59;
  assign out_40_58 = t_r40_c58_12 >> 4;

  assign t_r40_c59_0 = p_39_59 << 1;
  assign t_r40_c59_1 = p_40_58 << 1;
  assign t_r40_c59_2 = p_40_59 << 2;
  assign t_r40_c59_3 = p_40_60 << 1;
  assign t_r40_c59_4 = p_41_59 << 1;
  assign t_r40_c59_5 = t_r40_c59_0 + p_39_58;
  assign t_r40_c59_6 = t_r40_c59_1 + p_39_60;
  assign t_r40_c59_7 = t_r40_c59_2 + t_r40_c59_3;
  assign t_r40_c59_8 = t_r40_c59_4 + p_41_58;
  assign t_r40_c59_9 = t_r40_c59_5 + t_r40_c59_6;
  assign t_r40_c59_10 = t_r40_c59_7 + t_r40_c59_8;
  assign t_r40_c59_11 = t_r40_c59_9 + t_r40_c59_10;
  assign t_r40_c59_12 = t_r40_c59_11 + p_41_60;
  assign out_40_59 = t_r40_c59_12 >> 4;

  assign t_r40_c60_0 = p_39_60 << 1;
  assign t_r40_c60_1 = p_40_59 << 1;
  assign t_r40_c60_2 = p_40_60 << 2;
  assign t_r40_c60_3 = p_40_61 << 1;
  assign t_r40_c60_4 = p_41_60 << 1;
  assign t_r40_c60_5 = t_r40_c60_0 + p_39_59;
  assign t_r40_c60_6 = t_r40_c60_1 + p_39_61;
  assign t_r40_c60_7 = t_r40_c60_2 + t_r40_c60_3;
  assign t_r40_c60_8 = t_r40_c60_4 + p_41_59;
  assign t_r40_c60_9 = t_r40_c60_5 + t_r40_c60_6;
  assign t_r40_c60_10 = t_r40_c60_7 + t_r40_c60_8;
  assign t_r40_c60_11 = t_r40_c60_9 + t_r40_c60_10;
  assign t_r40_c60_12 = t_r40_c60_11 + p_41_61;
  assign out_40_60 = t_r40_c60_12 >> 4;

  assign t_r40_c61_0 = p_39_61 << 1;
  assign t_r40_c61_1 = p_40_60 << 1;
  assign t_r40_c61_2 = p_40_61 << 2;
  assign t_r40_c61_3 = p_40_62 << 1;
  assign t_r40_c61_4 = p_41_61 << 1;
  assign t_r40_c61_5 = t_r40_c61_0 + p_39_60;
  assign t_r40_c61_6 = t_r40_c61_1 + p_39_62;
  assign t_r40_c61_7 = t_r40_c61_2 + t_r40_c61_3;
  assign t_r40_c61_8 = t_r40_c61_4 + p_41_60;
  assign t_r40_c61_9 = t_r40_c61_5 + t_r40_c61_6;
  assign t_r40_c61_10 = t_r40_c61_7 + t_r40_c61_8;
  assign t_r40_c61_11 = t_r40_c61_9 + t_r40_c61_10;
  assign t_r40_c61_12 = t_r40_c61_11 + p_41_62;
  assign out_40_61 = t_r40_c61_12 >> 4;

  assign t_r40_c62_0 = p_39_62 << 1;
  assign t_r40_c62_1 = p_40_61 << 1;
  assign t_r40_c62_2 = p_40_62 << 2;
  assign t_r40_c62_3 = p_40_63 << 1;
  assign t_r40_c62_4 = p_41_62 << 1;
  assign t_r40_c62_5 = t_r40_c62_0 + p_39_61;
  assign t_r40_c62_6 = t_r40_c62_1 + p_39_63;
  assign t_r40_c62_7 = t_r40_c62_2 + t_r40_c62_3;
  assign t_r40_c62_8 = t_r40_c62_4 + p_41_61;
  assign t_r40_c62_9 = t_r40_c62_5 + t_r40_c62_6;
  assign t_r40_c62_10 = t_r40_c62_7 + t_r40_c62_8;
  assign t_r40_c62_11 = t_r40_c62_9 + t_r40_c62_10;
  assign t_r40_c62_12 = t_r40_c62_11 + p_41_63;
  assign out_40_62 = t_r40_c62_12 >> 4;

  assign t_r40_c63_0 = p_39_63 << 1;
  assign t_r40_c63_1 = p_40_62 << 1;
  assign t_r40_c63_2 = p_40_63 << 2;
  assign t_r40_c63_3 = p_40_64 << 1;
  assign t_r40_c63_4 = p_41_63 << 1;
  assign t_r40_c63_5 = t_r40_c63_0 + p_39_62;
  assign t_r40_c63_6 = t_r40_c63_1 + p_39_64;
  assign t_r40_c63_7 = t_r40_c63_2 + t_r40_c63_3;
  assign t_r40_c63_8 = t_r40_c63_4 + p_41_62;
  assign t_r40_c63_9 = t_r40_c63_5 + t_r40_c63_6;
  assign t_r40_c63_10 = t_r40_c63_7 + t_r40_c63_8;
  assign t_r40_c63_11 = t_r40_c63_9 + t_r40_c63_10;
  assign t_r40_c63_12 = t_r40_c63_11 + p_41_64;
  assign out_40_63 = t_r40_c63_12 >> 4;

  assign t_r40_c64_0 = p_39_64 << 1;
  assign t_r40_c64_1 = p_40_63 << 1;
  assign t_r40_c64_2 = p_40_64 << 2;
  assign t_r40_c64_3 = p_40_65 << 1;
  assign t_r40_c64_4 = p_41_64 << 1;
  assign t_r40_c64_5 = t_r40_c64_0 + p_39_63;
  assign t_r40_c64_6 = t_r40_c64_1 + p_39_65;
  assign t_r40_c64_7 = t_r40_c64_2 + t_r40_c64_3;
  assign t_r40_c64_8 = t_r40_c64_4 + p_41_63;
  assign t_r40_c64_9 = t_r40_c64_5 + t_r40_c64_6;
  assign t_r40_c64_10 = t_r40_c64_7 + t_r40_c64_8;
  assign t_r40_c64_11 = t_r40_c64_9 + t_r40_c64_10;
  assign t_r40_c64_12 = t_r40_c64_11 + p_41_65;
  assign out_40_64 = t_r40_c64_12 >> 4;

  assign t_r41_c1_0 = p_40_1 << 1;
  assign t_r41_c1_1 = p_41_0 << 1;
  assign t_r41_c1_2 = p_41_1 << 2;
  assign t_r41_c1_3 = p_41_2 << 1;
  assign t_r41_c1_4 = p_42_1 << 1;
  assign t_r41_c1_5 = t_r41_c1_0 + p_40_0;
  assign t_r41_c1_6 = t_r41_c1_1 + p_40_2;
  assign t_r41_c1_7 = t_r41_c1_2 + t_r41_c1_3;
  assign t_r41_c1_8 = t_r41_c1_4 + p_42_0;
  assign t_r41_c1_9 = t_r41_c1_5 + t_r41_c1_6;
  assign t_r41_c1_10 = t_r41_c1_7 + t_r41_c1_8;
  assign t_r41_c1_11 = t_r41_c1_9 + t_r41_c1_10;
  assign t_r41_c1_12 = t_r41_c1_11 + p_42_2;
  assign out_41_1 = t_r41_c1_12 >> 4;

  assign t_r41_c2_0 = p_40_2 << 1;
  assign t_r41_c2_1 = p_41_1 << 1;
  assign t_r41_c2_2 = p_41_2 << 2;
  assign t_r41_c2_3 = p_41_3 << 1;
  assign t_r41_c2_4 = p_42_2 << 1;
  assign t_r41_c2_5 = t_r41_c2_0 + p_40_1;
  assign t_r41_c2_6 = t_r41_c2_1 + p_40_3;
  assign t_r41_c2_7 = t_r41_c2_2 + t_r41_c2_3;
  assign t_r41_c2_8 = t_r41_c2_4 + p_42_1;
  assign t_r41_c2_9 = t_r41_c2_5 + t_r41_c2_6;
  assign t_r41_c2_10 = t_r41_c2_7 + t_r41_c2_8;
  assign t_r41_c2_11 = t_r41_c2_9 + t_r41_c2_10;
  assign t_r41_c2_12 = t_r41_c2_11 + p_42_3;
  assign out_41_2 = t_r41_c2_12 >> 4;

  assign t_r41_c3_0 = p_40_3 << 1;
  assign t_r41_c3_1 = p_41_2 << 1;
  assign t_r41_c3_2 = p_41_3 << 2;
  assign t_r41_c3_3 = p_41_4 << 1;
  assign t_r41_c3_4 = p_42_3 << 1;
  assign t_r41_c3_5 = t_r41_c3_0 + p_40_2;
  assign t_r41_c3_6 = t_r41_c3_1 + p_40_4;
  assign t_r41_c3_7 = t_r41_c3_2 + t_r41_c3_3;
  assign t_r41_c3_8 = t_r41_c3_4 + p_42_2;
  assign t_r41_c3_9 = t_r41_c3_5 + t_r41_c3_6;
  assign t_r41_c3_10 = t_r41_c3_7 + t_r41_c3_8;
  assign t_r41_c3_11 = t_r41_c3_9 + t_r41_c3_10;
  assign t_r41_c3_12 = t_r41_c3_11 + p_42_4;
  assign out_41_3 = t_r41_c3_12 >> 4;

  assign t_r41_c4_0 = p_40_4 << 1;
  assign t_r41_c4_1 = p_41_3 << 1;
  assign t_r41_c4_2 = p_41_4 << 2;
  assign t_r41_c4_3 = p_41_5 << 1;
  assign t_r41_c4_4 = p_42_4 << 1;
  assign t_r41_c4_5 = t_r41_c4_0 + p_40_3;
  assign t_r41_c4_6 = t_r41_c4_1 + p_40_5;
  assign t_r41_c4_7 = t_r41_c4_2 + t_r41_c4_3;
  assign t_r41_c4_8 = t_r41_c4_4 + p_42_3;
  assign t_r41_c4_9 = t_r41_c4_5 + t_r41_c4_6;
  assign t_r41_c4_10 = t_r41_c4_7 + t_r41_c4_8;
  assign t_r41_c4_11 = t_r41_c4_9 + t_r41_c4_10;
  assign t_r41_c4_12 = t_r41_c4_11 + p_42_5;
  assign out_41_4 = t_r41_c4_12 >> 4;

  assign t_r41_c5_0 = p_40_5 << 1;
  assign t_r41_c5_1 = p_41_4 << 1;
  assign t_r41_c5_2 = p_41_5 << 2;
  assign t_r41_c5_3 = p_41_6 << 1;
  assign t_r41_c5_4 = p_42_5 << 1;
  assign t_r41_c5_5 = t_r41_c5_0 + p_40_4;
  assign t_r41_c5_6 = t_r41_c5_1 + p_40_6;
  assign t_r41_c5_7 = t_r41_c5_2 + t_r41_c5_3;
  assign t_r41_c5_8 = t_r41_c5_4 + p_42_4;
  assign t_r41_c5_9 = t_r41_c5_5 + t_r41_c5_6;
  assign t_r41_c5_10 = t_r41_c5_7 + t_r41_c5_8;
  assign t_r41_c5_11 = t_r41_c5_9 + t_r41_c5_10;
  assign t_r41_c5_12 = t_r41_c5_11 + p_42_6;
  assign out_41_5 = t_r41_c5_12 >> 4;

  assign t_r41_c6_0 = p_40_6 << 1;
  assign t_r41_c6_1 = p_41_5 << 1;
  assign t_r41_c6_2 = p_41_6 << 2;
  assign t_r41_c6_3 = p_41_7 << 1;
  assign t_r41_c6_4 = p_42_6 << 1;
  assign t_r41_c6_5 = t_r41_c6_0 + p_40_5;
  assign t_r41_c6_6 = t_r41_c6_1 + p_40_7;
  assign t_r41_c6_7 = t_r41_c6_2 + t_r41_c6_3;
  assign t_r41_c6_8 = t_r41_c6_4 + p_42_5;
  assign t_r41_c6_9 = t_r41_c6_5 + t_r41_c6_6;
  assign t_r41_c6_10 = t_r41_c6_7 + t_r41_c6_8;
  assign t_r41_c6_11 = t_r41_c6_9 + t_r41_c6_10;
  assign t_r41_c6_12 = t_r41_c6_11 + p_42_7;
  assign out_41_6 = t_r41_c6_12 >> 4;

  assign t_r41_c7_0 = p_40_7 << 1;
  assign t_r41_c7_1 = p_41_6 << 1;
  assign t_r41_c7_2 = p_41_7 << 2;
  assign t_r41_c7_3 = p_41_8 << 1;
  assign t_r41_c7_4 = p_42_7 << 1;
  assign t_r41_c7_5 = t_r41_c7_0 + p_40_6;
  assign t_r41_c7_6 = t_r41_c7_1 + p_40_8;
  assign t_r41_c7_7 = t_r41_c7_2 + t_r41_c7_3;
  assign t_r41_c7_8 = t_r41_c7_4 + p_42_6;
  assign t_r41_c7_9 = t_r41_c7_5 + t_r41_c7_6;
  assign t_r41_c7_10 = t_r41_c7_7 + t_r41_c7_8;
  assign t_r41_c7_11 = t_r41_c7_9 + t_r41_c7_10;
  assign t_r41_c7_12 = t_r41_c7_11 + p_42_8;
  assign out_41_7 = t_r41_c7_12 >> 4;

  assign t_r41_c8_0 = p_40_8 << 1;
  assign t_r41_c8_1 = p_41_7 << 1;
  assign t_r41_c8_2 = p_41_8 << 2;
  assign t_r41_c8_3 = p_41_9 << 1;
  assign t_r41_c8_4 = p_42_8 << 1;
  assign t_r41_c8_5 = t_r41_c8_0 + p_40_7;
  assign t_r41_c8_6 = t_r41_c8_1 + p_40_9;
  assign t_r41_c8_7 = t_r41_c8_2 + t_r41_c8_3;
  assign t_r41_c8_8 = t_r41_c8_4 + p_42_7;
  assign t_r41_c8_9 = t_r41_c8_5 + t_r41_c8_6;
  assign t_r41_c8_10 = t_r41_c8_7 + t_r41_c8_8;
  assign t_r41_c8_11 = t_r41_c8_9 + t_r41_c8_10;
  assign t_r41_c8_12 = t_r41_c8_11 + p_42_9;
  assign out_41_8 = t_r41_c8_12 >> 4;

  assign t_r41_c9_0 = p_40_9 << 1;
  assign t_r41_c9_1 = p_41_8 << 1;
  assign t_r41_c9_2 = p_41_9 << 2;
  assign t_r41_c9_3 = p_41_10 << 1;
  assign t_r41_c9_4 = p_42_9 << 1;
  assign t_r41_c9_5 = t_r41_c9_0 + p_40_8;
  assign t_r41_c9_6 = t_r41_c9_1 + p_40_10;
  assign t_r41_c9_7 = t_r41_c9_2 + t_r41_c9_3;
  assign t_r41_c9_8 = t_r41_c9_4 + p_42_8;
  assign t_r41_c9_9 = t_r41_c9_5 + t_r41_c9_6;
  assign t_r41_c9_10 = t_r41_c9_7 + t_r41_c9_8;
  assign t_r41_c9_11 = t_r41_c9_9 + t_r41_c9_10;
  assign t_r41_c9_12 = t_r41_c9_11 + p_42_10;
  assign out_41_9 = t_r41_c9_12 >> 4;

  assign t_r41_c10_0 = p_40_10 << 1;
  assign t_r41_c10_1 = p_41_9 << 1;
  assign t_r41_c10_2 = p_41_10 << 2;
  assign t_r41_c10_3 = p_41_11 << 1;
  assign t_r41_c10_4 = p_42_10 << 1;
  assign t_r41_c10_5 = t_r41_c10_0 + p_40_9;
  assign t_r41_c10_6 = t_r41_c10_1 + p_40_11;
  assign t_r41_c10_7 = t_r41_c10_2 + t_r41_c10_3;
  assign t_r41_c10_8 = t_r41_c10_4 + p_42_9;
  assign t_r41_c10_9 = t_r41_c10_5 + t_r41_c10_6;
  assign t_r41_c10_10 = t_r41_c10_7 + t_r41_c10_8;
  assign t_r41_c10_11 = t_r41_c10_9 + t_r41_c10_10;
  assign t_r41_c10_12 = t_r41_c10_11 + p_42_11;
  assign out_41_10 = t_r41_c10_12 >> 4;

  assign t_r41_c11_0 = p_40_11 << 1;
  assign t_r41_c11_1 = p_41_10 << 1;
  assign t_r41_c11_2 = p_41_11 << 2;
  assign t_r41_c11_3 = p_41_12 << 1;
  assign t_r41_c11_4 = p_42_11 << 1;
  assign t_r41_c11_5 = t_r41_c11_0 + p_40_10;
  assign t_r41_c11_6 = t_r41_c11_1 + p_40_12;
  assign t_r41_c11_7 = t_r41_c11_2 + t_r41_c11_3;
  assign t_r41_c11_8 = t_r41_c11_4 + p_42_10;
  assign t_r41_c11_9 = t_r41_c11_5 + t_r41_c11_6;
  assign t_r41_c11_10 = t_r41_c11_7 + t_r41_c11_8;
  assign t_r41_c11_11 = t_r41_c11_9 + t_r41_c11_10;
  assign t_r41_c11_12 = t_r41_c11_11 + p_42_12;
  assign out_41_11 = t_r41_c11_12 >> 4;

  assign t_r41_c12_0 = p_40_12 << 1;
  assign t_r41_c12_1 = p_41_11 << 1;
  assign t_r41_c12_2 = p_41_12 << 2;
  assign t_r41_c12_3 = p_41_13 << 1;
  assign t_r41_c12_4 = p_42_12 << 1;
  assign t_r41_c12_5 = t_r41_c12_0 + p_40_11;
  assign t_r41_c12_6 = t_r41_c12_1 + p_40_13;
  assign t_r41_c12_7 = t_r41_c12_2 + t_r41_c12_3;
  assign t_r41_c12_8 = t_r41_c12_4 + p_42_11;
  assign t_r41_c12_9 = t_r41_c12_5 + t_r41_c12_6;
  assign t_r41_c12_10 = t_r41_c12_7 + t_r41_c12_8;
  assign t_r41_c12_11 = t_r41_c12_9 + t_r41_c12_10;
  assign t_r41_c12_12 = t_r41_c12_11 + p_42_13;
  assign out_41_12 = t_r41_c12_12 >> 4;

  assign t_r41_c13_0 = p_40_13 << 1;
  assign t_r41_c13_1 = p_41_12 << 1;
  assign t_r41_c13_2 = p_41_13 << 2;
  assign t_r41_c13_3 = p_41_14 << 1;
  assign t_r41_c13_4 = p_42_13 << 1;
  assign t_r41_c13_5 = t_r41_c13_0 + p_40_12;
  assign t_r41_c13_6 = t_r41_c13_1 + p_40_14;
  assign t_r41_c13_7 = t_r41_c13_2 + t_r41_c13_3;
  assign t_r41_c13_8 = t_r41_c13_4 + p_42_12;
  assign t_r41_c13_9 = t_r41_c13_5 + t_r41_c13_6;
  assign t_r41_c13_10 = t_r41_c13_7 + t_r41_c13_8;
  assign t_r41_c13_11 = t_r41_c13_9 + t_r41_c13_10;
  assign t_r41_c13_12 = t_r41_c13_11 + p_42_14;
  assign out_41_13 = t_r41_c13_12 >> 4;

  assign t_r41_c14_0 = p_40_14 << 1;
  assign t_r41_c14_1 = p_41_13 << 1;
  assign t_r41_c14_2 = p_41_14 << 2;
  assign t_r41_c14_3 = p_41_15 << 1;
  assign t_r41_c14_4 = p_42_14 << 1;
  assign t_r41_c14_5 = t_r41_c14_0 + p_40_13;
  assign t_r41_c14_6 = t_r41_c14_1 + p_40_15;
  assign t_r41_c14_7 = t_r41_c14_2 + t_r41_c14_3;
  assign t_r41_c14_8 = t_r41_c14_4 + p_42_13;
  assign t_r41_c14_9 = t_r41_c14_5 + t_r41_c14_6;
  assign t_r41_c14_10 = t_r41_c14_7 + t_r41_c14_8;
  assign t_r41_c14_11 = t_r41_c14_9 + t_r41_c14_10;
  assign t_r41_c14_12 = t_r41_c14_11 + p_42_15;
  assign out_41_14 = t_r41_c14_12 >> 4;

  assign t_r41_c15_0 = p_40_15 << 1;
  assign t_r41_c15_1 = p_41_14 << 1;
  assign t_r41_c15_2 = p_41_15 << 2;
  assign t_r41_c15_3 = p_41_16 << 1;
  assign t_r41_c15_4 = p_42_15 << 1;
  assign t_r41_c15_5 = t_r41_c15_0 + p_40_14;
  assign t_r41_c15_6 = t_r41_c15_1 + p_40_16;
  assign t_r41_c15_7 = t_r41_c15_2 + t_r41_c15_3;
  assign t_r41_c15_8 = t_r41_c15_4 + p_42_14;
  assign t_r41_c15_9 = t_r41_c15_5 + t_r41_c15_6;
  assign t_r41_c15_10 = t_r41_c15_7 + t_r41_c15_8;
  assign t_r41_c15_11 = t_r41_c15_9 + t_r41_c15_10;
  assign t_r41_c15_12 = t_r41_c15_11 + p_42_16;
  assign out_41_15 = t_r41_c15_12 >> 4;

  assign t_r41_c16_0 = p_40_16 << 1;
  assign t_r41_c16_1 = p_41_15 << 1;
  assign t_r41_c16_2 = p_41_16 << 2;
  assign t_r41_c16_3 = p_41_17 << 1;
  assign t_r41_c16_4 = p_42_16 << 1;
  assign t_r41_c16_5 = t_r41_c16_0 + p_40_15;
  assign t_r41_c16_6 = t_r41_c16_1 + p_40_17;
  assign t_r41_c16_7 = t_r41_c16_2 + t_r41_c16_3;
  assign t_r41_c16_8 = t_r41_c16_4 + p_42_15;
  assign t_r41_c16_9 = t_r41_c16_5 + t_r41_c16_6;
  assign t_r41_c16_10 = t_r41_c16_7 + t_r41_c16_8;
  assign t_r41_c16_11 = t_r41_c16_9 + t_r41_c16_10;
  assign t_r41_c16_12 = t_r41_c16_11 + p_42_17;
  assign out_41_16 = t_r41_c16_12 >> 4;

  assign t_r41_c17_0 = p_40_17 << 1;
  assign t_r41_c17_1 = p_41_16 << 1;
  assign t_r41_c17_2 = p_41_17 << 2;
  assign t_r41_c17_3 = p_41_18 << 1;
  assign t_r41_c17_4 = p_42_17 << 1;
  assign t_r41_c17_5 = t_r41_c17_0 + p_40_16;
  assign t_r41_c17_6 = t_r41_c17_1 + p_40_18;
  assign t_r41_c17_7 = t_r41_c17_2 + t_r41_c17_3;
  assign t_r41_c17_8 = t_r41_c17_4 + p_42_16;
  assign t_r41_c17_9 = t_r41_c17_5 + t_r41_c17_6;
  assign t_r41_c17_10 = t_r41_c17_7 + t_r41_c17_8;
  assign t_r41_c17_11 = t_r41_c17_9 + t_r41_c17_10;
  assign t_r41_c17_12 = t_r41_c17_11 + p_42_18;
  assign out_41_17 = t_r41_c17_12 >> 4;

  assign t_r41_c18_0 = p_40_18 << 1;
  assign t_r41_c18_1 = p_41_17 << 1;
  assign t_r41_c18_2 = p_41_18 << 2;
  assign t_r41_c18_3 = p_41_19 << 1;
  assign t_r41_c18_4 = p_42_18 << 1;
  assign t_r41_c18_5 = t_r41_c18_0 + p_40_17;
  assign t_r41_c18_6 = t_r41_c18_1 + p_40_19;
  assign t_r41_c18_7 = t_r41_c18_2 + t_r41_c18_3;
  assign t_r41_c18_8 = t_r41_c18_4 + p_42_17;
  assign t_r41_c18_9 = t_r41_c18_5 + t_r41_c18_6;
  assign t_r41_c18_10 = t_r41_c18_7 + t_r41_c18_8;
  assign t_r41_c18_11 = t_r41_c18_9 + t_r41_c18_10;
  assign t_r41_c18_12 = t_r41_c18_11 + p_42_19;
  assign out_41_18 = t_r41_c18_12 >> 4;

  assign t_r41_c19_0 = p_40_19 << 1;
  assign t_r41_c19_1 = p_41_18 << 1;
  assign t_r41_c19_2 = p_41_19 << 2;
  assign t_r41_c19_3 = p_41_20 << 1;
  assign t_r41_c19_4 = p_42_19 << 1;
  assign t_r41_c19_5 = t_r41_c19_0 + p_40_18;
  assign t_r41_c19_6 = t_r41_c19_1 + p_40_20;
  assign t_r41_c19_7 = t_r41_c19_2 + t_r41_c19_3;
  assign t_r41_c19_8 = t_r41_c19_4 + p_42_18;
  assign t_r41_c19_9 = t_r41_c19_5 + t_r41_c19_6;
  assign t_r41_c19_10 = t_r41_c19_7 + t_r41_c19_8;
  assign t_r41_c19_11 = t_r41_c19_9 + t_r41_c19_10;
  assign t_r41_c19_12 = t_r41_c19_11 + p_42_20;
  assign out_41_19 = t_r41_c19_12 >> 4;

  assign t_r41_c20_0 = p_40_20 << 1;
  assign t_r41_c20_1 = p_41_19 << 1;
  assign t_r41_c20_2 = p_41_20 << 2;
  assign t_r41_c20_3 = p_41_21 << 1;
  assign t_r41_c20_4 = p_42_20 << 1;
  assign t_r41_c20_5 = t_r41_c20_0 + p_40_19;
  assign t_r41_c20_6 = t_r41_c20_1 + p_40_21;
  assign t_r41_c20_7 = t_r41_c20_2 + t_r41_c20_3;
  assign t_r41_c20_8 = t_r41_c20_4 + p_42_19;
  assign t_r41_c20_9 = t_r41_c20_5 + t_r41_c20_6;
  assign t_r41_c20_10 = t_r41_c20_7 + t_r41_c20_8;
  assign t_r41_c20_11 = t_r41_c20_9 + t_r41_c20_10;
  assign t_r41_c20_12 = t_r41_c20_11 + p_42_21;
  assign out_41_20 = t_r41_c20_12 >> 4;

  assign t_r41_c21_0 = p_40_21 << 1;
  assign t_r41_c21_1 = p_41_20 << 1;
  assign t_r41_c21_2 = p_41_21 << 2;
  assign t_r41_c21_3 = p_41_22 << 1;
  assign t_r41_c21_4 = p_42_21 << 1;
  assign t_r41_c21_5 = t_r41_c21_0 + p_40_20;
  assign t_r41_c21_6 = t_r41_c21_1 + p_40_22;
  assign t_r41_c21_7 = t_r41_c21_2 + t_r41_c21_3;
  assign t_r41_c21_8 = t_r41_c21_4 + p_42_20;
  assign t_r41_c21_9 = t_r41_c21_5 + t_r41_c21_6;
  assign t_r41_c21_10 = t_r41_c21_7 + t_r41_c21_8;
  assign t_r41_c21_11 = t_r41_c21_9 + t_r41_c21_10;
  assign t_r41_c21_12 = t_r41_c21_11 + p_42_22;
  assign out_41_21 = t_r41_c21_12 >> 4;

  assign t_r41_c22_0 = p_40_22 << 1;
  assign t_r41_c22_1 = p_41_21 << 1;
  assign t_r41_c22_2 = p_41_22 << 2;
  assign t_r41_c22_3 = p_41_23 << 1;
  assign t_r41_c22_4 = p_42_22 << 1;
  assign t_r41_c22_5 = t_r41_c22_0 + p_40_21;
  assign t_r41_c22_6 = t_r41_c22_1 + p_40_23;
  assign t_r41_c22_7 = t_r41_c22_2 + t_r41_c22_3;
  assign t_r41_c22_8 = t_r41_c22_4 + p_42_21;
  assign t_r41_c22_9 = t_r41_c22_5 + t_r41_c22_6;
  assign t_r41_c22_10 = t_r41_c22_7 + t_r41_c22_8;
  assign t_r41_c22_11 = t_r41_c22_9 + t_r41_c22_10;
  assign t_r41_c22_12 = t_r41_c22_11 + p_42_23;
  assign out_41_22 = t_r41_c22_12 >> 4;

  assign t_r41_c23_0 = p_40_23 << 1;
  assign t_r41_c23_1 = p_41_22 << 1;
  assign t_r41_c23_2 = p_41_23 << 2;
  assign t_r41_c23_3 = p_41_24 << 1;
  assign t_r41_c23_4 = p_42_23 << 1;
  assign t_r41_c23_5 = t_r41_c23_0 + p_40_22;
  assign t_r41_c23_6 = t_r41_c23_1 + p_40_24;
  assign t_r41_c23_7 = t_r41_c23_2 + t_r41_c23_3;
  assign t_r41_c23_8 = t_r41_c23_4 + p_42_22;
  assign t_r41_c23_9 = t_r41_c23_5 + t_r41_c23_6;
  assign t_r41_c23_10 = t_r41_c23_7 + t_r41_c23_8;
  assign t_r41_c23_11 = t_r41_c23_9 + t_r41_c23_10;
  assign t_r41_c23_12 = t_r41_c23_11 + p_42_24;
  assign out_41_23 = t_r41_c23_12 >> 4;

  assign t_r41_c24_0 = p_40_24 << 1;
  assign t_r41_c24_1 = p_41_23 << 1;
  assign t_r41_c24_2 = p_41_24 << 2;
  assign t_r41_c24_3 = p_41_25 << 1;
  assign t_r41_c24_4 = p_42_24 << 1;
  assign t_r41_c24_5 = t_r41_c24_0 + p_40_23;
  assign t_r41_c24_6 = t_r41_c24_1 + p_40_25;
  assign t_r41_c24_7 = t_r41_c24_2 + t_r41_c24_3;
  assign t_r41_c24_8 = t_r41_c24_4 + p_42_23;
  assign t_r41_c24_9 = t_r41_c24_5 + t_r41_c24_6;
  assign t_r41_c24_10 = t_r41_c24_7 + t_r41_c24_8;
  assign t_r41_c24_11 = t_r41_c24_9 + t_r41_c24_10;
  assign t_r41_c24_12 = t_r41_c24_11 + p_42_25;
  assign out_41_24 = t_r41_c24_12 >> 4;

  assign t_r41_c25_0 = p_40_25 << 1;
  assign t_r41_c25_1 = p_41_24 << 1;
  assign t_r41_c25_2 = p_41_25 << 2;
  assign t_r41_c25_3 = p_41_26 << 1;
  assign t_r41_c25_4 = p_42_25 << 1;
  assign t_r41_c25_5 = t_r41_c25_0 + p_40_24;
  assign t_r41_c25_6 = t_r41_c25_1 + p_40_26;
  assign t_r41_c25_7 = t_r41_c25_2 + t_r41_c25_3;
  assign t_r41_c25_8 = t_r41_c25_4 + p_42_24;
  assign t_r41_c25_9 = t_r41_c25_5 + t_r41_c25_6;
  assign t_r41_c25_10 = t_r41_c25_7 + t_r41_c25_8;
  assign t_r41_c25_11 = t_r41_c25_9 + t_r41_c25_10;
  assign t_r41_c25_12 = t_r41_c25_11 + p_42_26;
  assign out_41_25 = t_r41_c25_12 >> 4;

  assign t_r41_c26_0 = p_40_26 << 1;
  assign t_r41_c26_1 = p_41_25 << 1;
  assign t_r41_c26_2 = p_41_26 << 2;
  assign t_r41_c26_3 = p_41_27 << 1;
  assign t_r41_c26_4 = p_42_26 << 1;
  assign t_r41_c26_5 = t_r41_c26_0 + p_40_25;
  assign t_r41_c26_6 = t_r41_c26_1 + p_40_27;
  assign t_r41_c26_7 = t_r41_c26_2 + t_r41_c26_3;
  assign t_r41_c26_8 = t_r41_c26_4 + p_42_25;
  assign t_r41_c26_9 = t_r41_c26_5 + t_r41_c26_6;
  assign t_r41_c26_10 = t_r41_c26_7 + t_r41_c26_8;
  assign t_r41_c26_11 = t_r41_c26_9 + t_r41_c26_10;
  assign t_r41_c26_12 = t_r41_c26_11 + p_42_27;
  assign out_41_26 = t_r41_c26_12 >> 4;

  assign t_r41_c27_0 = p_40_27 << 1;
  assign t_r41_c27_1 = p_41_26 << 1;
  assign t_r41_c27_2 = p_41_27 << 2;
  assign t_r41_c27_3 = p_41_28 << 1;
  assign t_r41_c27_4 = p_42_27 << 1;
  assign t_r41_c27_5 = t_r41_c27_0 + p_40_26;
  assign t_r41_c27_6 = t_r41_c27_1 + p_40_28;
  assign t_r41_c27_7 = t_r41_c27_2 + t_r41_c27_3;
  assign t_r41_c27_8 = t_r41_c27_4 + p_42_26;
  assign t_r41_c27_9 = t_r41_c27_5 + t_r41_c27_6;
  assign t_r41_c27_10 = t_r41_c27_7 + t_r41_c27_8;
  assign t_r41_c27_11 = t_r41_c27_9 + t_r41_c27_10;
  assign t_r41_c27_12 = t_r41_c27_11 + p_42_28;
  assign out_41_27 = t_r41_c27_12 >> 4;

  assign t_r41_c28_0 = p_40_28 << 1;
  assign t_r41_c28_1 = p_41_27 << 1;
  assign t_r41_c28_2 = p_41_28 << 2;
  assign t_r41_c28_3 = p_41_29 << 1;
  assign t_r41_c28_4 = p_42_28 << 1;
  assign t_r41_c28_5 = t_r41_c28_0 + p_40_27;
  assign t_r41_c28_6 = t_r41_c28_1 + p_40_29;
  assign t_r41_c28_7 = t_r41_c28_2 + t_r41_c28_3;
  assign t_r41_c28_8 = t_r41_c28_4 + p_42_27;
  assign t_r41_c28_9 = t_r41_c28_5 + t_r41_c28_6;
  assign t_r41_c28_10 = t_r41_c28_7 + t_r41_c28_8;
  assign t_r41_c28_11 = t_r41_c28_9 + t_r41_c28_10;
  assign t_r41_c28_12 = t_r41_c28_11 + p_42_29;
  assign out_41_28 = t_r41_c28_12 >> 4;

  assign t_r41_c29_0 = p_40_29 << 1;
  assign t_r41_c29_1 = p_41_28 << 1;
  assign t_r41_c29_2 = p_41_29 << 2;
  assign t_r41_c29_3 = p_41_30 << 1;
  assign t_r41_c29_4 = p_42_29 << 1;
  assign t_r41_c29_5 = t_r41_c29_0 + p_40_28;
  assign t_r41_c29_6 = t_r41_c29_1 + p_40_30;
  assign t_r41_c29_7 = t_r41_c29_2 + t_r41_c29_3;
  assign t_r41_c29_8 = t_r41_c29_4 + p_42_28;
  assign t_r41_c29_9 = t_r41_c29_5 + t_r41_c29_6;
  assign t_r41_c29_10 = t_r41_c29_7 + t_r41_c29_8;
  assign t_r41_c29_11 = t_r41_c29_9 + t_r41_c29_10;
  assign t_r41_c29_12 = t_r41_c29_11 + p_42_30;
  assign out_41_29 = t_r41_c29_12 >> 4;

  assign t_r41_c30_0 = p_40_30 << 1;
  assign t_r41_c30_1 = p_41_29 << 1;
  assign t_r41_c30_2 = p_41_30 << 2;
  assign t_r41_c30_3 = p_41_31 << 1;
  assign t_r41_c30_4 = p_42_30 << 1;
  assign t_r41_c30_5 = t_r41_c30_0 + p_40_29;
  assign t_r41_c30_6 = t_r41_c30_1 + p_40_31;
  assign t_r41_c30_7 = t_r41_c30_2 + t_r41_c30_3;
  assign t_r41_c30_8 = t_r41_c30_4 + p_42_29;
  assign t_r41_c30_9 = t_r41_c30_5 + t_r41_c30_6;
  assign t_r41_c30_10 = t_r41_c30_7 + t_r41_c30_8;
  assign t_r41_c30_11 = t_r41_c30_9 + t_r41_c30_10;
  assign t_r41_c30_12 = t_r41_c30_11 + p_42_31;
  assign out_41_30 = t_r41_c30_12 >> 4;

  assign t_r41_c31_0 = p_40_31 << 1;
  assign t_r41_c31_1 = p_41_30 << 1;
  assign t_r41_c31_2 = p_41_31 << 2;
  assign t_r41_c31_3 = p_41_32 << 1;
  assign t_r41_c31_4 = p_42_31 << 1;
  assign t_r41_c31_5 = t_r41_c31_0 + p_40_30;
  assign t_r41_c31_6 = t_r41_c31_1 + p_40_32;
  assign t_r41_c31_7 = t_r41_c31_2 + t_r41_c31_3;
  assign t_r41_c31_8 = t_r41_c31_4 + p_42_30;
  assign t_r41_c31_9 = t_r41_c31_5 + t_r41_c31_6;
  assign t_r41_c31_10 = t_r41_c31_7 + t_r41_c31_8;
  assign t_r41_c31_11 = t_r41_c31_9 + t_r41_c31_10;
  assign t_r41_c31_12 = t_r41_c31_11 + p_42_32;
  assign out_41_31 = t_r41_c31_12 >> 4;

  assign t_r41_c32_0 = p_40_32 << 1;
  assign t_r41_c32_1 = p_41_31 << 1;
  assign t_r41_c32_2 = p_41_32 << 2;
  assign t_r41_c32_3 = p_41_33 << 1;
  assign t_r41_c32_4 = p_42_32 << 1;
  assign t_r41_c32_5 = t_r41_c32_0 + p_40_31;
  assign t_r41_c32_6 = t_r41_c32_1 + p_40_33;
  assign t_r41_c32_7 = t_r41_c32_2 + t_r41_c32_3;
  assign t_r41_c32_8 = t_r41_c32_4 + p_42_31;
  assign t_r41_c32_9 = t_r41_c32_5 + t_r41_c32_6;
  assign t_r41_c32_10 = t_r41_c32_7 + t_r41_c32_8;
  assign t_r41_c32_11 = t_r41_c32_9 + t_r41_c32_10;
  assign t_r41_c32_12 = t_r41_c32_11 + p_42_33;
  assign out_41_32 = t_r41_c32_12 >> 4;

  assign t_r41_c33_0 = p_40_33 << 1;
  assign t_r41_c33_1 = p_41_32 << 1;
  assign t_r41_c33_2 = p_41_33 << 2;
  assign t_r41_c33_3 = p_41_34 << 1;
  assign t_r41_c33_4 = p_42_33 << 1;
  assign t_r41_c33_5 = t_r41_c33_0 + p_40_32;
  assign t_r41_c33_6 = t_r41_c33_1 + p_40_34;
  assign t_r41_c33_7 = t_r41_c33_2 + t_r41_c33_3;
  assign t_r41_c33_8 = t_r41_c33_4 + p_42_32;
  assign t_r41_c33_9 = t_r41_c33_5 + t_r41_c33_6;
  assign t_r41_c33_10 = t_r41_c33_7 + t_r41_c33_8;
  assign t_r41_c33_11 = t_r41_c33_9 + t_r41_c33_10;
  assign t_r41_c33_12 = t_r41_c33_11 + p_42_34;
  assign out_41_33 = t_r41_c33_12 >> 4;

  assign t_r41_c34_0 = p_40_34 << 1;
  assign t_r41_c34_1 = p_41_33 << 1;
  assign t_r41_c34_2 = p_41_34 << 2;
  assign t_r41_c34_3 = p_41_35 << 1;
  assign t_r41_c34_4 = p_42_34 << 1;
  assign t_r41_c34_5 = t_r41_c34_0 + p_40_33;
  assign t_r41_c34_6 = t_r41_c34_1 + p_40_35;
  assign t_r41_c34_7 = t_r41_c34_2 + t_r41_c34_3;
  assign t_r41_c34_8 = t_r41_c34_4 + p_42_33;
  assign t_r41_c34_9 = t_r41_c34_5 + t_r41_c34_6;
  assign t_r41_c34_10 = t_r41_c34_7 + t_r41_c34_8;
  assign t_r41_c34_11 = t_r41_c34_9 + t_r41_c34_10;
  assign t_r41_c34_12 = t_r41_c34_11 + p_42_35;
  assign out_41_34 = t_r41_c34_12 >> 4;

  assign t_r41_c35_0 = p_40_35 << 1;
  assign t_r41_c35_1 = p_41_34 << 1;
  assign t_r41_c35_2 = p_41_35 << 2;
  assign t_r41_c35_3 = p_41_36 << 1;
  assign t_r41_c35_4 = p_42_35 << 1;
  assign t_r41_c35_5 = t_r41_c35_0 + p_40_34;
  assign t_r41_c35_6 = t_r41_c35_1 + p_40_36;
  assign t_r41_c35_7 = t_r41_c35_2 + t_r41_c35_3;
  assign t_r41_c35_8 = t_r41_c35_4 + p_42_34;
  assign t_r41_c35_9 = t_r41_c35_5 + t_r41_c35_6;
  assign t_r41_c35_10 = t_r41_c35_7 + t_r41_c35_8;
  assign t_r41_c35_11 = t_r41_c35_9 + t_r41_c35_10;
  assign t_r41_c35_12 = t_r41_c35_11 + p_42_36;
  assign out_41_35 = t_r41_c35_12 >> 4;

  assign t_r41_c36_0 = p_40_36 << 1;
  assign t_r41_c36_1 = p_41_35 << 1;
  assign t_r41_c36_2 = p_41_36 << 2;
  assign t_r41_c36_3 = p_41_37 << 1;
  assign t_r41_c36_4 = p_42_36 << 1;
  assign t_r41_c36_5 = t_r41_c36_0 + p_40_35;
  assign t_r41_c36_6 = t_r41_c36_1 + p_40_37;
  assign t_r41_c36_7 = t_r41_c36_2 + t_r41_c36_3;
  assign t_r41_c36_8 = t_r41_c36_4 + p_42_35;
  assign t_r41_c36_9 = t_r41_c36_5 + t_r41_c36_6;
  assign t_r41_c36_10 = t_r41_c36_7 + t_r41_c36_8;
  assign t_r41_c36_11 = t_r41_c36_9 + t_r41_c36_10;
  assign t_r41_c36_12 = t_r41_c36_11 + p_42_37;
  assign out_41_36 = t_r41_c36_12 >> 4;

  assign t_r41_c37_0 = p_40_37 << 1;
  assign t_r41_c37_1 = p_41_36 << 1;
  assign t_r41_c37_2 = p_41_37 << 2;
  assign t_r41_c37_3 = p_41_38 << 1;
  assign t_r41_c37_4 = p_42_37 << 1;
  assign t_r41_c37_5 = t_r41_c37_0 + p_40_36;
  assign t_r41_c37_6 = t_r41_c37_1 + p_40_38;
  assign t_r41_c37_7 = t_r41_c37_2 + t_r41_c37_3;
  assign t_r41_c37_8 = t_r41_c37_4 + p_42_36;
  assign t_r41_c37_9 = t_r41_c37_5 + t_r41_c37_6;
  assign t_r41_c37_10 = t_r41_c37_7 + t_r41_c37_8;
  assign t_r41_c37_11 = t_r41_c37_9 + t_r41_c37_10;
  assign t_r41_c37_12 = t_r41_c37_11 + p_42_38;
  assign out_41_37 = t_r41_c37_12 >> 4;

  assign t_r41_c38_0 = p_40_38 << 1;
  assign t_r41_c38_1 = p_41_37 << 1;
  assign t_r41_c38_2 = p_41_38 << 2;
  assign t_r41_c38_3 = p_41_39 << 1;
  assign t_r41_c38_4 = p_42_38 << 1;
  assign t_r41_c38_5 = t_r41_c38_0 + p_40_37;
  assign t_r41_c38_6 = t_r41_c38_1 + p_40_39;
  assign t_r41_c38_7 = t_r41_c38_2 + t_r41_c38_3;
  assign t_r41_c38_8 = t_r41_c38_4 + p_42_37;
  assign t_r41_c38_9 = t_r41_c38_5 + t_r41_c38_6;
  assign t_r41_c38_10 = t_r41_c38_7 + t_r41_c38_8;
  assign t_r41_c38_11 = t_r41_c38_9 + t_r41_c38_10;
  assign t_r41_c38_12 = t_r41_c38_11 + p_42_39;
  assign out_41_38 = t_r41_c38_12 >> 4;

  assign t_r41_c39_0 = p_40_39 << 1;
  assign t_r41_c39_1 = p_41_38 << 1;
  assign t_r41_c39_2 = p_41_39 << 2;
  assign t_r41_c39_3 = p_41_40 << 1;
  assign t_r41_c39_4 = p_42_39 << 1;
  assign t_r41_c39_5 = t_r41_c39_0 + p_40_38;
  assign t_r41_c39_6 = t_r41_c39_1 + p_40_40;
  assign t_r41_c39_7 = t_r41_c39_2 + t_r41_c39_3;
  assign t_r41_c39_8 = t_r41_c39_4 + p_42_38;
  assign t_r41_c39_9 = t_r41_c39_5 + t_r41_c39_6;
  assign t_r41_c39_10 = t_r41_c39_7 + t_r41_c39_8;
  assign t_r41_c39_11 = t_r41_c39_9 + t_r41_c39_10;
  assign t_r41_c39_12 = t_r41_c39_11 + p_42_40;
  assign out_41_39 = t_r41_c39_12 >> 4;

  assign t_r41_c40_0 = p_40_40 << 1;
  assign t_r41_c40_1 = p_41_39 << 1;
  assign t_r41_c40_2 = p_41_40 << 2;
  assign t_r41_c40_3 = p_41_41 << 1;
  assign t_r41_c40_4 = p_42_40 << 1;
  assign t_r41_c40_5 = t_r41_c40_0 + p_40_39;
  assign t_r41_c40_6 = t_r41_c40_1 + p_40_41;
  assign t_r41_c40_7 = t_r41_c40_2 + t_r41_c40_3;
  assign t_r41_c40_8 = t_r41_c40_4 + p_42_39;
  assign t_r41_c40_9 = t_r41_c40_5 + t_r41_c40_6;
  assign t_r41_c40_10 = t_r41_c40_7 + t_r41_c40_8;
  assign t_r41_c40_11 = t_r41_c40_9 + t_r41_c40_10;
  assign t_r41_c40_12 = t_r41_c40_11 + p_42_41;
  assign out_41_40 = t_r41_c40_12 >> 4;

  assign t_r41_c41_0 = p_40_41 << 1;
  assign t_r41_c41_1 = p_41_40 << 1;
  assign t_r41_c41_2 = p_41_41 << 2;
  assign t_r41_c41_3 = p_41_42 << 1;
  assign t_r41_c41_4 = p_42_41 << 1;
  assign t_r41_c41_5 = t_r41_c41_0 + p_40_40;
  assign t_r41_c41_6 = t_r41_c41_1 + p_40_42;
  assign t_r41_c41_7 = t_r41_c41_2 + t_r41_c41_3;
  assign t_r41_c41_8 = t_r41_c41_4 + p_42_40;
  assign t_r41_c41_9 = t_r41_c41_5 + t_r41_c41_6;
  assign t_r41_c41_10 = t_r41_c41_7 + t_r41_c41_8;
  assign t_r41_c41_11 = t_r41_c41_9 + t_r41_c41_10;
  assign t_r41_c41_12 = t_r41_c41_11 + p_42_42;
  assign out_41_41 = t_r41_c41_12 >> 4;

  assign t_r41_c42_0 = p_40_42 << 1;
  assign t_r41_c42_1 = p_41_41 << 1;
  assign t_r41_c42_2 = p_41_42 << 2;
  assign t_r41_c42_3 = p_41_43 << 1;
  assign t_r41_c42_4 = p_42_42 << 1;
  assign t_r41_c42_5 = t_r41_c42_0 + p_40_41;
  assign t_r41_c42_6 = t_r41_c42_1 + p_40_43;
  assign t_r41_c42_7 = t_r41_c42_2 + t_r41_c42_3;
  assign t_r41_c42_8 = t_r41_c42_4 + p_42_41;
  assign t_r41_c42_9 = t_r41_c42_5 + t_r41_c42_6;
  assign t_r41_c42_10 = t_r41_c42_7 + t_r41_c42_8;
  assign t_r41_c42_11 = t_r41_c42_9 + t_r41_c42_10;
  assign t_r41_c42_12 = t_r41_c42_11 + p_42_43;
  assign out_41_42 = t_r41_c42_12 >> 4;

  assign t_r41_c43_0 = p_40_43 << 1;
  assign t_r41_c43_1 = p_41_42 << 1;
  assign t_r41_c43_2 = p_41_43 << 2;
  assign t_r41_c43_3 = p_41_44 << 1;
  assign t_r41_c43_4 = p_42_43 << 1;
  assign t_r41_c43_5 = t_r41_c43_0 + p_40_42;
  assign t_r41_c43_6 = t_r41_c43_1 + p_40_44;
  assign t_r41_c43_7 = t_r41_c43_2 + t_r41_c43_3;
  assign t_r41_c43_8 = t_r41_c43_4 + p_42_42;
  assign t_r41_c43_9 = t_r41_c43_5 + t_r41_c43_6;
  assign t_r41_c43_10 = t_r41_c43_7 + t_r41_c43_8;
  assign t_r41_c43_11 = t_r41_c43_9 + t_r41_c43_10;
  assign t_r41_c43_12 = t_r41_c43_11 + p_42_44;
  assign out_41_43 = t_r41_c43_12 >> 4;

  assign t_r41_c44_0 = p_40_44 << 1;
  assign t_r41_c44_1 = p_41_43 << 1;
  assign t_r41_c44_2 = p_41_44 << 2;
  assign t_r41_c44_3 = p_41_45 << 1;
  assign t_r41_c44_4 = p_42_44 << 1;
  assign t_r41_c44_5 = t_r41_c44_0 + p_40_43;
  assign t_r41_c44_6 = t_r41_c44_1 + p_40_45;
  assign t_r41_c44_7 = t_r41_c44_2 + t_r41_c44_3;
  assign t_r41_c44_8 = t_r41_c44_4 + p_42_43;
  assign t_r41_c44_9 = t_r41_c44_5 + t_r41_c44_6;
  assign t_r41_c44_10 = t_r41_c44_7 + t_r41_c44_8;
  assign t_r41_c44_11 = t_r41_c44_9 + t_r41_c44_10;
  assign t_r41_c44_12 = t_r41_c44_11 + p_42_45;
  assign out_41_44 = t_r41_c44_12 >> 4;

  assign t_r41_c45_0 = p_40_45 << 1;
  assign t_r41_c45_1 = p_41_44 << 1;
  assign t_r41_c45_2 = p_41_45 << 2;
  assign t_r41_c45_3 = p_41_46 << 1;
  assign t_r41_c45_4 = p_42_45 << 1;
  assign t_r41_c45_5 = t_r41_c45_0 + p_40_44;
  assign t_r41_c45_6 = t_r41_c45_1 + p_40_46;
  assign t_r41_c45_7 = t_r41_c45_2 + t_r41_c45_3;
  assign t_r41_c45_8 = t_r41_c45_4 + p_42_44;
  assign t_r41_c45_9 = t_r41_c45_5 + t_r41_c45_6;
  assign t_r41_c45_10 = t_r41_c45_7 + t_r41_c45_8;
  assign t_r41_c45_11 = t_r41_c45_9 + t_r41_c45_10;
  assign t_r41_c45_12 = t_r41_c45_11 + p_42_46;
  assign out_41_45 = t_r41_c45_12 >> 4;

  assign t_r41_c46_0 = p_40_46 << 1;
  assign t_r41_c46_1 = p_41_45 << 1;
  assign t_r41_c46_2 = p_41_46 << 2;
  assign t_r41_c46_3 = p_41_47 << 1;
  assign t_r41_c46_4 = p_42_46 << 1;
  assign t_r41_c46_5 = t_r41_c46_0 + p_40_45;
  assign t_r41_c46_6 = t_r41_c46_1 + p_40_47;
  assign t_r41_c46_7 = t_r41_c46_2 + t_r41_c46_3;
  assign t_r41_c46_8 = t_r41_c46_4 + p_42_45;
  assign t_r41_c46_9 = t_r41_c46_5 + t_r41_c46_6;
  assign t_r41_c46_10 = t_r41_c46_7 + t_r41_c46_8;
  assign t_r41_c46_11 = t_r41_c46_9 + t_r41_c46_10;
  assign t_r41_c46_12 = t_r41_c46_11 + p_42_47;
  assign out_41_46 = t_r41_c46_12 >> 4;

  assign t_r41_c47_0 = p_40_47 << 1;
  assign t_r41_c47_1 = p_41_46 << 1;
  assign t_r41_c47_2 = p_41_47 << 2;
  assign t_r41_c47_3 = p_41_48 << 1;
  assign t_r41_c47_4 = p_42_47 << 1;
  assign t_r41_c47_5 = t_r41_c47_0 + p_40_46;
  assign t_r41_c47_6 = t_r41_c47_1 + p_40_48;
  assign t_r41_c47_7 = t_r41_c47_2 + t_r41_c47_3;
  assign t_r41_c47_8 = t_r41_c47_4 + p_42_46;
  assign t_r41_c47_9 = t_r41_c47_5 + t_r41_c47_6;
  assign t_r41_c47_10 = t_r41_c47_7 + t_r41_c47_8;
  assign t_r41_c47_11 = t_r41_c47_9 + t_r41_c47_10;
  assign t_r41_c47_12 = t_r41_c47_11 + p_42_48;
  assign out_41_47 = t_r41_c47_12 >> 4;

  assign t_r41_c48_0 = p_40_48 << 1;
  assign t_r41_c48_1 = p_41_47 << 1;
  assign t_r41_c48_2 = p_41_48 << 2;
  assign t_r41_c48_3 = p_41_49 << 1;
  assign t_r41_c48_4 = p_42_48 << 1;
  assign t_r41_c48_5 = t_r41_c48_0 + p_40_47;
  assign t_r41_c48_6 = t_r41_c48_1 + p_40_49;
  assign t_r41_c48_7 = t_r41_c48_2 + t_r41_c48_3;
  assign t_r41_c48_8 = t_r41_c48_4 + p_42_47;
  assign t_r41_c48_9 = t_r41_c48_5 + t_r41_c48_6;
  assign t_r41_c48_10 = t_r41_c48_7 + t_r41_c48_8;
  assign t_r41_c48_11 = t_r41_c48_9 + t_r41_c48_10;
  assign t_r41_c48_12 = t_r41_c48_11 + p_42_49;
  assign out_41_48 = t_r41_c48_12 >> 4;

  assign t_r41_c49_0 = p_40_49 << 1;
  assign t_r41_c49_1 = p_41_48 << 1;
  assign t_r41_c49_2 = p_41_49 << 2;
  assign t_r41_c49_3 = p_41_50 << 1;
  assign t_r41_c49_4 = p_42_49 << 1;
  assign t_r41_c49_5 = t_r41_c49_0 + p_40_48;
  assign t_r41_c49_6 = t_r41_c49_1 + p_40_50;
  assign t_r41_c49_7 = t_r41_c49_2 + t_r41_c49_3;
  assign t_r41_c49_8 = t_r41_c49_4 + p_42_48;
  assign t_r41_c49_9 = t_r41_c49_5 + t_r41_c49_6;
  assign t_r41_c49_10 = t_r41_c49_7 + t_r41_c49_8;
  assign t_r41_c49_11 = t_r41_c49_9 + t_r41_c49_10;
  assign t_r41_c49_12 = t_r41_c49_11 + p_42_50;
  assign out_41_49 = t_r41_c49_12 >> 4;

  assign t_r41_c50_0 = p_40_50 << 1;
  assign t_r41_c50_1 = p_41_49 << 1;
  assign t_r41_c50_2 = p_41_50 << 2;
  assign t_r41_c50_3 = p_41_51 << 1;
  assign t_r41_c50_4 = p_42_50 << 1;
  assign t_r41_c50_5 = t_r41_c50_0 + p_40_49;
  assign t_r41_c50_6 = t_r41_c50_1 + p_40_51;
  assign t_r41_c50_7 = t_r41_c50_2 + t_r41_c50_3;
  assign t_r41_c50_8 = t_r41_c50_4 + p_42_49;
  assign t_r41_c50_9 = t_r41_c50_5 + t_r41_c50_6;
  assign t_r41_c50_10 = t_r41_c50_7 + t_r41_c50_8;
  assign t_r41_c50_11 = t_r41_c50_9 + t_r41_c50_10;
  assign t_r41_c50_12 = t_r41_c50_11 + p_42_51;
  assign out_41_50 = t_r41_c50_12 >> 4;

  assign t_r41_c51_0 = p_40_51 << 1;
  assign t_r41_c51_1 = p_41_50 << 1;
  assign t_r41_c51_2 = p_41_51 << 2;
  assign t_r41_c51_3 = p_41_52 << 1;
  assign t_r41_c51_4 = p_42_51 << 1;
  assign t_r41_c51_5 = t_r41_c51_0 + p_40_50;
  assign t_r41_c51_6 = t_r41_c51_1 + p_40_52;
  assign t_r41_c51_7 = t_r41_c51_2 + t_r41_c51_3;
  assign t_r41_c51_8 = t_r41_c51_4 + p_42_50;
  assign t_r41_c51_9 = t_r41_c51_5 + t_r41_c51_6;
  assign t_r41_c51_10 = t_r41_c51_7 + t_r41_c51_8;
  assign t_r41_c51_11 = t_r41_c51_9 + t_r41_c51_10;
  assign t_r41_c51_12 = t_r41_c51_11 + p_42_52;
  assign out_41_51 = t_r41_c51_12 >> 4;

  assign t_r41_c52_0 = p_40_52 << 1;
  assign t_r41_c52_1 = p_41_51 << 1;
  assign t_r41_c52_2 = p_41_52 << 2;
  assign t_r41_c52_3 = p_41_53 << 1;
  assign t_r41_c52_4 = p_42_52 << 1;
  assign t_r41_c52_5 = t_r41_c52_0 + p_40_51;
  assign t_r41_c52_6 = t_r41_c52_1 + p_40_53;
  assign t_r41_c52_7 = t_r41_c52_2 + t_r41_c52_3;
  assign t_r41_c52_8 = t_r41_c52_4 + p_42_51;
  assign t_r41_c52_9 = t_r41_c52_5 + t_r41_c52_6;
  assign t_r41_c52_10 = t_r41_c52_7 + t_r41_c52_8;
  assign t_r41_c52_11 = t_r41_c52_9 + t_r41_c52_10;
  assign t_r41_c52_12 = t_r41_c52_11 + p_42_53;
  assign out_41_52 = t_r41_c52_12 >> 4;

  assign t_r41_c53_0 = p_40_53 << 1;
  assign t_r41_c53_1 = p_41_52 << 1;
  assign t_r41_c53_2 = p_41_53 << 2;
  assign t_r41_c53_3 = p_41_54 << 1;
  assign t_r41_c53_4 = p_42_53 << 1;
  assign t_r41_c53_5 = t_r41_c53_0 + p_40_52;
  assign t_r41_c53_6 = t_r41_c53_1 + p_40_54;
  assign t_r41_c53_7 = t_r41_c53_2 + t_r41_c53_3;
  assign t_r41_c53_8 = t_r41_c53_4 + p_42_52;
  assign t_r41_c53_9 = t_r41_c53_5 + t_r41_c53_6;
  assign t_r41_c53_10 = t_r41_c53_7 + t_r41_c53_8;
  assign t_r41_c53_11 = t_r41_c53_9 + t_r41_c53_10;
  assign t_r41_c53_12 = t_r41_c53_11 + p_42_54;
  assign out_41_53 = t_r41_c53_12 >> 4;

  assign t_r41_c54_0 = p_40_54 << 1;
  assign t_r41_c54_1 = p_41_53 << 1;
  assign t_r41_c54_2 = p_41_54 << 2;
  assign t_r41_c54_3 = p_41_55 << 1;
  assign t_r41_c54_4 = p_42_54 << 1;
  assign t_r41_c54_5 = t_r41_c54_0 + p_40_53;
  assign t_r41_c54_6 = t_r41_c54_1 + p_40_55;
  assign t_r41_c54_7 = t_r41_c54_2 + t_r41_c54_3;
  assign t_r41_c54_8 = t_r41_c54_4 + p_42_53;
  assign t_r41_c54_9 = t_r41_c54_5 + t_r41_c54_6;
  assign t_r41_c54_10 = t_r41_c54_7 + t_r41_c54_8;
  assign t_r41_c54_11 = t_r41_c54_9 + t_r41_c54_10;
  assign t_r41_c54_12 = t_r41_c54_11 + p_42_55;
  assign out_41_54 = t_r41_c54_12 >> 4;

  assign t_r41_c55_0 = p_40_55 << 1;
  assign t_r41_c55_1 = p_41_54 << 1;
  assign t_r41_c55_2 = p_41_55 << 2;
  assign t_r41_c55_3 = p_41_56 << 1;
  assign t_r41_c55_4 = p_42_55 << 1;
  assign t_r41_c55_5 = t_r41_c55_0 + p_40_54;
  assign t_r41_c55_6 = t_r41_c55_1 + p_40_56;
  assign t_r41_c55_7 = t_r41_c55_2 + t_r41_c55_3;
  assign t_r41_c55_8 = t_r41_c55_4 + p_42_54;
  assign t_r41_c55_9 = t_r41_c55_5 + t_r41_c55_6;
  assign t_r41_c55_10 = t_r41_c55_7 + t_r41_c55_8;
  assign t_r41_c55_11 = t_r41_c55_9 + t_r41_c55_10;
  assign t_r41_c55_12 = t_r41_c55_11 + p_42_56;
  assign out_41_55 = t_r41_c55_12 >> 4;

  assign t_r41_c56_0 = p_40_56 << 1;
  assign t_r41_c56_1 = p_41_55 << 1;
  assign t_r41_c56_2 = p_41_56 << 2;
  assign t_r41_c56_3 = p_41_57 << 1;
  assign t_r41_c56_4 = p_42_56 << 1;
  assign t_r41_c56_5 = t_r41_c56_0 + p_40_55;
  assign t_r41_c56_6 = t_r41_c56_1 + p_40_57;
  assign t_r41_c56_7 = t_r41_c56_2 + t_r41_c56_3;
  assign t_r41_c56_8 = t_r41_c56_4 + p_42_55;
  assign t_r41_c56_9 = t_r41_c56_5 + t_r41_c56_6;
  assign t_r41_c56_10 = t_r41_c56_7 + t_r41_c56_8;
  assign t_r41_c56_11 = t_r41_c56_9 + t_r41_c56_10;
  assign t_r41_c56_12 = t_r41_c56_11 + p_42_57;
  assign out_41_56 = t_r41_c56_12 >> 4;

  assign t_r41_c57_0 = p_40_57 << 1;
  assign t_r41_c57_1 = p_41_56 << 1;
  assign t_r41_c57_2 = p_41_57 << 2;
  assign t_r41_c57_3 = p_41_58 << 1;
  assign t_r41_c57_4 = p_42_57 << 1;
  assign t_r41_c57_5 = t_r41_c57_0 + p_40_56;
  assign t_r41_c57_6 = t_r41_c57_1 + p_40_58;
  assign t_r41_c57_7 = t_r41_c57_2 + t_r41_c57_3;
  assign t_r41_c57_8 = t_r41_c57_4 + p_42_56;
  assign t_r41_c57_9 = t_r41_c57_5 + t_r41_c57_6;
  assign t_r41_c57_10 = t_r41_c57_7 + t_r41_c57_8;
  assign t_r41_c57_11 = t_r41_c57_9 + t_r41_c57_10;
  assign t_r41_c57_12 = t_r41_c57_11 + p_42_58;
  assign out_41_57 = t_r41_c57_12 >> 4;

  assign t_r41_c58_0 = p_40_58 << 1;
  assign t_r41_c58_1 = p_41_57 << 1;
  assign t_r41_c58_2 = p_41_58 << 2;
  assign t_r41_c58_3 = p_41_59 << 1;
  assign t_r41_c58_4 = p_42_58 << 1;
  assign t_r41_c58_5 = t_r41_c58_0 + p_40_57;
  assign t_r41_c58_6 = t_r41_c58_1 + p_40_59;
  assign t_r41_c58_7 = t_r41_c58_2 + t_r41_c58_3;
  assign t_r41_c58_8 = t_r41_c58_4 + p_42_57;
  assign t_r41_c58_9 = t_r41_c58_5 + t_r41_c58_6;
  assign t_r41_c58_10 = t_r41_c58_7 + t_r41_c58_8;
  assign t_r41_c58_11 = t_r41_c58_9 + t_r41_c58_10;
  assign t_r41_c58_12 = t_r41_c58_11 + p_42_59;
  assign out_41_58 = t_r41_c58_12 >> 4;

  assign t_r41_c59_0 = p_40_59 << 1;
  assign t_r41_c59_1 = p_41_58 << 1;
  assign t_r41_c59_2 = p_41_59 << 2;
  assign t_r41_c59_3 = p_41_60 << 1;
  assign t_r41_c59_4 = p_42_59 << 1;
  assign t_r41_c59_5 = t_r41_c59_0 + p_40_58;
  assign t_r41_c59_6 = t_r41_c59_1 + p_40_60;
  assign t_r41_c59_7 = t_r41_c59_2 + t_r41_c59_3;
  assign t_r41_c59_8 = t_r41_c59_4 + p_42_58;
  assign t_r41_c59_9 = t_r41_c59_5 + t_r41_c59_6;
  assign t_r41_c59_10 = t_r41_c59_7 + t_r41_c59_8;
  assign t_r41_c59_11 = t_r41_c59_9 + t_r41_c59_10;
  assign t_r41_c59_12 = t_r41_c59_11 + p_42_60;
  assign out_41_59 = t_r41_c59_12 >> 4;

  assign t_r41_c60_0 = p_40_60 << 1;
  assign t_r41_c60_1 = p_41_59 << 1;
  assign t_r41_c60_2 = p_41_60 << 2;
  assign t_r41_c60_3 = p_41_61 << 1;
  assign t_r41_c60_4 = p_42_60 << 1;
  assign t_r41_c60_5 = t_r41_c60_0 + p_40_59;
  assign t_r41_c60_6 = t_r41_c60_1 + p_40_61;
  assign t_r41_c60_7 = t_r41_c60_2 + t_r41_c60_3;
  assign t_r41_c60_8 = t_r41_c60_4 + p_42_59;
  assign t_r41_c60_9 = t_r41_c60_5 + t_r41_c60_6;
  assign t_r41_c60_10 = t_r41_c60_7 + t_r41_c60_8;
  assign t_r41_c60_11 = t_r41_c60_9 + t_r41_c60_10;
  assign t_r41_c60_12 = t_r41_c60_11 + p_42_61;
  assign out_41_60 = t_r41_c60_12 >> 4;

  assign t_r41_c61_0 = p_40_61 << 1;
  assign t_r41_c61_1 = p_41_60 << 1;
  assign t_r41_c61_2 = p_41_61 << 2;
  assign t_r41_c61_3 = p_41_62 << 1;
  assign t_r41_c61_4 = p_42_61 << 1;
  assign t_r41_c61_5 = t_r41_c61_0 + p_40_60;
  assign t_r41_c61_6 = t_r41_c61_1 + p_40_62;
  assign t_r41_c61_7 = t_r41_c61_2 + t_r41_c61_3;
  assign t_r41_c61_8 = t_r41_c61_4 + p_42_60;
  assign t_r41_c61_9 = t_r41_c61_5 + t_r41_c61_6;
  assign t_r41_c61_10 = t_r41_c61_7 + t_r41_c61_8;
  assign t_r41_c61_11 = t_r41_c61_9 + t_r41_c61_10;
  assign t_r41_c61_12 = t_r41_c61_11 + p_42_62;
  assign out_41_61 = t_r41_c61_12 >> 4;

  assign t_r41_c62_0 = p_40_62 << 1;
  assign t_r41_c62_1 = p_41_61 << 1;
  assign t_r41_c62_2 = p_41_62 << 2;
  assign t_r41_c62_3 = p_41_63 << 1;
  assign t_r41_c62_4 = p_42_62 << 1;
  assign t_r41_c62_5 = t_r41_c62_0 + p_40_61;
  assign t_r41_c62_6 = t_r41_c62_1 + p_40_63;
  assign t_r41_c62_7 = t_r41_c62_2 + t_r41_c62_3;
  assign t_r41_c62_8 = t_r41_c62_4 + p_42_61;
  assign t_r41_c62_9 = t_r41_c62_5 + t_r41_c62_6;
  assign t_r41_c62_10 = t_r41_c62_7 + t_r41_c62_8;
  assign t_r41_c62_11 = t_r41_c62_9 + t_r41_c62_10;
  assign t_r41_c62_12 = t_r41_c62_11 + p_42_63;
  assign out_41_62 = t_r41_c62_12 >> 4;

  assign t_r41_c63_0 = p_40_63 << 1;
  assign t_r41_c63_1 = p_41_62 << 1;
  assign t_r41_c63_2 = p_41_63 << 2;
  assign t_r41_c63_3 = p_41_64 << 1;
  assign t_r41_c63_4 = p_42_63 << 1;
  assign t_r41_c63_5 = t_r41_c63_0 + p_40_62;
  assign t_r41_c63_6 = t_r41_c63_1 + p_40_64;
  assign t_r41_c63_7 = t_r41_c63_2 + t_r41_c63_3;
  assign t_r41_c63_8 = t_r41_c63_4 + p_42_62;
  assign t_r41_c63_9 = t_r41_c63_5 + t_r41_c63_6;
  assign t_r41_c63_10 = t_r41_c63_7 + t_r41_c63_8;
  assign t_r41_c63_11 = t_r41_c63_9 + t_r41_c63_10;
  assign t_r41_c63_12 = t_r41_c63_11 + p_42_64;
  assign out_41_63 = t_r41_c63_12 >> 4;

  assign t_r41_c64_0 = p_40_64 << 1;
  assign t_r41_c64_1 = p_41_63 << 1;
  assign t_r41_c64_2 = p_41_64 << 2;
  assign t_r41_c64_3 = p_41_65 << 1;
  assign t_r41_c64_4 = p_42_64 << 1;
  assign t_r41_c64_5 = t_r41_c64_0 + p_40_63;
  assign t_r41_c64_6 = t_r41_c64_1 + p_40_65;
  assign t_r41_c64_7 = t_r41_c64_2 + t_r41_c64_3;
  assign t_r41_c64_8 = t_r41_c64_4 + p_42_63;
  assign t_r41_c64_9 = t_r41_c64_5 + t_r41_c64_6;
  assign t_r41_c64_10 = t_r41_c64_7 + t_r41_c64_8;
  assign t_r41_c64_11 = t_r41_c64_9 + t_r41_c64_10;
  assign t_r41_c64_12 = t_r41_c64_11 + p_42_65;
  assign out_41_64 = t_r41_c64_12 >> 4;

  assign t_r42_c1_0 = p_41_1 << 1;
  assign t_r42_c1_1 = p_42_0 << 1;
  assign t_r42_c1_2 = p_42_1 << 2;
  assign t_r42_c1_3 = p_42_2 << 1;
  assign t_r42_c1_4 = p_43_1 << 1;
  assign t_r42_c1_5 = t_r42_c1_0 + p_41_0;
  assign t_r42_c1_6 = t_r42_c1_1 + p_41_2;
  assign t_r42_c1_7 = t_r42_c1_2 + t_r42_c1_3;
  assign t_r42_c1_8 = t_r42_c1_4 + p_43_0;
  assign t_r42_c1_9 = t_r42_c1_5 + t_r42_c1_6;
  assign t_r42_c1_10 = t_r42_c1_7 + t_r42_c1_8;
  assign t_r42_c1_11 = t_r42_c1_9 + t_r42_c1_10;
  assign t_r42_c1_12 = t_r42_c1_11 + p_43_2;
  assign out_42_1 = t_r42_c1_12 >> 4;

  assign t_r42_c2_0 = p_41_2 << 1;
  assign t_r42_c2_1 = p_42_1 << 1;
  assign t_r42_c2_2 = p_42_2 << 2;
  assign t_r42_c2_3 = p_42_3 << 1;
  assign t_r42_c2_4 = p_43_2 << 1;
  assign t_r42_c2_5 = t_r42_c2_0 + p_41_1;
  assign t_r42_c2_6 = t_r42_c2_1 + p_41_3;
  assign t_r42_c2_7 = t_r42_c2_2 + t_r42_c2_3;
  assign t_r42_c2_8 = t_r42_c2_4 + p_43_1;
  assign t_r42_c2_9 = t_r42_c2_5 + t_r42_c2_6;
  assign t_r42_c2_10 = t_r42_c2_7 + t_r42_c2_8;
  assign t_r42_c2_11 = t_r42_c2_9 + t_r42_c2_10;
  assign t_r42_c2_12 = t_r42_c2_11 + p_43_3;
  assign out_42_2 = t_r42_c2_12 >> 4;

  assign t_r42_c3_0 = p_41_3 << 1;
  assign t_r42_c3_1 = p_42_2 << 1;
  assign t_r42_c3_2 = p_42_3 << 2;
  assign t_r42_c3_3 = p_42_4 << 1;
  assign t_r42_c3_4 = p_43_3 << 1;
  assign t_r42_c3_5 = t_r42_c3_0 + p_41_2;
  assign t_r42_c3_6 = t_r42_c3_1 + p_41_4;
  assign t_r42_c3_7 = t_r42_c3_2 + t_r42_c3_3;
  assign t_r42_c3_8 = t_r42_c3_4 + p_43_2;
  assign t_r42_c3_9 = t_r42_c3_5 + t_r42_c3_6;
  assign t_r42_c3_10 = t_r42_c3_7 + t_r42_c3_8;
  assign t_r42_c3_11 = t_r42_c3_9 + t_r42_c3_10;
  assign t_r42_c3_12 = t_r42_c3_11 + p_43_4;
  assign out_42_3 = t_r42_c3_12 >> 4;

  assign t_r42_c4_0 = p_41_4 << 1;
  assign t_r42_c4_1 = p_42_3 << 1;
  assign t_r42_c4_2 = p_42_4 << 2;
  assign t_r42_c4_3 = p_42_5 << 1;
  assign t_r42_c4_4 = p_43_4 << 1;
  assign t_r42_c4_5 = t_r42_c4_0 + p_41_3;
  assign t_r42_c4_6 = t_r42_c4_1 + p_41_5;
  assign t_r42_c4_7 = t_r42_c4_2 + t_r42_c4_3;
  assign t_r42_c4_8 = t_r42_c4_4 + p_43_3;
  assign t_r42_c4_9 = t_r42_c4_5 + t_r42_c4_6;
  assign t_r42_c4_10 = t_r42_c4_7 + t_r42_c4_8;
  assign t_r42_c4_11 = t_r42_c4_9 + t_r42_c4_10;
  assign t_r42_c4_12 = t_r42_c4_11 + p_43_5;
  assign out_42_4 = t_r42_c4_12 >> 4;

  assign t_r42_c5_0 = p_41_5 << 1;
  assign t_r42_c5_1 = p_42_4 << 1;
  assign t_r42_c5_2 = p_42_5 << 2;
  assign t_r42_c5_3 = p_42_6 << 1;
  assign t_r42_c5_4 = p_43_5 << 1;
  assign t_r42_c5_5 = t_r42_c5_0 + p_41_4;
  assign t_r42_c5_6 = t_r42_c5_1 + p_41_6;
  assign t_r42_c5_7 = t_r42_c5_2 + t_r42_c5_3;
  assign t_r42_c5_8 = t_r42_c5_4 + p_43_4;
  assign t_r42_c5_9 = t_r42_c5_5 + t_r42_c5_6;
  assign t_r42_c5_10 = t_r42_c5_7 + t_r42_c5_8;
  assign t_r42_c5_11 = t_r42_c5_9 + t_r42_c5_10;
  assign t_r42_c5_12 = t_r42_c5_11 + p_43_6;
  assign out_42_5 = t_r42_c5_12 >> 4;

  assign t_r42_c6_0 = p_41_6 << 1;
  assign t_r42_c6_1 = p_42_5 << 1;
  assign t_r42_c6_2 = p_42_6 << 2;
  assign t_r42_c6_3 = p_42_7 << 1;
  assign t_r42_c6_4 = p_43_6 << 1;
  assign t_r42_c6_5 = t_r42_c6_0 + p_41_5;
  assign t_r42_c6_6 = t_r42_c6_1 + p_41_7;
  assign t_r42_c6_7 = t_r42_c6_2 + t_r42_c6_3;
  assign t_r42_c6_8 = t_r42_c6_4 + p_43_5;
  assign t_r42_c6_9 = t_r42_c6_5 + t_r42_c6_6;
  assign t_r42_c6_10 = t_r42_c6_7 + t_r42_c6_8;
  assign t_r42_c6_11 = t_r42_c6_9 + t_r42_c6_10;
  assign t_r42_c6_12 = t_r42_c6_11 + p_43_7;
  assign out_42_6 = t_r42_c6_12 >> 4;

  assign t_r42_c7_0 = p_41_7 << 1;
  assign t_r42_c7_1 = p_42_6 << 1;
  assign t_r42_c7_2 = p_42_7 << 2;
  assign t_r42_c7_3 = p_42_8 << 1;
  assign t_r42_c7_4 = p_43_7 << 1;
  assign t_r42_c7_5 = t_r42_c7_0 + p_41_6;
  assign t_r42_c7_6 = t_r42_c7_1 + p_41_8;
  assign t_r42_c7_7 = t_r42_c7_2 + t_r42_c7_3;
  assign t_r42_c7_8 = t_r42_c7_4 + p_43_6;
  assign t_r42_c7_9 = t_r42_c7_5 + t_r42_c7_6;
  assign t_r42_c7_10 = t_r42_c7_7 + t_r42_c7_8;
  assign t_r42_c7_11 = t_r42_c7_9 + t_r42_c7_10;
  assign t_r42_c7_12 = t_r42_c7_11 + p_43_8;
  assign out_42_7 = t_r42_c7_12 >> 4;

  assign t_r42_c8_0 = p_41_8 << 1;
  assign t_r42_c8_1 = p_42_7 << 1;
  assign t_r42_c8_2 = p_42_8 << 2;
  assign t_r42_c8_3 = p_42_9 << 1;
  assign t_r42_c8_4 = p_43_8 << 1;
  assign t_r42_c8_5 = t_r42_c8_0 + p_41_7;
  assign t_r42_c8_6 = t_r42_c8_1 + p_41_9;
  assign t_r42_c8_7 = t_r42_c8_2 + t_r42_c8_3;
  assign t_r42_c8_8 = t_r42_c8_4 + p_43_7;
  assign t_r42_c8_9 = t_r42_c8_5 + t_r42_c8_6;
  assign t_r42_c8_10 = t_r42_c8_7 + t_r42_c8_8;
  assign t_r42_c8_11 = t_r42_c8_9 + t_r42_c8_10;
  assign t_r42_c8_12 = t_r42_c8_11 + p_43_9;
  assign out_42_8 = t_r42_c8_12 >> 4;

  assign t_r42_c9_0 = p_41_9 << 1;
  assign t_r42_c9_1 = p_42_8 << 1;
  assign t_r42_c9_2 = p_42_9 << 2;
  assign t_r42_c9_3 = p_42_10 << 1;
  assign t_r42_c9_4 = p_43_9 << 1;
  assign t_r42_c9_5 = t_r42_c9_0 + p_41_8;
  assign t_r42_c9_6 = t_r42_c9_1 + p_41_10;
  assign t_r42_c9_7 = t_r42_c9_2 + t_r42_c9_3;
  assign t_r42_c9_8 = t_r42_c9_4 + p_43_8;
  assign t_r42_c9_9 = t_r42_c9_5 + t_r42_c9_6;
  assign t_r42_c9_10 = t_r42_c9_7 + t_r42_c9_8;
  assign t_r42_c9_11 = t_r42_c9_9 + t_r42_c9_10;
  assign t_r42_c9_12 = t_r42_c9_11 + p_43_10;
  assign out_42_9 = t_r42_c9_12 >> 4;

  assign t_r42_c10_0 = p_41_10 << 1;
  assign t_r42_c10_1 = p_42_9 << 1;
  assign t_r42_c10_2 = p_42_10 << 2;
  assign t_r42_c10_3 = p_42_11 << 1;
  assign t_r42_c10_4 = p_43_10 << 1;
  assign t_r42_c10_5 = t_r42_c10_0 + p_41_9;
  assign t_r42_c10_6 = t_r42_c10_1 + p_41_11;
  assign t_r42_c10_7 = t_r42_c10_2 + t_r42_c10_3;
  assign t_r42_c10_8 = t_r42_c10_4 + p_43_9;
  assign t_r42_c10_9 = t_r42_c10_5 + t_r42_c10_6;
  assign t_r42_c10_10 = t_r42_c10_7 + t_r42_c10_8;
  assign t_r42_c10_11 = t_r42_c10_9 + t_r42_c10_10;
  assign t_r42_c10_12 = t_r42_c10_11 + p_43_11;
  assign out_42_10 = t_r42_c10_12 >> 4;

  assign t_r42_c11_0 = p_41_11 << 1;
  assign t_r42_c11_1 = p_42_10 << 1;
  assign t_r42_c11_2 = p_42_11 << 2;
  assign t_r42_c11_3 = p_42_12 << 1;
  assign t_r42_c11_4 = p_43_11 << 1;
  assign t_r42_c11_5 = t_r42_c11_0 + p_41_10;
  assign t_r42_c11_6 = t_r42_c11_1 + p_41_12;
  assign t_r42_c11_7 = t_r42_c11_2 + t_r42_c11_3;
  assign t_r42_c11_8 = t_r42_c11_4 + p_43_10;
  assign t_r42_c11_9 = t_r42_c11_5 + t_r42_c11_6;
  assign t_r42_c11_10 = t_r42_c11_7 + t_r42_c11_8;
  assign t_r42_c11_11 = t_r42_c11_9 + t_r42_c11_10;
  assign t_r42_c11_12 = t_r42_c11_11 + p_43_12;
  assign out_42_11 = t_r42_c11_12 >> 4;

  assign t_r42_c12_0 = p_41_12 << 1;
  assign t_r42_c12_1 = p_42_11 << 1;
  assign t_r42_c12_2 = p_42_12 << 2;
  assign t_r42_c12_3 = p_42_13 << 1;
  assign t_r42_c12_4 = p_43_12 << 1;
  assign t_r42_c12_5 = t_r42_c12_0 + p_41_11;
  assign t_r42_c12_6 = t_r42_c12_1 + p_41_13;
  assign t_r42_c12_7 = t_r42_c12_2 + t_r42_c12_3;
  assign t_r42_c12_8 = t_r42_c12_4 + p_43_11;
  assign t_r42_c12_9 = t_r42_c12_5 + t_r42_c12_6;
  assign t_r42_c12_10 = t_r42_c12_7 + t_r42_c12_8;
  assign t_r42_c12_11 = t_r42_c12_9 + t_r42_c12_10;
  assign t_r42_c12_12 = t_r42_c12_11 + p_43_13;
  assign out_42_12 = t_r42_c12_12 >> 4;

  assign t_r42_c13_0 = p_41_13 << 1;
  assign t_r42_c13_1 = p_42_12 << 1;
  assign t_r42_c13_2 = p_42_13 << 2;
  assign t_r42_c13_3 = p_42_14 << 1;
  assign t_r42_c13_4 = p_43_13 << 1;
  assign t_r42_c13_5 = t_r42_c13_0 + p_41_12;
  assign t_r42_c13_6 = t_r42_c13_1 + p_41_14;
  assign t_r42_c13_7 = t_r42_c13_2 + t_r42_c13_3;
  assign t_r42_c13_8 = t_r42_c13_4 + p_43_12;
  assign t_r42_c13_9 = t_r42_c13_5 + t_r42_c13_6;
  assign t_r42_c13_10 = t_r42_c13_7 + t_r42_c13_8;
  assign t_r42_c13_11 = t_r42_c13_9 + t_r42_c13_10;
  assign t_r42_c13_12 = t_r42_c13_11 + p_43_14;
  assign out_42_13 = t_r42_c13_12 >> 4;

  assign t_r42_c14_0 = p_41_14 << 1;
  assign t_r42_c14_1 = p_42_13 << 1;
  assign t_r42_c14_2 = p_42_14 << 2;
  assign t_r42_c14_3 = p_42_15 << 1;
  assign t_r42_c14_4 = p_43_14 << 1;
  assign t_r42_c14_5 = t_r42_c14_0 + p_41_13;
  assign t_r42_c14_6 = t_r42_c14_1 + p_41_15;
  assign t_r42_c14_7 = t_r42_c14_2 + t_r42_c14_3;
  assign t_r42_c14_8 = t_r42_c14_4 + p_43_13;
  assign t_r42_c14_9 = t_r42_c14_5 + t_r42_c14_6;
  assign t_r42_c14_10 = t_r42_c14_7 + t_r42_c14_8;
  assign t_r42_c14_11 = t_r42_c14_9 + t_r42_c14_10;
  assign t_r42_c14_12 = t_r42_c14_11 + p_43_15;
  assign out_42_14 = t_r42_c14_12 >> 4;

  assign t_r42_c15_0 = p_41_15 << 1;
  assign t_r42_c15_1 = p_42_14 << 1;
  assign t_r42_c15_2 = p_42_15 << 2;
  assign t_r42_c15_3 = p_42_16 << 1;
  assign t_r42_c15_4 = p_43_15 << 1;
  assign t_r42_c15_5 = t_r42_c15_0 + p_41_14;
  assign t_r42_c15_6 = t_r42_c15_1 + p_41_16;
  assign t_r42_c15_7 = t_r42_c15_2 + t_r42_c15_3;
  assign t_r42_c15_8 = t_r42_c15_4 + p_43_14;
  assign t_r42_c15_9 = t_r42_c15_5 + t_r42_c15_6;
  assign t_r42_c15_10 = t_r42_c15_7 + t_r42_c15_8;
  assign t_r42_c15_11 = t_r42_c15_9 + t_r42_c15_10;
  assign t_r42_c15_12 = t_r42_c15_11 + p_43_16;
  assign out_42_15 = t_r42_c15_12 >> 4;

  assign t_r42_c16_0 = p_41_16 << 1;
  assign t_r42_c16_1 = p_42_15 << 1;
  assign t_r42_c16_2 = p_42_16 << 2;
  assign t_r42_c16_3 = p_42_17 << 1;
  assign t_r42_c16_4 = p_43_16 << 1;
  assign t_r42_c16_5 = t_r42_c16_0 + p_41_15;
  assign t_r42_c16_6 = t_r42_c16_1 + p_41_17;
  assign t_r42_c16_7 = t_r42_c16_2 + t_r42_c16_3;
  assign t_r42_c16_8 = t_r42_c16_4 + p_43_15;
  assign t_r42_c16_9 = t_r42_c16_5 + t_r42_c16_6;
  assign t_r42_c16_10 = t_r42_c16_7 + t_r42_c16_8;
  assign t_r42_c16_11 = t_r42_c16_9 + t_r42_c16_10;
  assign t_r42_c16_12 = t_r42_c16_11 + p_43_17;
  assign out_42_16 = t_r42_c16_12 >> 4;

  assign t_r42_c17_0 = p_41_17 << 1;
  assign t_r42_c17_1 = p_42_16 << 1;
  assign t_r42_c17_2 = p_42_17 << 2;
  assign t_r42_c17_3 = p_42_18 << 1;
  assign t_r42_c17_4 = p_43_17 << 1;
  assign t_r42_c17_5 = t_r42_c17_0 + p_41_16;
  assign t_r42_c17_6 = t_r42_c17_1 + p_41_18;
  assign t_r42_c17_7 = t_r42_c17_2 + t_r42_c17_3;
  assign t_r42_c17_8 = t_r42_c17_4 + p_43_16;
  assign t_r42_c17_9 = t_r42_c17_5 + t_r42_c17_6;
  assign t_r42_c17_10 = t_r42_c17_7 + t_r42_c17_8;
  assign t_r42_c17_11 = t_r42_c17_9 + t_r42_c17_10;
  assign t_r42_c17_12 = t_r42_c17_11 + p_43_18;
  assign out_42_17 = t_r42_c17_12 >> 4;

  assign t_r42_c18_0 = p_41_18 << 1;
  assign t_r42_c18_1 = p_42_17 << 1;
  assign t_r42_c18_2 = p_42_18 << 2;
  assign t_r42_c18_3 = p_42_19 << 1;
  assign t_r42_c18_4 = p_43_18 << 1;
  assign t_r42_c18_5 = t_r42_c18_0 + p_41_17;
  assign t_r42_c18_6 = t_r42_c18_1 + p_41_19;
  assign t_r42_c18_7 = t_r42_c18_2 + t_r42_c18_3;
  assign t_r42_c18_8 = t_r42_c18_4 + p_43_17;
  assign t_r42_c18_9 = t_r42_c18_5 + t_r42_c18_6;
  assign t_r42_c18_10 = t_r42_c18_7 + t_r42_c18_8;
  assign t_r42_c18_11 = t_r42_c18_9 + t_r42_c18_10;
  assign t_r42_c18_12 = t_r42_c18_11 + p_43_19;
  assign out_42_18 = t_r42_c18_12 >> 4;

  assign t_r42_c19_0 = p_41_19 << 1;
  assign t_r42_c19_1 = p_42_18 << 1;
  assign t_r42_c19_2 = p_42_19 << 2;
  assign t_r42_c19_3 = p_42_20 << 1;
  assign t_r42_c19_4 = p_43_19 << 1;
  assign t_r42_c19_5 = t_r42_c19_0 + p_41_18;
  assign t_r42_c19_6 = t_r42_c19_1 + p_41_20;
  assign t_r42_c19_7 = t_r42_c19_2 + t_r42_c19_3;
  assign t_r42_c19_8 = t_r42_c19_4 + p_43_18;
  assign t_r42_c19_9 = t_r42_c19_5 + t_r42_c19_6;
  assign t_r42_c19_10 = t_r42_c19_7 + t_r42_c19_8;
  assign t_r42_c19_11 = t_r42_c19_9 + t_r42_c19_10;
  assign t_r42_c19_12 = t_r42_c19_11 + p_43_20;
  assign out_42_19 = t_r42_c19_12 >> 4;

  assign t_r42_c20_0 = p_41_20 << 1;
  assign t_r42_c20_1 = p_42_19 << 1;
  assign t_r42_c20_2 = p_42_20 << 2;
  assign t_r42_c20_3 = p_42_21 << 1;
  assign t_r42_c20_4 = p_43_20 << 1;
  assign t_r42_c20_5 = t_r42_c20_0 + p_41_19;
  assign t_r42_c20_6 = t_r42_c20_1 + p_41_21;
  assign t_r42_c20_7 = t_r42_c20_2 + t_r42_c20_3;
  assign t_r42_c20_8 = t_r42_c20_4 + p_43_19;
  assign t_r42_c20_9 = t_r42_c20_5 + t_r42_c20_6;
  assign t_r42_c20_10 = t_r42_c20_7 + t_r42_c20_8;
  assign t_r42_c20_11 = t_r42_c20_9 + t_r42_c20_10;
  assign t_r42_c20_12 = t_r42_c20_11 + p_43_21;
  assign out_42_20 = t_r42_c20_12 >> 4;

  assign t_r42_c21_0 = p_41_21 << 1;
  assign t_r42_c21_1 = p_42_20 << 1;
  assign t_r42_c21_2 = p_42_21 << 2;
  assign t_r42_c21_3 = p_42_22 << 1;
  assign t_r42_c21_4 = p_43_21 << 1;
  assign t_r42_c21_5 = t_r42_c21_0 + p_41_20;
  assign t_r42_c21_6 = t_r42_c21_1 + p_41_22;
  assign t_r42_c21_7 = t_r42_c21_2 + t_r42_c21_3;
  assign t_r42_c21_8 = t_r42_c21_4 + p_43_20;
  assign t_r42_c21_9 = t_r42_c21_5 + t_r42_c21_6;
  assign t_r42_c21_10 = t_r42_c21_7 + t_r42_c21_8;
  assign t_r42_c21_11 = t_r42_c21_9 + t_r42_c21_10;
  assign t_r42_c21_12 = t_r42_c21_11 + p_43_22;
  assign out_42_21 = t_r42_c21_12 >> 4;

  assign t_r42_c22_0 = p_41_22 << 1;
  assign t_r42_c22_1 = p_42_21 << 1;
  assign t_r42_c22_2 = p_42_22 << 2;
  assign t_r42_c22_3 = p_42_23 << 1;
  assign t_r42_c22_4 = p_43_22 << 1;
  assign t_r42_c22_5 = t_r42_c22_0 + p_41_21;
  assign t_r42_c22_6 = t_r42_c22_1 + p_41_23;
  assign t_r42_c22_7 = t_r42_c22_2 + t_r42_c22_3;
  assign t_r42_c22_8 = t_r42_c22_4 + p_43_21;
  assign t_r42_c22_9 = t_r42_c22_5 + t_r42_c22_6;
  assign t_r42_c22_10 = t_r42_c22_7 + t_r42_c22_8;
  assign t_r42_c22_11 = t_r42_c22_9 + t_r42_c22_10;
  assign t_r42_c22_12 = t_r42_c22_11 + p_43_23;
  assign out_42_22 = t_r42_c22_12 >> 4;

  assign t_r42_c23_0 = p_41_23 << 1;
  assign t_r42_c23_1 = p_42_22 << 1;
  assign t_r42_c23_2 = p_42_23 << 2;
  assign t_r42_c23_3 = p_42_24 << 1;
  assign t_r42_c23_4 = p_43_23 << 1;
  assign t_r42_c23_5 = t_r42_c23_0 + p_41_22;
  assign t_r42_c23_6 = t_r42_c23_1 + p_41_24;
  assign t_r42_c23_7 = t_r42_c23_2 + t_r42_c23_3;
  assign t_r42_c23_8 = t_r42_c23_4 + p_43_22;
  assign t_r42_c23_9 = t_r42_c23_5 + t_r42_c23_6;
  assign t_r42_c23_10 = t_r42_c23_7 + t_r42_c23_8;
  assign t_r42_c23_11 = t_r42_c23_9 + t_r42_c23_10;
  assign t_r42_c23_12 = t_r42_c23_11 + p_43_24;
  assign out_42_23 = t_r42_c23_12 >> 4;

  assign t_r42_c24_0 = p_41_24 << 1;
  assign t_r42_c24_1 = p_42_23 << 1;
  assign t_r42_c24_2 = p_42_24 << 2;
  assign t_r42_c24_3 = p_42_25 << 1;
  assign t_r42_c24_4 = p_43_24 << 1;
  assign t_r42_c24_5 = t_r42_c24_0 + p_41_23;
  assign t_r42_c24_6 = t_r42_c24_1 + p_41_25;
  assign t_r42_c24_7 = t_r42_c24_2 + t_r42_c24_3;
  assign t_r42_c24_8 = t_r42_c24_4 + p_43_23;
  assign t_r42_c24_9 = t_r42_c24_5 + t_r42_c24_6;
  assign t_r42_c24_10 = t_r42_c24_7 + t_r42_c24_8;
  assign t_r42_c24_11 = t_r42_c24_9 + t_r42_c24_10;
  assign t_r42_c24_12 = t_r42_c24_11 + p_43_25;
  assign out_42_24 = t_r42_c24_12 >> 4;

  assign t_r42_c25_0 = p_41_25 << 1;
  assign t_r42_c25_1 = p_42_24 << 1;
  assign t_r42_c25_2 = p_42_25 << 2;
  assign t_r42_c25_3 = p_42_26 << 1;
  assign t_r42_c25_4 = p_43_25 << 1;
  assign t_r42_c25_5 = t_r42_c25_0 + p_41_24;
  assign t_r42_c25_6 = t_r42_c25_1 + p_41_26;
  assign t_r42_c25_7 = t_r42_c25_2 + t_r42_c25_3;
  assign t_r42_c25_8 = t_r42_c25_4 + p_43_24;
  assign t_r42_c25_9 = t_r42_c25_5 + t_r42_c25_6;
  assign t_r42_c25_10 = t_r42_c25_7 + t_r42_c25_8;
  assign t_r42_c25_11 = t_r42_c25_9 + t_r42_c25_10;
  assign t_r42_c25_12 = t_r42_c25_11 + p_43_26;
  assign out_42_25 = t_r42_c25_12 >> 4;

  assign t_r42_c26_0 = p_41_26 << 1;
  assign t_r42_c26_1 = p_42_25 << 1;
  assign t_r42_c26_2 = p_42_26 << 2;
  assign t_r42_c26_3 = p_42_27 << 1;
  assign t_r42_c26_4 = p_43_26 << 1;
  assign t_r42_c26_5 = t_r42_c26_0 + p_41_25;
  assign t_r42_c26_6 = t_r42_c26_1 + p_41_27;
  assign t_r42_c26_7 = t_r42_c26_2 + t_r42_c26_3;
  assign t_r42_c26_8 = t_r42_c26_4 + p_43_25;
  assign t_r42_c26_9 = t_r42_c26_5 + t_r42_c26_6;
  assign t_r42_c26_10 = t_r42_c26_7 + t_r42_c26_8;
  assign t_r42_c26_11 = t_r42_c26_9 + t_r42_c26_10;
  assign t_r42_c26_12 = t_r42_c26_11 + p_43_27;
  assign out_42_26 = t_r42_c26_12 >> 4;

  assign t_r42_c27_0 = p_41_27 << 1;
  assign t_r42_c27_1 = p_42_26 << 1;
  assign t_r42_c27_2 = p_42_27 << 2;
  assign t_r42_c27_3 = p_42_28 << 1;
  assign t_r42_c27_4 = p_43_27 << 1;
  assign t_r42_c27_5 = t_r42_c27_0 + p_41_26;
  assign t_r42_c27_6 = t_r42_c27_1 + p_41_28;
  assign t_r42_c27_7 = t_r42_c27_2 + t_r42_c27_3;
  assign t_r42_c27_8 = t_r42_c27_4 + p_43_26;
  assign t_r42_c27_9 = t_r42_c27_5 + t_r42_c27_6;
  assign t_r42_c27_10 = t_r42_c27_7 + t_r42_c27_8;
  assign t_r42_c27_11 = t_r42_c27_9 + t_r42_c27_10;
  assign t_r42_c27_12 = t_r42_c27_11 + p_43_28;
  assign out_42_27 = t_r42_c27_12 >> 4;

  assign t_r42_c28_0 = p_41_28 << 1;
  assign t_r42_c28_1 = p_42_27 << 1;
  assign t_r42_c28_2 = p_42_28 << 2;
  assign t_r42_c28_3 = p_42_29 << 1;
  assign t_r42_c28_4 = p_43_28 << 1;
  assign t_r42_c28_5 = t_r42_c28_0 + p_41_27;
  assign t_r42_c28_6 = t_r42_c28_1 + p_41_29;
  assign t_r42_c28_7 = t_r42_c28_2 + t_r42_c28_3;
  assign t_r42_c28_8 = t_r42_c28_4 + p_43_27;
  assign t_r42_c28_9 = t_r42_c28_5 + t_r42_c28_6;
  assign t_r42_c28_10 = t_r42_c28_7 + t_r42_c28_8;
  assign t_r42_c28_11 = t_r42_c28_9 + t_r42_c28_10;
  assign t_r42_c28_12 = t_r42_c28_11 + p_43_29;
  assign out_42_28 = t_r42_c28_12 >> 4;

  assign t_r42_c29_0 = p_41_29 << 1;
  assign t_r42_c29_1 = p_42_28 << 1;
  assign t_r42_c29_2 = p_42_29 << 2;
  assign t_r42_c29_3 = p_42_30 << 1;
  assign t_r42_c29_4 = p_43_29 << 1;
  assign t_r42_c29_5 = t_r42_c29_0 + p_41_28;
  assign t_r42_c29_6 = t_r42_c29_1 + p_41_30;
  assign t_r42_c29_7 = t_r42_c29_2 + t_r42_c29_3;
  assign t_r42_c29_8 = t_r42_c29_4 + p_43_28;
  assign t_r42_c29_9 = t_r42_c29_5 + t_r42_c29_6;
  assign t_r42_c29_10 = t_r42_c29_7 + t_r42_c29_8;
  assign t_r42_c29_11 = t_r42_c29_9 + t_r42_c29_10;
  assign t_r42_c29_12 = t_r42_c29_11 + p_43_30;
  assign out_42_29 = t_r42_c29_12 >> 4;

  assign t_r42_c30_0 = p_41_30 << 1;
  assign t_r42_c30_1 = p_42_29 << 1;
  assign t_r42_c30_2 = p_42_30 << 2;
  assign t_r42_c30_3 = p_42_31 << 1;
  assign t_r42_c30_4 = p_43_30 << 1;
  assign t_r42_c30_5 = t_r42_c30_0 + p_41_29;
  assign t_r42_c30_6 = t_r42_c30_1 + p_41_31;
  assign t_r42_c30_7 = t_r42_c30_2 + t_r42_c30_3;
  assign t_r42_c30_8 = t_r42_c30_4 + p_43_29;
  assign t_r42_c30_9 = t_r42_c30_5 + t_r42_c30_6;
  assign t_r42_c30_10 = t_r42_c30_7 + t_r42_c30_8;
  assign t_r42_c30_11 = t_r42_c30_9 + t_r42_c30_10;
  assign t_r42_c30_12 = t_r42_c30_11 + p_43_31;
  assign out_42_30 = t_r42_c30_12 >> 4;

  assign t_r42_c31_0 = p_41_31 << 1;
  assign t_r42_c31_1 = p_42_30 << 1;
  assign t_r42_c31_2 = p_42_31 << 2;
  assign t_r42_c31_3 = p_42_32 << 1;
  assign t_r42_c31_4 = p_43_31 << 1;
  assign t_r42_c31_5 = t_r42_c31_0 + p_41_30;
  assign t_r42_c31_6 = t_r42_c31_1 + p_41_32;
  assign t_r42_c31_7 = t_r42_c31_2 + t_r42_c31_3;
  assign t_r42_c31_8 = t_r42_c31_4 + p_43_30;
  assign t_r42_c31_9 = t_r42_c31_5 + t_r42_c31_6;
  assign t_r42_c31_10 = t_r42_c31_7 + t_r42_c31_8;
  assign t_r42_c31_11 = t_r42_c31_9 + t_r42_c31_10;
  assign t_r42_c31_12 = t_r42_c31_11 + p_43_32;
  assign out_42_31 = t_r42_c31_12 >> 4;

  assign t_r42_c32_0 = p_41_32 << 1;
  assign t_r42_c32_1 = p_42_31 << 1;
  assign t_r42_c32_2 = p_42_32 << 2;
  assign t_r42_c32_3 = p_42_33 << 1;
  assign t_r42_c32_4 = p_43_32 << 1;
  assign t_r42_c32_5 = t_r42_c32_0 + p_41_31;
  assign t_r42_c32_6 = t_r42_c32_1 + p_41_33;
  assign t_r42_c32_7 = t_r42_c32_2 + t_r42_c32_3;
  assign t_r42_c32_8 = t_r42_c32_4 + p_43_31;
  assign t_r42_c32_9 = t_r42_c32_5 + t_r42_c32_6;
  assign t_r42_c32_10 = t_r42_c32_7 + t_r42_c32_8;
  assign t_r42_c32_11 = t_r42_c32_9 + t_r42_c32_10;
  assign t_r42_c32_12 = t_r42_c32_11 + p_43_33;
  assign out_42_32 = t_r42_c32_12 >> 4;

  assign t_r42_c33_0 = p_41_33 << 1;
  assign t_r42_c33_1 = p_42_32 << 1;
  assign t_r42_c33_2 = p_42_33 << 2;
  assign t_r42_c33_3 = p_42_34 << 1;
  assign t_r42_c33_4 = p_43_33 << 1;
  assign t_r42_c33_5 = t_r42_c33_0 + p_41_32;
  assign t_r42_c33_6 = t_r42_c33_1 + p_41_34;
  assign t_r42_c33_7 = t_r42_c33_2 + t_r42_c33_3;
  assign t_r42_c33_8 = t_r42_c33_4 + p_43_32;
  assign t_r42_c33_9 = t_r42_c33_5 + t_r42_c33_6;
  assign t_r42_c33_10 = t_r42_c33_7 + t_r42_c33_8;
  assign t_r42_c33_11 = t_r42_c33_9 + t_r42_c33_10;
  assign t_r42_c33_12 = t_r42_c33_11 + p_43_34;
  assign out_42_33 = t_r42_c33_12 >> 4;

  assign t_r42_c34_0 = p_41_34 << 1;
  assign t_r42_c34_1 = p_42_33 << 1;
  assign t_r42_c34_2 = p_42_34 << 2;
  assign t_r42_c34_3 = p_42_35 << 1;
  assign t_r42_c34_4 = p_43_34 << 1;
  assign t_r42_c34_5 = t_r42_c34_0 + p_41_33;
  assign t_r42_c34_6 = t_r42_c34_1 + p_41_35;
  assign t_r42_c34_7 = t_r42_c34_2 + t_r42_c34_3;
  assign t_r42_c34_8 = t_r42_c34_4 + p_43_33;
  assign t_r42_c34_9 = t_r42_c34_5 + t_r42_c34_6;
  assign t_r42_c34_10 = t_r42_c34_7 + t_r42_c34_8;
  assign t_r42_c34_11 = t_r42_c34_9 + t_r42_c34_10;
  assign t_r42_c34_12 = t_r42_c34_11 + p_43_35;
  assign out_42_34 = t_r42_c34_12 >> 4;

  assign t_r42_c35_0 = p_41_35 << 1;
  assign t_r42_c35_1 = p_42_34 << 1;
  assign t_r42_c35_2 = p_42_35 << 2;
  assign t_r42_c35_3 = p_42_36 << 1;
  assign t_r42_c35_4 = p_43_35 << 1;
  assign t_r42_c35_5 = t_r42_c35_0 + p_41_34;
  assign t_r42_c35_6 = t_r42_c35_1 + p_41_36;
  assign t_r42_c35_7 = t_r42_c35_2 + t_r42_c35_3;
  assign t_r42_c35_8 = t_r42_c35_4 + p_43_34;
  assign t_r42_c35_9 = t_r42_c35_5 + t_r42_c35_6;
  assign t_r42_c35_10 = t_r42_c35_7 + t_r42_c35_8;
  assign t_r42_c35_11 = t_r42_c35_9 + t_r42_c35_10;
  assign t_r42_c35_12 = t_r42_c35_11 + p_43_36;
  assign out_42_35 = t_r42_c35_12 >> 4;

  assign t_r42_c36_0 = p_41_36 << 1;
  assign t_r42_c36_1 = p_42_35 << 1;
  assign t_r42_c36_2 = p_42_36 << 2;
  assign t_r42_c36_3 = p_42_37 << 1;
  assign t_r42_c36_4 = p_43_36 << 1;
  assign t_r42_c36_5 = t_r42_c36_0 + p_41_35;
  assign t_r42_c36_6 = t_r42_c36_1 + p_41_37;
  assign t_r42_c36_7 = t_r42_c36_2 + t_r42_c36_3;
  assign t_r42_c36_8 = t_r42_c36_4 + p_43_35;
  assign t_r42_c36_9 = t_r42_c36_5 + t_r42_c36_6;
  assign t_r42_c36_10 = t_r42_c36_7 + t_r42_c36_8;
  assign t_r42_c36_11 = t_r42_c36_9 + t_r42_c36_10;
  assign t_r42_c36_12 = t_r42_c36_11 + p_43_37;
  assign out_42_36 = t_r42_c36_12 >> 4;

  assign t_r42_c37_0 = p_41_37 << 1;
  assign t_r42_c37_1 = p_42_36 << 1;
  assign t_r42_c37_2 = p_42_37 << 2;
  assign t_r42_c37_3 = p_42_38 << 1;
  assign t_r42_c37_4 = p_43_37 << 1;
  assign t_r42_c37_5 = t_r42_c37_0 + p_41_36;
  assign t_r42_c37_6 = t_r42_c37_1 + p_41_38;
  assign t_r42_c37_7 = t_r42_c37_2 + t_r42_c37_3;
  assign t_r42_c37_8 = t_r42_c37_4 + p_43_36;
  assign t_r42_c37_9 = t_r42_c37_5 + t_r42_c37_6;
  assign t_r42_c37_10 = t_r42_c37_7 + t_r42_c37_8;
  assign t_r42_c37_11 = t_r42_c37_9 + t_r42_c37_10;
  assign t_r42_c37_12 = t_r42_c37_11 + p_43_38;
  assign out_42_37 = t_r42_c37_12 >> 4;

  assign t_r42_c38_0 = p_41_38 << 1;
  assign t_r42_c38_1 = p_42_37 << 1;
  assign t_r42_c38_2 = p_42_38 << 2;
  assign t_r42_c38_3 = p_42_39 << 1;
  assign t_r42_c38_4 = p_43_38 << 1;
  assign t_r42_c38_5 = t_r42_c38_0 + p_41_37;
  assign t_r42_c38_6 = t_r42_c38_1 + p_41_39;
  assign t_r42_c38_7 = t_r42_c38_2 + t_r42_c38_3;
  assign t_r42_c38_8 = t_r42_c38_4 + p_43_37;
  assign t_r42_c38_9 = t_r42_c38_5 + t_r42_c38_6;
  assign t_r42_c38_10 = t_r42_c38_7 + t_r42_c38_8;
  assign t_r42_c38_11 = t_r42_c38_9 + t_r42_c38_10;
  assign t_r42_c38_12 = t_r42_c38_11 + p_43_39;
  assign out_42_38 = t_r42_c38_12 >> 4;

  assign t_r42_c39_0 = p_41_39 << 1;
  assign t_r42_c39_1 = p_42_38 << 1;
  assign t_r42_c39_2 = p_42_39 << 2;
  assign t_r42_c39_3 = p_42_40 << 1;
  assign t_r42_c39_4 = p_43_39 << 1;
  assign t_r42_c39_5 = t_r42_c39_0 + p_41_38;
  assign t_r42_c39_6 = t_r42_c39_1 + p_41_40;
  assign t_r42_c39_7 = t_r42_c39_2 + t_r42_c39_3;
  assign t_r42_c39_8 = t_r42_c39_4 + p_43_38;
  assign t_r42_c39_9 = t_r42_c39_5 + t_r42_c39_6;
  assign t_r42_c39_10 = t_r42_c39_7 + t_r42_c39_8;
  assign t_r42_c39_11 = t_r42_c39_9 + t_r42_c39_10;
  assign t_r42_c39_12 = t_r42_c39_11 + p_43_40;
  assign out_42_39 = t_r42_c39_12 >> 4;

  assign t_r42_c40_0 = p_41_40 << 1;
  assign t_r42_c40_1 = p_42_39 << 1;
  assign t_r42_c40_2 = p_42_40 << 2;
  assign t_r42_c40_3 = p_42_41 << 1;
  assign t_r42_c40_4 = p_43_40 << 1;
  assign t_r42_c40_5 = t_r42_c40_0 + p_41_39;
  assign t_r42_c40_6 = t_r42_c40_1 + p_41_41;
  assign t_r42_c40_7 = t_r42_c40_2 + t_r42_c40_3;
  assign t_r42_c40_8 = t_r42_c40_4 + p_43_39;
  assign t_r42_c40_9 = t_r42_c40_5 + t_r42_c40_6;
  assign t_r42_c40_10 = t_r42_c40_7 + t_r42_c40_8;
  assign t_r42_c40_11 = t_r42_c40_9 + t_r42_c40_10;
  assign t_r42_c40_12 = t_r42_c40_11 + p_43_41;
  assign out_42_40 = t_r42_c40_12 >> 4;

  assign t_r42_c41_0 = p_41_41 << 1;
  assign t_r42_c41_1 = p_42_40 << 1;
  assign t_r42_c41_2 = p_42_41 << 2;
  assign t_r42_c41_3 = p_42_42 << 1;
  assign t_r42_c41_4 = p_43_41 << 1;
  assign t_r42_c41_5 = t_r42_c41_0 + p_41_40;
  assign t_r42_c41_6 = t_r42_c41_1 + p_41_42;
  assign t_r42_c41_7 = t_r42_c41_2 + t_r42_c41_3;
  assign t_r42_c41_8 = t_r42_c41_4 + p_43_40;
  assign t_r42_c41_9 = t_r42_c41_5 + t_r42_c41_6;
  assign t_r42_c41_10 = t_r42_c41_7 + t_r42_c41_8;
  assign t_r42_c41_11 = t_r42_c41_9 + t_r42_c41_10;
  assign t_r42_c41_12 = t_r42_c41_11 + p_43_42;
  assign out_42_41 = t_r42_c41_12 >> 4;

  assign t_r42_c42_0 = p_41_42 << 1;
  assign t_r42_c42_1 = p_42_41 << 1;
  assign t_r42_c42_2 = p_42_42 << 2;
  assign t_r42_c42_3 = p_42_43 << 1;
  assign t_r42_c42_4 = p_43_42 << 1;
  assign t_r42_c42_5 = t_r42_c42_0 + p_41_41;
  assign t_r42_c42_6 = t_r42_c42_1 + p_41_43;
  assign t_r42_c42_7 = t_r42_c42_2 + t_r42_c42_3;
  assign t_r42_c42_8 = t_r42_c42_4 + p_43_41;
  assign t_r42_c42_9 = t_r42_c42_5 + t_r42_c42_6;
  assign t_r42_c42_10 = t_r42_c42_7 + t_r42_c42_8;
  assign t_r42_c42_11 = t_r42_c42_9 + t_r42_c42_10;
  assign t_r42_c42_12 = t_r42_c42_11 + p_43_43;
  assign out_42_42 = t_r42_c42_12 >> 4;

  assign t_r42_c43_0 = p_41_43 << 1;
  assign t_r42_c43_1 = p_42_42 << 1;
  assign t_r42_c43_2 = p_42_43 << 2;
  assign t_r42_c43_3 = p_42_44 << 1;
  assign t_r42_c43_4 = p_43_43 << 1;
  assign t_r42_c43_5 = t_r42_c43_0 + p_41_42;
  assign t_r42_c43_6 = t_r42_c43_1 + p_41_44;
  assign t_r42_c43_7 = t_r42_c43_2 + t_r42_c43_3;
  assign t_r42_c43_8 = t_r42_c43_4 + p_43_42;
  assign t_r42_c43_9 = t_r42_c43_5 + t_r42_c43_6;
  assign t_r42_c43_10 = t_r42_c43_7 + t_r42_c43_8;
  assign t_r42_c43_11 = t_r42_c43_9 + t_r42_c43_10;
  assign t_r42_c43_12 = t_r42_c43_11 + p_43_44;
  assign out_42_43 = t_r42_c43_12 >> 4;

  assign t_r42_c44_0 = p_41_44 << 1;
  assign t_r42_c44_1 = p_42_43 << 1;
  assign t_r42_c44_2 = p_42_44 << 2;
  assign t_r42_c44_3 = p_42_45 << 1;
  assign t_r42_c44_4 = p_43_44 << 1;
  assign t_r42_c44_5 = t_r42_c44_0 + p_41_43;
  assign t_r42_c44_6 = t_r42_c44_1 + p_41_45;
  assign t_r42_c44_7 = t_r42_c44_2 + t_r42_c44_3;
  assign t_r42_c44_8 = t_r42_c44_4 + p_43_43;
  assign t_r42_c44_9 = t_r42_c44_5 + t_r42_c44_6;
  assign t_r42_c44_10 = t_r42_c44_7 + t_r42_c44_8;
  assign t_r42_c44_11 = t_r42_c44_9 + t_r42_c44_10;
  assign t_r42_c44_12 = t_r42_c44_11 + p_43_45;
  assign out_42_44 = t_r42_c44_12 >> 4;

  assign t_r42_c45_0 = p_41_45 << 1;
  assign t_r42_c45_1 = p_42_44 << 1;
  assign t_r42_c45_2 = p_42_45 << 2;
  assign t_r42_c45_3 = p_42_46 << 1;
  assign t_r42_c45_4 = p_43_45 << 1;
  assign t_r42_c45_5 = t_r42_c45_0 + p_41_44;
  assign t_r42_c45_6 = t_r42_c45_1 + p_41_46;
  assign t_r42_c45_7 = t_r42_c45_2 + t_r42_c45_3;
  assign t_r42_c45_8 = t_r42_c45_4 + p_43_44;
  assign t_r42_c45_9 = t_r42_c45_5 + t_r42_c45_6;
  assign t_r42_c45_10 = t_r42_c45_7 + t_r42_c45_8;
  assign t_r42_c45_11 = t_r42_c45_9 + t_r42_c45_10;
  assign t_r42_c45_12 = t_r42_c45_11 + p_43_46;
  assign out_42_45 = t_r42_c45_12 >> 4;

  assign t_r42_c46_0 = p_41_46 << 1;
  assign t_r42_c46_1 = p_42_45 << 1;
  assign t_r42_c46_2 = p_42_46 << 2;
  assign t_r42_c46_3 = p_42_47 << 1;
  assign t_r42_c46_4 = p_43_46 << 1;
  assign t_r42_c46_5 = t_r42_c46_0 + p_41_45;
  assign t_r42_c46_6 = t_r42_c46_1 + p_41_47;
  assign t_r42_c46_7 = t_r42_c46_2 + t_r42_c46_3;
  assign t_r42_c46_8 = t_r42_c46_4 + p_43_45;
  assign t_r42_c46_9 = t_r42_c46_5 + t_r42_c46_6;
  assign t_r42_c46_10 = t_r42_c46_7 + t_r42_c46_8;
  assign t_r42_c46_11 = t_r42_c46_9 + t_r42_c46_10;
  assign t_r42_c46_12 = t_r42_c46_11 + p_43_47;
  assign out_42_46 = t_r42_c46_12 >> 4;

  assign t_r42_c47_0 = p_41_47 << 1;
  assign t_r42_c47_1 = p_42_46 << 1;
  assign t_r42_c47_2 = p_42_47 << 2;
  assign t_r42_c47_3 = p_42_48 << 1;
  assign t_r42_c47_4 = p_43_47 << 1;
  assign t_r42_c47_5 = t_r42_c47_0 + p_41_46;
  assign t_r42_c47_6 = t_r42_c47_1 + p_41_48;
  assign t_r42_c47_7 = t_r42_c47_2 + t_r42_c47_3;
  assign t_r42_c47_8 = t_r42_c47_4 + p_43_46;
  assign t_r42_c47_9 = t_r42_c47_5 + t_r42_c47_6;
  assign t_r42_c47_10 = t_r42_c47_7 + t_r42_c47_8;
  assign t_r42_c47_11 = t_r42_c47_9 + t_r42_c47_10;
  assign t_r42_c47_12 = t_r42_c47_11 + p_43_48;
  assign out_42_47 = t_r42_c47_12 >> 4;

  assign t_r42_c48_0 = p_41_48 << 1;
  assign t_r42_c48_1 = p_42_47 << 1;
  assign t_r42_c48_2 = p_42_48 << 2;
  assign t_r42_c48_3 = p_42_49 << 1;
  assign t_r42_c48_4 = p_43_48 << 1;
  assign t_r42_c48_5 = t_r42_c48_0 + p_41_47;
  assign t_r42_c48_6 = t_r42_c48_1 + p_41_49;
  assign t_r42_c48_7 = t_r42_c48_2 + t_r42_c48_3;
  assign t_r42_c48_8 = t_r42_c48_4 + p_43_47;
  assign t_r42_c48_9 = t_r42_c48_5 + t_r42_c48_6;
  assign t_r42_c48_10 = t_r42_c48_7 + t_r42_c48_8;
  assign t_r42_c48_11 = t_r42_c48_9 + t_r42_c48_10;
  assign t_r42_c48_12 = t_r42_c48_11 + p_43_49;
  assign out_42_48 = t_r42_c48_12 >> 4;

  assign t_r42_c49_0 = p_41_49 << 1;
  assign t_r42_c49_1 = p_42_48 << 1;
  assign t_r42_c49_2 = p_42_49 << 2;
  assign t_r42_c49_3 = p_42_50 << 1;
  assign t_r42_c49_4 = p_43_49 << 1;
  assign t_r42_c49_5 = t_r42_c49_0 + p_41_48;
  assign t_r42_c49_6 = t_r42_c49_1 + p_41_50;
  assign t_r42_c49_7 = t_r42_c49_2 + t_r42_c49_3;
  assign t_r42_c49_8 = t_r42_c49_4 + p_43_48;
  assign t_r42_c49_9 = t_r42_c49_5 + t_r42_c49_6;
  assign t_r42_c49_10 = t_r42_c49_7 + t_r42_c49_8;
  assign t_r42_c49_11 = t_r42_c49_9 + t_r42_c49_10;
  assign t_r42_c49_12 = t_r42_c49_11 + p_43_50;
  assign out_42_49 = t_r42_c49_12 >> 4;

  assign t_r42_c50_0 = p_41_50 << 1;
  assign t_r42_c50_1 = p_42_49 << 1;
  assign t_r42_c50_2 = p_42_50 << 2;
  assign t_r42_c50_3 = p_42_51 << 1;
  assign t_r42_c50_4 = p_43_50 << 1;
  assign t_r42_c50_5 = t_r42_c50_0 + p_41_49;
  assign t_r42_c50_6 = t_r42_c50_1 + p_41_51;
  assign t_r42_c50_7 = t_r42_c50_2 + t_r42_c50_3;
  assign t_r42_c50_8 = t_r42_c50_4 + p_43_49;
  assign t_r42_c50_9 = t_r42_c50_5 + t_r42_c50_6;
  assign t_r42_c50_10 = t_r42_c50_7 + t_r42_c50_8;
  assign t_r42_c50_11 = t_r42_c50_9 + t_r42_c50_10;
  assign t_r42_c50_12 = t_r42_c50_11 + p_43_51;
  assign out_42_50 = t_r42_c50_12 >> 4;

  assign t_r42_c51_0 = p_41_51 << 1;
  assign t_r42_c51_1 = p_42_50 << 1;
  assign t_r42_c51_2 = p_42_51 << 2;
  assign t_r42_c51_3 = p_42_52 << 1;
  assign t_r42_c51_4 = p_43_51 << 1;
  assign t_r42_c51_5 = t_r42_c51_0 + p_41_50;
  assign t_r42_c51_6 = t_r42_c51_1 + p_41_52;
  assign t_r42_c51_7 = t_r42_c51_2 + t_r42_c51_3;
  assign t_r42_c51_8 = t_r42_c51_4 + p_43_50;
  assign t_r42_c51_9 = t_r42_c51_5 + t_r42_c51_6;
  assign t_r42_c51_10 = t_r42_c51_7 + t_r42_c51_8;
  assign t_r42_c51_11 = t_r42_c51_9 + t_r42_c51_10;
  assign t_r42_c51_12 = t_r42_c51_11 + p_43_52;
  assign out_42_51 = t_r42_c51_12 >> 4;

  assign t_r42_c52_0 = p_41_52 << 1;
  assign t_r42_c52_1 = p_42_51 << 1;
  assign t_r42_c52_2 = p_42_52 << 2;
  assign t_r42_c52_3 = p_42_53 << 1;
  assign t_r42_c52_4 = p_43_52 << 1;
  assign t_r42_c52_5 = t_r42_c52_0 + p_41_51;
  assign t_r42_c52_6 = t_r42_c52_1 + p_41_53;
  assign t_r42_c52_7 = t_r42_c52_2 + t_r42_c52_3;
  assign t_r42_c52_8 = t_r42_c52_4 + p_43_51;
  assign t_r42_c52_9 = t_r42_c52_5 + t_r42_c52_6;
  assign t_r42_c52_10 = t_r42_c52_7 + t_r42_c52_8;
  assign t_r42_c52_11 = t_r42_c52_9 + t_r42_c52_10;
  assign t_r42_c52_12 = t_r42_c52_11 + p_43_53;
  assign out_42_52 = t_r42_c52_12 >> 4;

  assign t_r42_c53_0 = p_41_53 << 1;
  assign t_r42_c53_1 = p_42_52 << 1;
  assign t_r42_c53_2 = p_42_53 << 2;
  assign t_r42_c53_3 = p_42_54 << 1;
  assign t_r42_c53_4 = p_43_53 << 1;
  assign t_r42_c53_5 = t_r42_c53_0 + p_41_52;
  assign t_r42_c53_6 = t_r42_c53_1 + p_41_54;
  assign t_r42_c53_7 = t_r42_c53_2 + t_r42_c53_3;
  assign t_r42_c53_8 = t_r42_c53_4 + p_43_52;
  assign t_r42_c53_9 = t_r42_c53_5 + t_r42_c53_6;
  assign t_r42_c53_10 = t_r42_c53_7 + t_r42_c53_8;
  assign t_r42_c53_11 = t_r42_c53_9 + t_r42_c53_10;
  assign t_r42_c53_12 = t_r42_c53_11 + p_43_54;
  assign out_42_53 = t_r42_c53_12 >> 4;

  assign t_r42_c54_0 = p_41_54 << 1;
  assign t_r42_c54_1 = p_42_53 << 1;
  assign t_r42_c54_2 = p_42_54 << 2;
  assign t_r42_c54_3 = p_42_55 << 1;
  assign t_r42_c54_4 = p_43_54 << 1;
  assign t_r42_c54_5 = t_r42_c54_0 + p_41_53;
  assign t_r42_c54_6 = t_r42_c54_1 + p_41_55;
  assign t_r42_c54_7 = t_r42_c54_2 + t_r42_c54_3;
  assign t_r42_c54_8 = t_r42_c54_4 + p_43_53;
  assign t_r42_c54_9 = t_r42_c54_5 + t_r42_c54_6;
  assign t_r42_c54_10 = t_r42_c54_7 + t_r42_c54_8;
  assign t_r42_c54_11 = t_r42_c54_9 + t_r42_c54_10;
  assign t_r42_c54_12 = t_r42_c54_11 + p_43_55;
  assign out_42_54 = t_r42_c54_12 >> 4;

  assign t_r42_c55_0 = p_41_55 << 1;
  assign t_r42_c55_1 = p_42_54 << 1;
  assign t_r42_c55_2 = p_42_55 << 2;
  assign t_r42_c55_3 = p_42_56 << 1;
  assign t_r42_c55_4 = p_43_55 << 1;
  assign t_r42_c55_5 = t_r42_c55_0 + p_41_54;
  assign t_r42_c55_6 = t_r42_c55_1 + p_41_56;
  assign t_r42_c55_7 = t_r42_c55_2 + t_r42_c55_3;
  assign t_r42_c55_8 = t_r42_c55_4 + p_43_54;
  assign t_r42_c55_9 = t_r42_c55_5 + t_r42_c55_6;
  assign t_r42_c55_10 = t_r42_c55_7 + t_r42_c55_8;
  assign t_r42_c55_11 = t_r42_c55_9 + t_r42_c55_10;
  assign t_r42_c55_12 = t_r42_c55_11 + p_43_56;
  assign out_42_55 = t_r42_c55_12 >> 4;

  assign t_r42_c56_0 = p_41_56 << 1;
  assign t_r42_c56_1 = p_42_55 << 1;
  assign t_r42_c56_2 = p_42_56 << 2;
  assign t_r42_c56_3 = p_42_57 << 1;
  assign t_r42_c56_4 = p_43_56 << 1;
  assign t_r42_c56_5 = t_r42_c56_0 + p_41_55;
  assign t_r42_c56_6 = t_r42_c56_1 + p_41_57;
  assign t_r42_c56_7 = t_r42_c56_2 + t_r42_c56_3;
  assign t_r42_c56_8 = t_r42_c56_4 + p_43_55;
  assign t_r42_c56_9 = t_r42_c56_5 + t_r42_c56_6;
  assign t_r42_c56_10 = t_r42_c56_7 + t_r42_c56_8;
  assign t_r42_c56_11 = t_r42_c56_9 + t_r42_c56_10;
  assign t_r42_c56_12 = t_r42_c56_11 + p_43_57;
  assign out_42_56 = t_r42_c56_12 >> 4;

  assign t_r42_c57_0 = p_41_57 << 1;
  assign t_r42_c57_1 = p_42_56 << 1;
  assign t_r42_c57_2 = p_42_57 << 2;
  assign t_r42_c57_3 = p_42_58 << 1;
  assign t_r42_c57_4 = p_43_57 << 1;
  assign t_r42_c57_5 = t_r42_c57_0 + p_41_56;
  assign t_r42_c57_6 = t_r42_c57_1 + p_41_58;
  assign t_r42_c57_7 = t_r42_c57_2 + t_r42_c57_3;
  assign t_r42_c57_8 = t_r42_c57_4 + p_43_56;
  assign t_r42_c57_9 = t_r42_c57_5 + t_r42_c57_6;
  assign t_r42_c57_10 = t_r42_c57_7 + t_r42_c57_8;
  assign t_r42_c57_11 = t_r42_c57_9 + t_r42_c57_10;
  assign t_r42_c57_12 = t_r42_c57_11 + p_43_58;
  assign out_42_57 = t_r42_c57_12 >> 4;

  assign t_r42_c58_0 = p_41_58 << 1;
  assign t_r42_c58_1 = p_42_57 << 1;
  assign t_r42_c58_2 = p_42_58 << 2;
  assign t_r42_c58_3 = p_42_59 << 1;
  assign t_r42_c58_4 = p_43_58 << 1;
  assign t_r42_c58_5 = t_r42_c58_0 + p_41_57;
  assign t_r42_c58_6 = t_r42_c58_1 + p_41_59;
  assign t_r42_c58_7 = t_r42_c58_2 + t_r42_c58_3;
  assign t_r42_c58_8 = t_r42_c58_4 + p_43_57;
  assign t_r42_c58_9 = t_r42_c58_5 + t_r42_c58_6;
  assign t_r42_c58_10 = t_r42_c58_7 + t_r42_c58_8;
  assign t_r42_c58_11 = t_r42_c58_9 + t_r42_c58_10;
  assign t_r42_c58_12 = t_r42_c58_11 + p_43_59;
  assign out_42_58 = t_r42_c58_12 >> 4;

  assign t_r42_c59_0 = p_41_59 << 1;
  assign t_r42_c59_1 = p_42_58 << 1;
  assign t_r42_c59_2 = p_42_59 << 2;
  assign t_r42_c59_3 = p_42_60 << 1;
  assign t_r42_c59_4 = p_43_59 << 1;
  assign t_r42_c59_5 = t_r42_c59_0 + p_41_58;
  assign t_r42_c59_6 = t_r42_c59_1 + p_41_60;
  assign t_r42_c59_7 = t_r42_c59_2 + t_r42_c59_3;
  assign t_r42_c59_8 = t_r42_c59_4 + p_43_58;
  assign t_r42_c59_9 = t_r42_c59_5 + t_r42_c59_6;
  assign t_r42_c59_10 = t_r42_c59_7 + t_r42_c59_8;
  assign t_r42_c59_11 = t_r42_c59_9 + t_r42_c59_10;
  assign t_r42_c59_12 = t_r42_c59_11 + p_43_60;
  assign out_42_59 = t_r42_c59_12 >> 4;

  assign t_r42_c60_0 = p_41_60 << 1;
  assign t_r42_c60_1 = p_42_59 << 1;
  assign t_r42_c60_2 = p_42_60 << 2;
  assign t_r42_c60_3 = p_42_61 << 1;
  assign t_r42_c60_4 = p_43_60 << 1;
  assign t_r42_c60_5 = t_r42_c60_0 + p_41_59;
  assign t_r42_c60_6 = t_r42_c60_1 + p_41_61;
  assign t_r42_c60_7 = t_r42_c60_2 + t_r42_c60_3;
  assign t_r42_c60_8 = t_r42_c60_4 + p_43_59;
  assign t_r42_c60_9 = t_r42_c60_5 + t_r42_c60_6;
  assign t_r42_c60_10 = t_r42_c60_7 + t_r42_c60_8;
  assign t_r42_c60_11 = t_r42_c60_9 + t_r42_c60_10;
  assign t_r42_c60_12 = t_r42_c60_11 + p_43_61;
  assign out_42_60 = t_r42_c60_12 >> 4;

  assign t_r42_c61_0 = p_41_61 << 1;
  assign t_r42_c61_1 = p_42_60 << 1;
  assign t_r42_c61_2 = p_42_61 << 2;
  assign t_r42_c61_3 = p_42_62 << 1;
  assign t_r42_c61_4 = p_43_61 << 1;
  assign t_r42_c61_5 = t_r42_c61_0 + p_41_60;
  assign t_r42_c61_6 = t_r42_c61_1 + p_41_62;
  assign t_r42_c61_7 = t_r42_c61_2 + t_r42_c61_3;
  assign t_r42_c61_8 = t_r42_c61_4 + p_43_60;
  assign t_r42_c61_9 = t_r42_c61_5 + t_r42_c61_6;
  assign t_r42_c61_10 = t_r42_c61_7 + t_r42_c61_8;
  assign t_r42_c61_11 = t_r42_c61_9 + t_r42_c61_10;
  assign t_r42_c61_12 = t_r42_c61_11 + p_43_62;
  assign out_42_61 = t_r42_c61_12 >> 4;

  assign t_r42_c62_0 = p_41_62 << 1;
  assign t_r42_c62_1 = p_42_61 << 1;
  assign t_r42_c62_2 = p_42_62 << 2;
  assign t_r42_c62_3 = p_42_63 << 1;
  assign t_r42_c62_4 = p_43_62 << 1;
  assign t_r42_c62_5 = t_r42_c62_0 + p_41_61;
  assign t_r42_c62_6 = t_r42_c62_1 + p_41_63;
  assign t_r42_c62_7 = t_r42_c62_2 + t_r42_c62_3;
  assign t_r42_c62_8 = t_r42_c62_4 + p_43_61;
  assign t_r42_c62_9 = t_r42_c62_5 + t_r42_c62_6;
  assign t_r42_c62_10 = t_r42_c62_7 + t_r42_c62_8;
  assign t_r42_c62_11 = t_r42_c62_9 + t_r42_c62_10;
  assign t_r42_c62_12 = t_r42_c62_11 + p_43_63;
  assign out_42_62 = t_r42_c62_12 >> 4;

  assign t_r42_c63_0 = p_41_63 << 1;
  assign t_r42_c63_1 = p_42_62 << 1;
  assign t_r42_c63_2 = p_42_63 << 2;
  assign t_r42_c63_3 = p_42_64 << 1;
  assign t_r42_c63_4 = p_43_63 << 1;
  assign t_r42_c63_5 = t_r42_c63_0 + p_41_62;
  assign t_r42_c63_6 = t_r42_c63_1 + p_41_64;
  assign t_r42_c63_7 = t_r42_c63_2 + t_r42_c63_3;
  assign t_r42_c63_8 = t_r42_c63_4 + p_43_62;
  assign t_r42_c63_9 = t_r42_c63_5 + t_r42_c63_6;
  assign t_r42_c63_10 = t_r42_c63_7 + t_r42_c63_8;
  assign t_r42_c63_11 = t_r42_c63_9 + t_r42_c63_10;
  assign t_r42_c63_12 = t_r42_c63_11 + p_43_64;
  assign out_42_63 = t_r42_c63_12 >> 4;

  assign t_r42_c64_0 = p_41_64 << 1;
  assign t_r42_c64_1 = p_42_63 << 1;
  assign t_r42_c64_2 = p_42_64 << 2;
  assign t_r42_c64_3 = p_42_65 << 1;
  assign t_r42_c64_4 = p_43_64 << 1;
  assign t_r42_c64_5 = t_r42_c64_0 + p_41_63;
  assign t_r42_c64_6 = t_r42_c64_1 + p_41_65;
  assign t_r42_c64_7 = t_r42_c64_2 + t_r42_c64_3;
  assign t_r42_c64_8 = t_r42_c64_4 + p_43_63;
  assign t_r42_c64_9 = t_r42_c64_5 + t_r42_c64_6;
  assign t_r42_c64_10 = t_r42_c64_7 + t_r42_c64_8;
  assign t_r42_c64_11 = t_r42_c64_9 + t_r42_c64_10;
  assign t_r42_c64_12 = t_r42_c64_11 + p_43_65;
  assign out_42_64 = t_r42_c64_12 >> 4;

  assign t_r43_c1_0 = p_42_1 << 1;
  assign t_r43_c1_1 = p_43_0 << 1;
  assign t_r43_c1_2 = p_43_1 << 2;
  assign t_r43_c1_3 = p_43_2 << 1;
  assign t_r43_c1_4 = p_44_1 << 1;
  assign t_r43_c1_5 = t_r43_c1_0 + p_42_0;
  assign t_r43_c1_6 = t_r43_c1_1 + p_42_2;
  assign t_r43_c1_7 = t_r43_c1_2 + t_r43_c1_3;
  assign t_r43_c1_8 = t_r43_c1_4 + p_44_0;
  assign t_r43_c1_9 = t_r43_c1_5 + t_r43_c1_6;
  assign t_r43_c1_10 = t_r43_c1_7 + t_r43_c1_8;
  assign t_r43_c1_11 = t_r43_c1_9 + t_r43_c1_10;
  assign t_r43_c1_12 = t_r43_c1_11 + p_44_2;
  assign out_43_1 = t_r43_c1_12 >> 4;

  assign t_r43_c2_0 = p_42_2 << 1;
  assign t_r43_c2_1 = p_43_1 << 1;
  assign t_r43_c2_2 = p_43_2 << 2;
  assign t_r43_c2_3 = p_43_3 << 1;
  assign t_r43_c2_4 = p_44_2 << 1;
  assign t_r43_c2_5 = t_r43_c2_0 + p_42_1;
  assign t_r43_c2_6 = t_r43_c2_1 + p_42_3;
  assign t_r43_c2_7 = t_r43_c2_2 + t_r43_c2_3;
  assign t_r43_c2_8 = t_r43_c2_4 + p_44_1;
  assign t_r43_c2_9 = t_r43_c2_5 + t_r43_c2_6;
  assign t_r43_c2_10 = t_r43_c2_7 + t_r43_c2_8;
  assign t_r43_c2_11 = t_r43_c2_9 + t_r43_c2_10;
  assign t_r43_c2_12 = t_r43_c2_11 + p_44_3;
  assign out_43_2 = t_r43_c2_12 >> 4;

  assign t_r43_c3_0 = p_42_3 << 1;
  assign t_r43_c3_1 = p_43_2 << 1;
  assign t_r43_c3_2 = p_43_3 << 2;
  assign t_r43_c3_3 = p_43_4 << 1;
  assign t_r43_c3_4 = p_44_3 << 1;
  assign t_r43_c3_5 = t_r43_c3_0 + p_42_2;
  assign t_r43_c3_6 = t_r43_c3_1 + p_42_4;
  assign t_r43_c3_7 = t_r43_c3_2 + t_r43_c3_3;
  assign t_r43_c3_8 = t_r43_c3_4 + p_44_2;
  assign t_r43_c3_9 = t_r43_c3_5 + t_r43_c3_6;
  assign t_r43_c3_10 = t_r43_c3_7 + t_r43_c3_8;
  assign t_r43_c3_11 = t_r43_c3_9 + t_r43_c3_10;
  assign t_r43_c3_12 = t_r43_c3_11 + p_44_4;
  assign out_43_3 = t_r43_c3_12 >> 4;

  assign t_r43_c4_0 = p_42_4 << 1;
  assign t_r43_c4_1 = p_43_3 << 1;
  assign t_r43_c4_2 = p_43_4 << 2;
  assign t_r43_c4_3 = p_43_5 << 1;
  assign t_r43_c4_4 = p_44_4 << 1;
  assign t_r43_c4_5 = t_r43_c4_0 + p_42_3;
  assign t_r43_c4_6 = t_r43_c4_1 + p_42_5;
  assign t_r43_c4_7 = t_r43_c4_2 + t_r43_c4_3;
  assign t_r43_c4_8 = t_r43_c4_4 + p_44_3;
  assign t_r43_c4_9 = t_r43_c4_5 + t_r43_c4_6;
  assign t_r43_c4_10 = t_r43_c4_7 + t_r43_c4_8;
  assign t_r43_c4_11 = t_r43_c4_9 + t_r43_c4_10;
  assign t_r43_c4_12 = t_r43_c4_11 + p_44_5;
  assign out_43_4 = t_r43_c4_12 >> 4;

  assign t_r43_c5_0 = p_42_5 << 1;
  assign t_r43_c5_1 = p_43_4 << 1;
  assign t_r43_c5_2 = p_43_5 << 2;
  assign t_r43_c5_3 = p_43_6 << 1;
  assign t_r43_c5_4 = p_44_5 << 1;
  assign t_r43_c5_5 = t_r43_c5_0 + p_42_4;
  assign t_r43_c5_6 = t_r43_c5_1 + p_42_6;
  assign t_r43_c5_7 = t_r43_c5_2 + t_r43_c5_3;
  assign t_r43_c5_8 = t_r43_c5_4 + p_44_4;
  assign t_r43_c5_9 = t_r43_c5_5 + t_r43_c5_6;
  assign t_r43_c5_10 = t_r43_c5_7 + t_r43_c5_8;
  assign t_r43_c5_11 = t_r43_c5_9 + t_r43_c5_10;
  assign t_r43_c5_12 = t_r43_c5_11 + p_44_6;
  assign out_43_5 = t_r43_c5_12 >> 4;

  assign t_r43_c6_0 = p_42_6 << 1;
  assign t_r43_c6_1 = p_43_5 << 1;
  assign t_r43_c6_2 = p_43_6 << 2;
  assign t_r43_c6_3 = p_43_7 << 1;
  assign t_r43_c6_4 = p_44_6 << 1;
  assign t_r43_c6_5 = t_r43_c6_0 + p_42_5;
  assign t_r43_c6_6 = t_r43_c6_1 + p_42_7;
  assign t_r43_c6_7 = t_r43_c6_2 + t_r43_c6_3;
  assign t_r43_c6_8 = t_r43_c6_4 + p_44_5;
  assign t_r43_c6_9 = t_r43_c6_5 + t_r43_c6_6;
  assign t_r43_c6_10 = t_r43_c6_7 + t_r43_c6_8;
  assign t_r43_c6_11 = t_r43_c6_9 + t_r43_c6_10;
  assign t_r43_c6_12 = t_r43_c6_11 + p_44_7;
  assign out_43_6 = t_r43_c6_12 >> 4;

  assign t_r43_c7_0 = p_42_7 << 1;
  assign t_r43_c7_1 = p_43_6 << 1;
  assign t_r43_c7_2 = p_43_7 << 2;
  assign t_r43_c7_3 = p_43_8 << 1;
  assign t_r43_c7_4 = p_44_7 << 1;
  assign t_r43_c7_5 = t_r43_c7_0 + p_42_6;
  assign t_r43_c7_6 = t_r43_c7_1 + p_42_8;
  assign t_r43_c7_7 = t_r43_c7_2 + t_r43_c7_3;
  assign t_r43_c7_8 = t_r43_c7_4 + p_44_6;
  assign t_r43_c7_9 = t_r43_c7_5 + t_r43_c7_6;
  assign t_r43_c7_10 = t_r43_c7_7 + t_r43_c7_8;
  assign t_r43_c7_11 = t_r43_c7_9 + t_r43_c7_10;
  assign t_r43_c7_12 = t_r43_c7_11 + p_44_8;
  assign out_43_7 = t_r43_c7_12 >> 4;

  assign t_r43_c8_0 = p_42_8 << 1;
  assign t_r43_c8_1 = p_43_7 << 1;
  assign t_r43_c8_2 = p_43_8 << 2;
  assign t_r43_c8_3 = p_43_9 << 1;
  assign t_r43_c8_4 = p_44_8 << 1;
  assign t_r43_c8_5 = t_r43_c8_0 + p_42_7;
  assign t_r43_c8_6 = t_r43_c8_1 + p_42_9;
  assign t_r43_c8_7 = t_r43_c8_2 + t_r43_c8_3;
  assign t_r43_c8_8 = t_r43_c8_4 + p_44_7;
  assign t_r43_c8_9 = t_r43_c8_5 + t_r43_c8_6;
  assign t_r43_c8_10 = t_r43_c8_7 + t_r43_c8_8;
  assign t_r43_c8_11 = t_r43_c8_9 + t_r43_c8_10;
  assign t_r43_c8_12 = t_r43_c8_11 + p_44_9;
  assign out_43_8 = t_r43_c8_12 >> 4;

  assign t_r43_c9_0 = p_42_9 << 1;
  assign t_r43_c9_1 = p_43_8 << 1;
  assign t_r43_c9_2 = p_43_9 << 2;
  assign t_r43_c9_3 = p_43_10 << 1;
  assign t_r43_c9_4 = p_44_9 << 1;
  assign t_r43_c9_5 = t_r43_c9_0 + p_42_8;
  assign t_r43_c9_6 = t_r43_c9_1 + p_42_10;
  assign t_r43_c9_7 = t_r43_c9_2 + t_r43_c9_3;
  assign t_r43_c9_8 = t_r43_c9_4 + p_44_8;
  assign t_r43_c9_9 = t_r43_c9_5 + t_r43_c9_6;
  assign t_r43_c9_10 = t_r43_c9_7 + t_r43_c9_8;
  assign t_r43_c9_11 = t_r43_c9_9 + t_r43_c9_10;
  assign t_r43_c9_12 = t_r43_c9_11 + p_44_10;
  assign out_43_9 = t_r43_c9_12 >> 4;

  assign t_r43_c10_0 = p_42_10 << 1;
  assign t_r43_c10_1 = p_43_9 << 1;
  assign t_r43_c10_2 = p_43_10 << 2;
  assign t_r43_c10_3 = p_43_11 << 1;
  assign t_r43_c10_4 = p_44_10 << 1;
  assign t_r43_c10_5 = t_r43_c10_0 + p_42_9;
  assign t_r43_c10_6 = t_r43_c10_1 + p_42_11;
  assign t_r43_c10_7 = t_r43_c10_2 + t_r43_c10_3;
  assign t_r43_c10_8 = t_r43_c10_4 + p_44_9;
  assign t_r43_c10_9 = t_r43_c10_5 + t_r43_c10_6;
  assign t_r43_c10_10 = t_r43_c10_7 + t_r43_c10_8;
  assign t_r43_c10_11 = t_r43_c10_9 + t_r43_c10_10;
  assign t_r43_c10_12 = t_r43_c10_11 + p_44_11;
  assign out_43_10 = t_r43_c10_12 >> 4;

  assign t_r43_c11_0 = p_42_11 << 1;
  assign t_r43_c11_1 = p_43_10 << 1;
  assign t_r43_c11_2 = p_43_11 << 2;
  assign t_r43_c11_3 = p_43_12 << 1;
  assign t_r43_c11_4 = p_44_11 << 1;
  assign t_r43_c11_5 = t_r43_c11_0 + p_42_10;
  assign t_r43_c11_6 = t_r43_c11_1 + p_42_12;
  assign t_r43_c11_7 = t_r43_c11_2 + t_r43_c11_3;
  assign t_r43_c11_8 = t_r43_c11_4 + p_44_10;
  assign t_r43_c11_9 = t_r43_c11_5 + t_r43_c11_6;
  assign t_r43_c11_10 = t_r43_c11_7 + t_r43_c11_8;
  assign t_r43_c11_11 = t_r43_c11_9 + t_r43_c11_10;
  assign t_r43_c11_12 = t_r43_c11_11 + p_44_12;
  assign out_43_11 = t_r43_c11_12 >> 4;

  assign t_r43_c12_0 = p_42_12 << 1;
  assign t_r43_c12_1 = p_43_11 << 1;
  assign t_r43_c12_2 = p_43_12 << 2;
  assign t_r43_c12_3 = p_43_13 << 1;
  assign t_r43_c12_4 = p_44_12 << 1;
  assign t_r43_c12_5 = t_r43_c12_0 + p_42_11;
  assign t_r43_c12_6 = t_r43_c12_1 + p_42_13;
  assign t_r43_c12_7 = t_r43_c12_2 + t_r43_c12_3;
  assign t_r43_c12_8 = t_r43_c12_4 + p_44_11;
  assign t_r43_c12_9 = t_r43_c12_5 + t_r43_c12_6;
  assign t_r43_c12_10 = t_r43_c12_7 + t_r43_c12_8;
  assign t_r43_c12_11 = t_r43_c12_9 + t_r43_c12_10;
  assign t_r43_c12_12 = t_r43_c12_11 + p_44_13;
  assign out_43_12 = t_r43_c12_12 >> 4;

  assign t_r43_c13_0 = p_42_13 << 1;
  assign t_r43_c13_1 = p_43_12 << 1;
  assign t_r43_c13_2 = p_43_13 << 2;
  assign t_r43_c13_3 = p_43_14 << 1;
  assign t_r43_c13_4 = p_44_13 << 1;
  assign t_r43_c13_5 = t_r43_c13_0 + p_42_12;
  assign t_r43_c13_6 = t_r43_c13_1 + p_42_14;
  assign t_r43_c13_7 = t_r43_c13_2 + t_r43_c13_3;
  assign t_r43_c13_8 = t_r43_c13_4 + p_44_12;
  assign t_r43_c13_9 = t_r43_c13_5 + t_r43_c13_6;
  assign t_r43_c13_10 = t_r43_c13_7 + t_r43_c13_8;
  assign t_r43_c13_11 = t_r43_c13_9 + t_r43_c13_10;
  assign t_r43_c13_12 = t_r43_c13_11 + p_44_14;
  assign out_43_13 = t_r43_c13_12 >> 4;

  assign t_r43_c14_0 = p_42_14 << 1;
  assign t_r43_c14_1 = p_43_13 << 1;
  assign t_r43_c14_2 = p_43_14 << 2;
  assign t_r43_c14_3 = p_43_15 << 1;
  assign t_r43_c14_4 = p_44_14 << 1;
  assign t_r43_c14_5 = t_r43_c14_0 + p_42_13;
  assign t_r43_c14_6 = t_r43_c14_1 + p_42_15;
  assign t_r43_c14_7 = t_r43_c14_2 + t_r43_c14_3;
  assign t_r43_c14_8 = t_r43_c14_4 + p_44_13;
  assign t_r43_c14_9 = t_r43_c14_5 + t_r43_c14_6;
  assign t_r43_c14_10 = t_r43_c14_7 + t_r43_c14_8;
  assign t_r43_c14_11 = t_r43_c14_9 + t_r43_c14_10;
  assign t_r43_c14_12 = t_r43_c14_11 + p_44_15;
  assign out_43_14 = t_r43_c14_12 >> 4;

  assign t_r43_c15_0 = p_42_15 << 1;
  assign t_r43_c15_1 = p_43_14 << 1;
  assign t_r43_c15_2 = p_43_15 << 2;
  assign t_r43_c15_3 = p_43_16 << 1;
  assign t_r43_c15_4 = p_44_15 << 1;
  assign t_r43_c15_5 = t_r43_c15_0 + p_42_14;
  assign t_r43_c15_6 = t_r43_c15_1 + p_42_16;
  assign t_r43_c15_7 = t_r43_c15_2 + t_r43_c15_3;
  assign t_r43_c15_8 = t_r43_c15_4 + p_44_14;
  assign t_r43_c15_9 = t_r43_c15_5 + t_r43_c15_6;
  assign t_r43_c15_10 = t_r43_c15_7 + t_r43_c15_8;
  assign t_r43_c15_11 = t_r43_c15_9 + t_r43_c15_10;
  assign t_r43_c15_12 = t_r43_c15_11 + p_44_16;
  assign out_43_15 = t_r43_c15_12 >> 4;

  assign t_r43_c16_0 = p_42_16 << 1;
  assign t_r43_c16_1 = p_43_15 << 1;
  assign t_r43_c16_2 = p_43_16 << 2;
  assign t_r43_c16_3 = p_43_17 << 1;
  assign t_r43_c16_4 = p_44_16 << 1;
  assign t_r43_c16_5 = t_r43_c16_0 + p_42_15;
  assign t_r43_c16_6 = t_r43_c16_1 + p_42_17;
  assign t_r43_c16_7 = t_r43_c16_2 + t_r43_c16_3;
  assign t_r43_c16_8 = t_r43_c16_4 + p_44_15;
  assign t_r43_c16_9 = t_r43_c16_5 + t_r43_c16_6;
  assign t_r43_c16_10 = t_r43_c16_7 + t_r43_c16_8;
  assign t_r43_c16_11 = t_r43_c16_9 + t_r43_c16_10;
  assign t_r43_c16_12 = t_r43_c16_11 + p_44_17;
  assign out_43_16 = t_r43_c16_12 >> 4;

  assign t_r43_c17_0 = p_42_17 << 1;
  assign t_r43_c17_1 = p_43_16 << 1;
  assign t_r43_c17_2 = p_43_17 << 2;
  assign t_r43_c17_3 = p_43_18 << 1;
  assign t_r43_c17_4 = p_44_17 << 1;
  assign t_r43_c17_5 = t_r43_c17_0 + p_42_16;
  assign t_r43_c17_6 = t_r43_c17_1 + p_42_18;
  assign t_r43_c17_7 = t_r43_c17_2 + t_r43_c17_3;
  assign t_r43_c17_8 = t_r43_c17_4 + p_44_16;
  assign t_r43_c17_9 = t_r43_c17_5 + t_r43_c17_6;
  assign t_r43_c17_10 = t_r43_c17_7 + t_r43_c17_8;
  assign t_r43_c17_11 = t_r43_c17_9 + t_r43_c17_10;
  assign t_r43_c17_12 = t_r43_c17_11 + p_44_18;
  assign out_43_17 = t_r43_c17_12 >> 4;

  assign t_r43_c18_0 = p_42_18 << 1;
  assign t_r43_c18_1 = p_43_17 << 1;
  assign t_r43_c18_2 = p_43_18 << 2;
  assign t_r43_c18_3 = p_43_19 << 1;
  assign t_r43_c18_4 = p_44_18 << 1;
  assign t_r43_c18_5 = t_r43_c18_0 + p_42_17;
  assign t_r43_c18_6 = t_r43_c18_1 + p_42_19;
  assign t_r43_c18_7 = t_r43_c18_2 + t_r43_c18_3;
  assign t_r43_c18_8 = t_r43_c18_4 + p_44_17;
  assign t_r43_c18_9 = t_r43_c18_5 + t_r43_c18_6;
  assign t_r43_c18_10 = t_r43_c18_7 + t_r43_c18_8;
  assign t_r43_c18_11 = t_r43_c18_9 + t_r43_c18_10;
  assign t_r43_c18_12 = t_r43_c18_11 + p_44_19;
  assign out_43_18 = t_r43_c18_12 >> 4;

  assign t_r43_c19_0 = p_42_19 << 1;
  assign t_r43_c19_1 = p_43_18 << 1;
  assign t_r43_c19_2 = p_43_19 << 2;
  assign t_r43_c19_3 = p_43_20 << 1;
  assign t_r43_c19_4 = p_44_19 << 1;
  assign t_r43_c19_5 = t_r43_c19_0 + p_42_18;
  assign t_r43_c19_6 = t_r43_c19_1 + p_42_20;
  assign t_r43_c19_7 = t_r43_c19_2 + t_r43_c19_3;
  assign t_r43_c19_8 = t_r43_c19_4 + p_44_18;
  assign t_r43_c19_9 = t_r43_c19_5 + t_r43_c19_6;
  assign t_r43_c19_10 = t_r43_c19_7 + t_r43_c19_8;
  assign t_r43_c19_11 = t_r43_c19_9 + t_r43_c19_10;
  assign t_r43_c19_12 = t_r43_c19_11 + p_44_20;
  assign out_43_19 = t_r43_c19_12 >> 4;

  assign t_r43_c20_0 = p_42_20 << 1;
  assign t_r43_c20_1 = p_43_19 << 1;
  assign t_r43_c20_2 = p_43_20 << 2;
  assign t_r43_c20_3 = p_43_21 << 1;
  assign t_r43_c20_4 = p_44_20 << 1;
  assign t_r43_c20_5 = t_r43_c20_0 + p_42_19;
  assign t_r43_c20_6 = t_r43_c20_1 + p_42_21;
  assign t_r43_c20_7 = t_r43_c20_2 + t_r43_c20_3;
  assign t_r43_c20_8 = t_r43_c20_4 + p_44_19;
  assign t_r43_c20_9 = t_r43_c20_5 + t_r43_c20_6;
  assign t_r43_c20_10 = t_r43_c20_7 + t_r43_c20_8;
  assign t_r43_c20_11 = t_r43_c20_9 + t_r43_c20_10;
  assign t_r43_c20_12 = t_r43_c20_11 + p_44_21;
  assign out_43_20 = t_r43_c20_12 >> 4;

  assign t_r43_c21_0 = p_42_21 << 1;
  assign t_r43_c21_1 = p_43_20 << 1;
  assign t_r43_c21_2 = p_43_21 << 2;
  assign t_r43_c21_3 = p_43_22 << 1;
  assign t_r43_c21_4 = p_44_21 << 1;
  assign t_r43_c21_5 = t_r43_c21_0 + p_42_20;
  assign t_r43_c21_6 = t_r43_c21_1 + p_42_22;
  assign t_r43_c21_7 = t_r43_c21_2 + t_r43_c21_3;
  assign t_r43_c21_8 = t_r43_c21_4 + p_44_20;
  assign t_r43_c21_9 = t_r43_c21_5 + t_r43_c21_6;
  assign t_r43_c21_10 = t_r43_c21_7 + t_r43_c21_8;
  assign t_r43_c21_11 = t_r43_c21_9 + t_r43_c21_10;
  assign t_r43_c21_12 = t_r43_c21_11 + p_44_22;
  assign out_43_21 = t_r43_c21_12 >> 4;

  assign t_r43_c22_0 = p_42_22 << 1;
  assign t_r43_c22_1 = p_43_21 << 1;
  assign t_r43_c22_2 = p_43_22 << 2;
  assign t_r43_c22_3 = p_43_23 << 1;
  assign t_r43_c22_4 = p_44_22 << 1;
  assign t_r43_c22_5 = t_r43_c22_0 + p_42_21;
  assign t_r43_c22_6 = t_r43_c22_1 + p_42_23;
  assign t_r43_c22_7 = t_r43_c22_2 + t_r43_c22_3;
  assign t_r43_c22_8 = t_r43_c22_4 + p_44_21;
  assign t_r43_c22_9 = t_r43_c22_5 + t_r43_c22_6;
  assign t_r43_c22_10 = t_r43_c22_7 + t_r43_c22_8;
  assign t_r43_c22_11 = t_r43_c22_9 + t_r43_c22_10;
  assign t_r43_c22_12 = t_r43_c22_11 + p_44_23;
  assign out_43_22 = t_r43_c22_12 >> 4;

  assign t_r43_c23_0 = p_42_23 << 1;
  assign t_r43_c23_1 = p_43_22 << 1;
  assign t_r43_c23_2 = p_43_23 << 2;
  assign t_r43_c23_3 = p_43_24 << 1;
  assign t_r43_c23_4 = p_44_23 << 1;
  assign t_r43_c23_5 = t_r43_c23_0 + p_42_22;
  assign t_r43_c23_6 = t_r43_c23_1 + p_42_24;
  assign t_r43_c23_7 = t_r43_c23_2 + t_r43_c23_3;
  assign t_r43_c23_8 = t_r43_c23_4 + p_44_22;
  assign t_r43_c23_9 = t_r43_c23_5 + t_r43_c23_6;
  assign t_r43_c23_10 = t_r43_c23_7 + t_r43_c23_8;
  assign t_r43_c23_11 = t_r43_c23_9 + t_r43_c23_10;
  assign t_r43_c23_12 = t_r43_c23_11 + p_44_24;
  assign out_43_23 = t_r43_c23_12 >> 4;

  assign t_r43_c24_0 = p_42_24 << 1;
  assign t_r43_c24_1 = p_43_23 << 1;
  assign t_r43_c24_2 = p_43_24 << 2;
  assign t_r43_c24_3 = p_43_25 << 1;
  assign t_r43_c24_4 = p_44_24 << 1;
  assign t_r43_c24_5 = t_r43_c24_0 + p_42_23;
  assign t_r43_c24_6 = t_r43_c24_1 + p_42_25;
  assign t_r43_c24_7 = t_r43_c24_2 + t_r43_c24_3;
  assign t_r43_c24_8 = t_r43_c24_4 + p_44_23;
  assign t_r43_c24_9 = t_r43_c24_5 + t_r43_c24_6;
  assign t_r43_c24_10 = t_r43_c24_7 + t_r43_c24_8;
  assign t_r43_c24_11 = t_r43_c24_9 + t_r43_c24_10;
  assign t_r43_c24_12 = t_r43_c24_11 + p_44_25;
  assign out_43_24 = t_r43_c24_12 >> 4;

  assign t_r43_c25_0 = p_42_25 << 1;
  assign t_r43_c25_1 = p_43_24 << 1;
  assign t_r43_c25_2 = p_43_25 << 2;
  assign t_r43_c25_3 = p_43_26 << 1;
  assign t_r43_c25_4 = p_44_25 << 1;
  assign t_r43_c25_5 = t_r43_c25_0 + p_42_24;
  assign t_r43_c25_6 = t_r43_c25_1 + p_42_26;
  assign t_r43_c25_7 = t_r43_c25_2 + t_r43_c25_3;
  assign t_r43_c25_8 = t_r43_c25_4 + p_44_24;
  assign t_r43_c25_9 = t_r43_c25_5 + t_r43_c25_6;
  assign t_r43_c25_10 = t_r43_c25_7 + t_r43_c25_8;
  assign t_r43_c25_11 = t_r43_c25_9 + t_r43_c25_10;
  assign t_r43_c25_12 = t_r43_c25_11 + p_44_26;
  assign out_43_25 = t_r43_c25_12 >> 4;

  assign t_r43_c26_0 = p_42_26 << 1;
  assign t_r43_c26_1 = p_43_25 << 1;
  assign t_r43_c26_2 = p_43_26 << 2;
  assign t_r43_c26_3 = p_43_27 << 1;
  assign t_r43_c26_4 = p_44_26 << 1;
  assign t_r43_c26_5 = t_r43_c26_0 + p_42_25;
  assign t_r43_c26_6 = t_r43_c26_1 + p_42_27;
  assign t_r43_c26_7 = t_r43_c26_2 + t_r43_c26_3;
  assign t_r43_c26_8 = t_r43_c26_4 + p_44_25;
  assign t_r43_c26_9 = t_r43_c26_5 + t_r43_c26_6;
  assign t_r43_c26_10 = t_r43_c26_7 + t_r43_c26_8;
  assign t_r43_c26_11 = t_r43_c26_9 + t_r43_c26_10;
  assign t_r43_c26_12 = t_r43_c26_11 + p_44_27;
  assign out_43_26 = t_r43_c26_12 >> 4;

  assign t_r43_c27_0 = p_42_27 << 1;
  assign t_r43_c27_1 = p_43_26 << 1;
  assign t_r43_c27_2 = p_43_27 << 2;
  assign t_r43_c27_3 = p_43_28 << 1;
  assign t_r43_c27_4 = p_44_27 << 1;
  assign t_r43_c27_5 = t_r43_c27_0 + p_42_26;
  assign t_r43_c27_6 = t_r43_c27_1 + p_42_28;
  assign t_r43_c27_7 = t_r43_c27_2 + t_r43_c27_3;
  assign t_r43_c27_8 = t_r43_c27_4 + p_44_26;
  assign t_r43_c27_9 = t_r43_c27_5 + t_r43_c27_6;
  assign t_r43_c27_10 = t_r43_c27_7 + t_r43_c27_8;
  assign t_r43_c27_11 = t_r43_c27_9 + t_r43_c27_10;
  assign t_r43_c27_12 = t_r43_c27_11 + p_44_28;
  assign out_43_27 = t_r43_c27_12 >> 4;

  assign t_r43_c28_0 = p_42_28 << 1;
  assign t_r43_c28_1 = p_43_27 << 1;
  assign t_r43_c28_2 = p_43_28 << 2;
  assign t_r43_c28_3 = p_43_29 << 1;
  assign t_r43_c28_4 = p_44_28 << 1;
  assign t_r43_c28_5 = t_r43_c28_0 + p_42_27;
  assign t_r43_c28_6 = t_r43_c28_1 + p_42_29;
  assign t_r43_c28_7 = t_r43_c28_2 + t_r43_c28_3;
  assign t_r43_c28_8 = t_r43_c28_4 + p_44_27;
  assign t_r43_c28_9 = t_r43_c28_5 + t_r43_c28_6;
  assign t_r43_c28_10 = t_r43_c28_7 + t_r43_c28_8;
  assign t_r43_c28_11 = t_r43_c28_9 + t_r43_c28_10;
  assign t_r43_c28_12 = t_r43_c28_11 + p_44_29;
  assign out_43_28 = t_r43_c28_12 >> 4;

  assign t_r43_c29_0 = p_42_29 << 1;
  assign t_r43_c29_1 = p_43_28 << 1;
  assign t_r43_c29_2 = p_43_29 << 2;
  assign t_r43_c29_3 = p_43_30 << 1;
  assign t_r43_c29_4 = p_44_29 << 1;
  assign t_r43_c29_5 = t_r43_c29_0 + p_42_28;
  assign t_r43_c29_6 = t_r43_c29_1 + p_42_30;
  assign t_r43_c29_7 = t_r43_c29_2 + t_r43_c29_3;
  assign t_r43_c29_8 = t_r43_c29_4 + p_44_28;
  assign t_r43_c29_9 = t_r43_c29_5 + t_r43_c29_6;
  assign t_r43_c29_10 = t_r43_c29_7 + t_r43_c29_8;
  assign t_r43_c29_11 = t_r43_c29_9 + t_r43_c29_10;
  assign t_r43_c29_12 = t_r43_c29_11 + p_44_30;
  assign out_43_29 = t_r43_c29_12 >> 4;

  assign t_r43_c30_0 = p_42_30 << 1;
  assign t_r43_c30_1 = p_43_29 << 1;
  assign t_r43_c30_2 = p_43_30 << 2;
  assign t_r43_c30_3 = p_43_31 << 1;
  assign t_r43_c30_4 = p_44_30 << 1;
  assign t_r43_c30_5 = t_r43_c30_0 + p_42_29;
  assign t_r43_c30_6 = t_r43_c30_1 + p_42_31;
  assign t_r43_c30_7 = t_r43_c30_2 + t_r43_c30_3;
  assign t_r43_c30_8 = t_r43_c30_4 + p_44_29;
  assign t_r43_c30_9 = t_r43_c30_5 + t_r43_c30_6;
  assign t_r43_c30_10 = t_r43_c30_7 + t_r43_c30_8;
  assign t_r43_c30_11 = t_r43_c30_9 + t_r43_c30_10;
  assign t_r43_c30_12 = t_r43_c30_11 + p_44_31;
  assign out_43_30 = t_r43_c30_12 >> 4;

  assign t_r43_c31_0 = p_42_31 << 1;
  assign t_r43_c31_1 = p_43_30 << 1;
  assign t_r43_c31_2 = p_43_31 << 2;
  assign t_r43_c31_3 = p_43_32 << 1;
  assign t_r43_c31_4 = p_44_31 << 1;
  assign t_r43_c31_5 = t_r43_c31_0 + p_42_30;
  assign t_r43_c31_6 = t_r43_c31_1 + p_42_32;
  assign t_r43_c31_7 = t_r43_c31_2 + t_r43_c31_3;
  assign t_r43_c31_8 = t_r43_c31_4 + p_44_30;
  assign t_r43_c31_9 = t_r43_c31_5 + t_r43_c31_6;
  assign t_r43_c31_10 = t_r43_c31_7 + t_r43_c31_8;
  assign t_r43_c31_11 = t_r43_c31_9 + t_r43_c31_10;
  assign t_r43_c31_12 = t_r43_c31_11 + p_44_32;
  assign out_43_31 = t_r43_c31_12 >> 4;

  assign t_r43_c32_0 = p_42_32 << 1;
  assign t_r43_c32_1 = p_43_31 << 1;
  assign t_r43_c32_2 = p_43_32 << 2;
  assign t_r43_c32_3 = p_43_33 << 1;
  assign t_r43_c32_4 = p_44_32 << 1;
  assign t_r43_c32_5 = t_r43_c32_0 + p_42_31;
  assign t_r43_c32_6 = t_r43_c32_1 + p_42_33;
  assign t_r43_c32_7 = t_r43_c32_2 + t_r43_c32_3;
  assign t_r43_c32_8 = t_r43_c32_4 + p_44_31;
  assign t_r43_c32_9 = t_r43_c32_5 + t_r43_c32_6;
  assign t_r43_c32_10 = t_r43_c32_7 + t_r43_c32_8;
  assign t_r43_c32_11 = t_r43_c32_9 + t_r43_c32_10;
  assign t_r43_c32_12 = t_r43_c32_11 + p_44_33;
  assign out_43_32 = t_r43_c32_12 >> 4;

  assign t_r43_c33_0 = p_42_33 << 1;
  assign t_r43_c33_1 = p_43_32 << 1;
  assign t_r43_c33_2 = p_43_33 << 2;
  assign t_r43_c33_3 = p_43_34 << 1;
  assign t_r43_c33_4 = p_44_33 << 1;
  assign t_r43_c33_5 = t_r43_c33_0 + p_42_32;
  assign t_r43_c33_6 = t_r43_c33_1 + p_42_34;
  assign t_r43_c33_7 = t_r43_c33_2 + t_r43_c33_3;
  assign t_r43_c33_8 = t_r43_c33_4 + p_44_32;
  assign t_r43_c33_9 = t_r43_c33_5 + t_r43_c33_6;
  assign t_r43_c33_10 = t_r43_c33_7 + t_r43_c33_8;
  assign t_r43_c33_11 = t_r43_c33_9 + t_r43_c33_10;
  assign t_r43_c33_12 = t_r43_c33_11 + p_44_34;
  assign out_43_33 = t_r43_c33_12 >> 4;

  assign t_r43_c34_0 = p_42_34 << 1;
  assign t_r43_c34_1 = p_43_33 << 1;
  assign t_r43_c34_2 = p_43_34 << 2;
  assign t_r43_c34_3 = p_43_35 << 1;
  assign t_r43_c34_4 = p_44_34 << 1;
  assign t_r43_c34_5 = t_r43_c34_0 + p_42_33;
  assign t_r43_c34_6 = t_r43_c34_1 + p_42_35;
  assign t_r43_c34_7 = t_r43_c34_2 + t_r43_c34_3;
  assign t_r43_c34_8 = t_r43_c34_4 + p_44_33;
  assign t_r43_c34_9 = t_r43_c34_5 + t_r43_c34_6;
  assign t_r43_c34_10 = t_r43_c34_7 + t_r43_c34_8;
  assign t_r43_c34_11 = t_r43_c34_9 + t_r43_c34_10;
  assign t_r43_c34_12 = t_r43_c34_11 + p_44_35;
  assign out_43_34 = t_r43_c34_12 >> 4;

  assign t_r43_c35_0 = p_42_35 << 1;
  assign t_r43_c35_1 = p_43_34 << 1;
  assign t_r43_c35_2 = p_43_35 << 2;
  assign t_r43_c35_3 = p_43_36 << 1;
  assign t_r43_c35_4 = p_44_35 << 1;
  assign t_r43_c35_5 = t_r43_c35_0 + p_42_34;
  assign t_r43_c35_6 = t_r43_c35_1 + p_42_36;
  assign t_r43_c35_7 = t_r43_c35_2 + t_r43_c35_3;
  assign t_r43_c35_8 = t_r43_c35_4 + p_44_34;
  assign t_r43_c35_9 = t_r43_c35_5 + t_r43_c35_6;
  assign t_r43_c35_10 = t_r43_c35_7 + t_r43_c35_8;
  assign t_r43_c35_11 = t_r43_c35_9 + t_r43_c35_10;
  assign t_r43_c35_12 = t_r43_c35_11 + p_44_36;
  assign out_43_35 = t_r43_c35_12 >> 4;

  assign t_r43_c36_0 = p_42_36 << 1;
  assign t_r43_c36_1 = p_43_35 << 1;
  assign t_r43_c36_2 = p_43_36 << 2;
  assign t_r43_c36_3 = p_43_37 << 1;
  assign t_r43_c36_4 = p_44_36 << 1;
  assign t_r43_c36_5 = t_r43_c36_0 + p_42_35;
  assign t_r43_c36_6 = t_r43_c36_1 + p_42_37;
  assign t_r43_c36_7 = t_r43_c36_2 + t_r43_c36_3;
  assign t_r43_c36_8 = t_r43_c36_4 + p_44_35;
  assign t_r43_c36_9 = t_r43_c36_5 + t_r43_c36_6;
  assign t_r43_c36_10 = t_r43_c36_7 + t_r43_c36_8;
  assign t_r43_c36_11 = t_r43_c36_9 + t_r43_c36_10;
  assign t_r43_c36_12 = t_r43_c36_11 + p_44_37;
  assign out_43_36 = t_r43_c36_12 >> 4;

  assign t_r43_c37_0 = p_42_37 << 1;
  assign t_r43_c37_1 = p_43_36 << 1;
  assign t_r43_c37_2 = p_43_37 << 2;
  assign t_r43_c37_3 = p_43_38 << 1;
  assign t_r43_c37_4 = p_44_37 << 1;
  assign t_r43_c37_5 = t_r43_c37_0 + p_42_36;
  assign t_r43_c37_6 = t_r43_c37_1 + p_42_38;
  assign t_r43_c37_7 = t_r43_c37_2 + t_r43_c37_3;
  assign t_r43_c37_8 = t_r43_c37_4 + p_44_36;
  assign t_r43_c37_9 = t_r43_c37_5 + t_r43_c37_6;
  assign t_r43_c37_10 = t_r43_c37_7 + t_r43_c37_8;
  assign t_r43_c37_11 = t_r43_c37_9 + t_r43_c37_10;
  assign t_r43_c37_12 = t_r43_c37_11 + p_44_38;
  assign out_43_37 = t_r43_c37_12 >> 4;

  assign t_r43_c38_0 = p_42_38 << 1;
  assign t_r43_c38_1 = p_43_37 << 1;
  assign t_r43_c38_2 = p_43_38 << 2;
  assign t_r43_c38_3 = p_43_39 << 1;
  assign t_r43_c38_4 = p_44_38 << 1;
  assign t_r43_c38_5 = t_r43_c38_0 + p_42_37;
  assign t_r43_c38_6 = t_r43_c38_1 + p_42_39;
  assign t_r43_c38_7 = t_r43_c38_2 + t_r43_c38_3;
  assign t_r43_c38_8 = t_r43_c38_4 + p_44_37;
  assign t_r43_c38_9 = t_r43_c38_5 + t_r43_c38_6;
  assign t_r43_c38_10 = t_r43_c38_7 + t_r43_c38_8;
  assign t_r43_c38_11 = t_r43_c38_9 + t_r43_c38_10;
  assign t_r43_c38_12 = t_r43_c38_11 + p_44_39;
  assign out_43_38 = t_r43_c38_12 >> 4;

  assign t_r43_c39_0 = p_42_39 << 1;
  assign t_r43_c39_1 = p_43_38 << 1;
  assign t_r43_c39_2 = p_43_39 << 2;
  assign t_r43_c39_3 = p_43_40 << 1;
  assign t_r43_c39_4 = p_44_39 << 1;
  assign t_r43_c39_5 = t_r43_c39_0 + p_42_38;
  assign t_r43_c39_6 = t_r43_c39_1 + p_42_40;
  assign t_r43_c39_7 = t_r43_c39_2 + t_r43_c39_3;
  assign t_r43_c39_8 = t_r43_c39_4 + p_44_38;
  assign t_r43_c39_9 = t_r43_c39_5 + t_r43_c39_6;
  assign t_r43_c39_10 = t_r43_c39_7 + t_r43_c39_8;
  assign t_r43_c39_11 = t_r43_c39_9 + t_r43_c39_10;
  assign t_r43_c39_12 = t_r43_c39_11 + p_44_40;
  assign out_43_39 = t_r43_c39_12 >> 4;

  assign t_r43_c40_0 = p_42_40 << 1;
  assign t_r43_c40_1 = p_43_39 << 1;
  assign t_r43_c40_2 = p_43_40 << 2;
  assign t_r43_c40_3 = p_43_41 << 1;
  assign t_r43_c40_4 = p_44_40 << 1;
  assign t_r43_c40_5 = t_r43_c40_0 + p_42_39;
  assign t_r43_c40_6 = t_r43_c40_1 + p_42_41;
  assign t_r43_c40_7 = t_r43_c40_2 + t_r43_c40_3;
  assign t_r43_c40_8 = t_r43_c40_4 + p_44_39;
  assign t_r43_c40_9 = t_r43_c40_5 + t_r43_c40_6;
  assign t_r43_c40_10 = t_r43_c40_7 + t_r43_c40_8;
  assign t_r43_c40_11 = t_r43_c40_9 + t_r43_c40_10;
  assign t_r43_c40_12 = t_r43_c40_11 + p_44_41;
  assign out_43_40 = t_r43_c40_12 >> 4;

  assign t_r43_c41_0 = p_42_41 << 1;
  assign t_r43_c41_1 = p_43_40 << 1;
  assign t_r43_c41_2 = p_43_41 << 2;
  assign t_r43_c41_3 = p_43_42 << 1;
  assign t_r43_c41_4 = p_44_41 << 1;
  assign t_r43_c41_5 = t_r43_c41_0 + p_42_40;
  assign t_r43_c41_6 = t_r43_c41_1 + p_42_42;
  assign t_r43_c41_7 = t_r43_c41_2 + t_r43_c41_3;
  assign t_r43_c41_8 = t_r43_c41_4 + p_44_40;
  assign t_r43_c41_9 = t_r43_c41_5 + t_r43_c41_6;
  assign t_r43_c41_10 = t_r43_c41_7 + t_r43_c41_8;
  assign t_r43_c41_11 = t_r43_c41_9 + t_r43_c41_10;
  assign t_r43_c41_12 = t_r43_c41_11 + p_44_42;
  assign out_43_41 = t_r43_c41_12 >> 4;

  assign t_r43_c42_0 = p_42_42 << 1;
  assign t_r43_c42_1 = p_43_41 << 1;
  assign t_r43_c42_2 = p_43_42 << 2;
  assign t_r43_c42_3 = p_43_43 << 1;
  assign t_r43_c42_4 = p_44_42 << 1;
  assign t_r43_c42_5 = t_r43_c42_0 + p_42_41;
  assign t_r43_c42_6 = t_r43_c42_1 + p_42_43;
  assign t_r43_c42_7 = t_r43_c42_2 + t_r43_c42_3;
  assign t_r43_c42_8 = t_r43_c42_4 + p_44_41;
  assign t_r43_c42_9 = t_r43_c42_5 + t_r43_c42_6;
  assign t_r43_c42_10 = t_r43_c42_7 + t_r43_c42_8;
  assign t_r43_c42_11 = t_r43_c42_9 + t_r43_c42_10;
  assign t_r43_c42_12 = t_r43_c42_11 + p_44_43;
  assign out_43_42 = t_r43_c42_12 >> 4;

  assign t_r43_c43_0 = p_42_43 << 1;
  assign t_r43_c43_1 = p_43_42 << 1;
  assign t_r43_c43_2 = p_43_43 << 2;
  assign t_r43_c43_3 = p_43_44 << 1;
  assign t_r43_c43_4 = p_44_43 << 1;
  assign t_r43_c43_5 = t_r43_c43_0 + p_42_42;
  assign t_r43_c43_6 = t_r43_c43_1 + p_42_44;
  assign t_r43_c43_7 = t_r43_c43_2 + t_r43_c43_3;
  assign t_r43_c43_8 = t_r43_c43_4 + p_44_42;
  assign t_r43_c43_9 = t_r43_c43_5 + t_r43_c43_6;
  assign t_r43_c43_10 = t_r43_c43_7 + t_r43_c43_8;
  assign t_r43_c43_11 = t_r43_c43_9 + t_r43_c43_10;
  assign t_r43_c43_12 = t_r43_c43_11 + p_44_44;
  assign out_43_43 = t_r43_c43_12 >> 4;

  assign t_r43_c44_0 = p_42_44 << 1;
  assign t_r43_c44_1 = p_43_43 << 1;
  assign t_r43_c44_2 = p_43_44 << 2;
  assign t_r43_c44_3 = p_43_45 << 1;
  assign t_r43_c44_4 = p_44_44 << 1;
  assign t_r43_c44_5 = t_r43_c44_0 + p_42_43;
  assign t_r43_c44_6 = t_r43_c44_1 + p_42_45;
  assign t_r43_c44_7 = t_r43_c44_2 + t_r43_c44_3;
  assign t_r43_c44_8 = t_r43_c44_4 + p_44_43;
  assign t_r43_c44_9 = t_r43_c44_5 + t_r43_c44_6;
  assign t_r43_c44_10 = t_r43_c44_7 + t_r43_c44_8;
  assign t_r43_c44_11 = t_r43_c44_9 + t_r43_c44_10;
  assign t_r43_c44_12 = t_r43_c44_11 + p_44_45;
  assign out_43_44 = t_r43_c44_12 >> 4;

  assign t_r43_c45_0 = p_42_45 << 1;
  assign t_r43_c45_1 = p_43_44 << 1;
  assign t_r43_c45_2 = p_43_45 << 2;
  assign t_r43_c45_3 = p_43_46 << 1;
  assign t_r43_c45_4 = p_44_45 << 1;
  assign t_r43_c45_5 = t_r43_c45_0 + p_42_44;
  assign t_r43_c45_6 = t_r43_c45_1 + p_42_46;
  assign t_r43_c45_7 = t_r43_c45_2 + t_r43_c45_3;
  assign t_r43_c45_8 = t_r43_c45_4 + p_44_44;
  assign t_r43_c45_9 = t_r43_c45_5 + t_r43_c45_6;
  assign t_r43_c45_10 = t_r43_c45_7 + t_r43_c45_8;
  assign t_r43_c45_11 = t_r43_c45_9 + t_r43_c45_10;
  assign t_r43_c45_12 = t_r43_c45_11 + p_44_46;
  assign out_43_45 = t_r43_c45_12 >> 4;

  assign t_r43_c46_0 = p_42_46 << 1;
  assign t_r43_c46_1 = p_43_45 << 1;
  assign t_r43_c46_2 = p_43_46 << 2;
  assign t_r43_c46_3 = p_43_47 << 1;
  assign t_r43_c46_4 = p_44_46 << 1;
  assign t_r43_c46_5 = t_r43_c46_0 + p_42_45;
  assign t_r43_c46_6 = t_r43_c46_1 + p_42_47;
  assign t_r43_c46_7 = t_r43_c46_2 + t_r43_c46_3;
  assign t_r43_c46_8 = t_r43_c46_4 + p_44_45;
  assign t_r43_c46_9 = t_r43_c46_5 + t_r43_c46_6;
  assign t_r43_c46_10 = t_r43_c46_7 + t_r43_c46_8;
  assign t_r43_c46_11 = t_r43_c46_9 + t_r43_c46_10;
  assign t_r43_c46_12 = t_r43_c46_11 + p_44_47;
  assign out_43_46 = t_r43_c46_12 >> 4;

  assign t_r43_c47_0 = p_42_47 << 1;
  assign t_r43_c47_1 = p_43_46 << 1;
  assign t_r43_c47_2 = p_43_47 << 2;
  assign t_r43_c47_3 = p_43_48 << 1;
  assign t_r43_c47_4 = p_44_47 << 1;
  assign t_r43_c47_5 = t_r43_c47_0 + p_42_46;
  assign t_r43_c47_6 = t_r43_c47_1 + p_42_48;
  assign t_r43_c47_7 = t_r43_c47_2 + t_r43_c47_3;
  assign t_r43_c47_8 = t_r43_c47_4 + p_44_46;
  assign t_r43_c47_9 = t_r43_c47_5 + t_r43_c47_6;
  assign t_r43_c47_10 = t_r43_c47_7 + t_r43_c47_8;
  assign t_r43_c47_11 = t_r43_c47_9 + t_r43_c47_10;
  assign t_r43_c47_12 = t_r43_c47_11 + p_44_48;
  assign out_43_47 = t_r43_c47_12 >> 4;

  assign t_r43_c48_0 = p_42_48 << 1;
  assign t_r43_c48_1 = p_43_47 << 1;
  assign t_r43_c48_2 = p_43_48 << 2;
  assign t_r43_c48_3 = p_43_49 << 1;
  assign t_r43_c48_4 = p_44_48 << 1;
  assign t_r43_c48_5 = t_r43_c48_0 + p_42_47;
  assign t_r43_c48_6 = t_r43_c48_1 + p_42_49;
  assign t_r43_c48_7 = t_r43_c48_2 + t_r43_c48_3;
  assign t_r43_c48_8 = t_r43_c48_4 + p_44_47;
  assign t_r43_c48_9 = t_r43_c48_5 + t_r43_c48_6;
  assign t_r43_c48_10 = t_r43_c48_7 + t_r43_c48_8;
  assign t_r43_c48_11 = t_r43_c48_9 + t_r43_c48_10;
  assign t_r43_c48_12 = t_r43_c48_11 + p_44_49;
  assign out_43_48 = t_r43_c48_12 >> 4;

  assign t_r43_c49_0 = p_42_49 << 1;
  assign t_r43_c49_1 = p_43_48 << 1;
  assign t_r43_c49_2 = p_43_49 << 2;
  assign t_r43_c49_3 = p_43_50 << 1;
  assign t_r43_c49_4 = p_44_49 << 1;
  assign t_r43_c49_5 = t_r43_c49_0 + p_42_48;
  assign t_r43_c49_6 = t_r43_c49_1 + p_42_50;
  assign t_r43_c49_7 = t_r43_c49_2 + t_r43_c49_3;
  assign t_r43_c49_8 = t_r43_c49_4 + p_44_48;
  assign t_r43_c49_9 = t_r43_c49_5 + t_r43_c49_6;
  assign t_r43_c49_10 = t_r43_c49_7 + t_r43_c49_8;
  assign t_r43_c49_11 = t_r43_c49_9 + t_r43_c49_10;
  assign t_r43_c49_12 = t_r43_c49_11 + p_44_50;
  assign out_43_49 = t_r43_c49_12 >> 4;

  assign t_r43_c50_0 = p_42_50 << 1;
  assign t_r43_c50_1 = p_43_49 << 1;
  assign t_r43_c50_2 = p_43_50 << 2;
  assign t_r43_c50_3 = p_43_51 << 1;
  assign t_r43_c50_4 = p_44_50 << 1;
  assign t_r43_c50_5 = t_r43_c50_0 + p_42_49;
  assign t_r43_c50_6 = t_r43_c50_1 + p_42_51;
  assign t_r43_c50_7 = t_r43_c50_2 + t_r43_c50_3;
  assign t_r43_c50_8 = t_r43_c50_4 + p_44_49;
  assign t_r43_c50_9 = t_r43_c50_5 + t_r43_c50_6;
  assign t_r43_c50_10 = t_r43_c50_7 + t_r43_c50_8;
  assign t_r43_c50_11 = t_r43_c50_9 + t_r43_c50_10;
  assign t_r43_c50_12 = t_r43_c50_11 + p_44_51;
  assign out_43_50 = t_r43_c50_12 >> 4;

  assign t_r43_c51_0 = p_42_51 << 1;
  assign t_r43_c51_1 = p_43_50 << 1;
  assign t_r43_c51_2 = p_43_51 << 2;
  assign t_r43_c51_3 = p_43_52 << 1;
  assign t_r43_c51_4 = p_44_51 << 1;
  assign t_r43_c51_5 = t_r43_c51_0 + p_42_50;
  assign t_r43_c51_6 = t_r43_c51_1 + p_42_52;
  assign t_r43_c51_7 = t_r43_c51_2 + t_r43_c51_3;
  assign t_r43_c51_8 = t_r43_c51_4 + p_44_50;
  assign t_r43_c51_9 = t_r43_c51_5 + t_r43_c51_6;
  assign t_r43_c51_10 = t_r43_c51_7 + t_r43_c51_8;
  assign t_r43_c51_11 = t_r43_c51_9 + t_r43_c51_10;
  assign t_r43_c51_12 = t_r43_c51_11 + p_44_52;
  assign out_43_51 = t_r43_c51_12 >> 4;

  assign t_r43_c52_0 = p_42_52 << 1;
  assign t_r43_c52_1 = p_43_51 << 1;
  assign t_r43_c52_2 = p_43_52 << 2;
  assign t_r43_c52_3 = p_43_53 << 1;
  assign t_r43_c52_4 = p_44_52 << 1;
  assign t_r43_c52_5 = t_r43_c52_0 + p_42_51;
  assign t_r43_c52_6 = t_r43_c52_1 + p_42_53;
  assign t_r43_c52_7 = t_r43_c52_2 + t_r43_c52_3;
  assign t_r43_c52_8 = t_r43_c52_4 + p_44_51;
  assign t_r43_c52_9 = t_r43_c52_5 + t_r43_c52_6;
  assign t_r43_c52_10 = t_r43_c52_7 + t_r43_c52_8;
  assign t_r43_c52_11 = t_r43_c52_9 + t_r43_c52_10;
  assign t_r43_c52_12 = t_r43_c52_11 + p_44_53;
  assign out_43_52 = t_r43_c52_12 >> 4;

  assign t_r43_c53_0 = p_42_53 << 1;
  assign t_r43_c53_1 = p_43_52 << 1;
  assign t_r43_c53_2 = p_43_53 << 2;
  assign t_r43_c53_3 = p_43_54 << 1;
  assign t_r43_c53_4 = p_44_53 << 1;
  assign t_r43_c53_5 = t_r43_c53_0 + p_42_52;
  assign t_r43_c53_6 = t_r43_c53_1 + p_42_54;
  assign t_r43_c53_7 = t_r43_c53_2 + t_r43_c53_3;
  assign t_r43_c53_8 = t_r43_c53_4 + p_44_52;
  assign t_r43_c53_9 = t_r43_c53_5 + t_r43_c53_6;
  assign t_r43_c53_10 = t_r43_c53_7 + t_r43_c53_8;
  assign t_r43_c53_11 = t_r43_c53_9 + t_r43_c53_10;
  assign t_r43_c53_12 = t_r43_c53_11 + p_44_54;
  assign out_43_53 = t_r43_c53_12 >> 4;

  assign t_r43_c54_0 = p_42_54 << 1;
  assign t_r43_c54_1 = p_43_53 << 1;
  assign t_r43_c54_2 = p_43_54 << 2;
  assign t_r43_c54_3 = p_43_55 << 1;
  assign t_r43_c54_4 = p_44_54 << 1;
  assign t_r43_c54_5 = t_r43_c54_0 + p_42_53;
  assign t_r43_c54_6 = t_r43_c54_1 + p_42_55;
  assign t_r43_c54_7 = t_r43_c54_2 + t_r43_c54_3;
  assign t_r43_c54_8 = t_r43_c54_4 + p_44_53;
  assign t_r43_c54_9 = t_r43_c54_5 + t_r43_c54_6;
  assign t_r43_c54_10 = t_r43_c54_7 + t_r43_c54_8;
  assign t_r43_c54_11 = t_r43_c54_9 + t_r43_c54_10;
  assign t_r43_c54_12 = t_r43_c54_11 + p_44_55;
  assign out_43_54 = t_r43_c54_12 >> 4;

  assign t_r43_c55_0 = p_42_55 << 1;
  assign t_r43_c55_1 = p_43_54 << 1;
  assign t_r43_c55_2 = p_43_55 << 2;
  assign t_r43_c55_3 = p_43_56 << 1;
  assign t_r43_c55_4 = p_44_55 << 1;
  assign t_r43_c55_5 = t_r43_c55_0 + p_42_54;
  assign t_r43_c55_6 = t_r43_c55_1 + p_42_56;
  assign t_r43_c55_7 = t_r43_c55_2 + t_r43_c55_3;
  assign t_r43_c55_8 = t_r43_c55_4 + p_44_54;
  assign t_r43_c55_9 = t_r43_c55_5 + t_r43_c55_6;
  assign t_r43_c55_10 = t_r43_c55_7 + t_r43_c55_8;
  assign t_r43_c55_11 = t_r43_c55_9 + t_r43_c55_10;
  assign t_r43_c55_12 = t_r43_c55_11 + p_44_56;
  assign out_43_55 = t_r43_c55_12 >> 4;

  assign t_r43_c56_0 = p_42_56 << 1;
  assign t_r43_c56_1 = p_43_55 << 1;
  assign t_r43_c56_2 = p_43_56 << 2;
  assign t_r43_c56_3 = p_43_57 << 1;
  assign t_r43_c56_4 = p_44_56 << 1;
  assign t_r43_c56_5 = t_r43_c56_0 + p_42_55;
  assign t_r43_c56_6 = t_r43_c56_1 + p_42_57;
  assign t_r43_c56_7 = t_r43_c56_2 + t_r43_c56_3;
  assign t_r43_c56_8 = t_r43_c56_4 + p_44_55;
  assign t_r43_c56_9 = t_r43_c56_5 + t_r43_c56_6;
  assign t_r43_c56_10 = t_r43_c56_7 + t_r43_c56_8;
  assign t_r43_c56_11 = t_r43_c56_9 + t_r43_c56_10;
  assign t_r43_c56_12 = t_r43_c56_11 + p_44_57;
  assign out_43_56 = t_r43_c56_12 >> 4;

  assign t_r43_c57_0 = p_42_57 << 1;
  assign t_r43_c57_1 = p_43_56 << 1;
  assign t_r43_c57_2 = p_43_57 << 2;
  assign t_r43_c57_3 = p_43_58 << 1;
  assign t_r43_c57_4 = p_44_57 << 1;
  assign t_r43_c57_5 = t_r43_c57_0 + p_42_56;
  assign t_r43_c57_6 = t_r43_c57_1 + p_42_58;
  assign t_r43_c57_7 = t_r43_c57_2 + t_r43_c57_3;
  assign t_r43_c57_8 = t_r43_c57_4 + p_44_56;
  assign t_r43_c57_9 = t_r43_c57_5 + t_r43_c57_6;
  assign t_r43_c57_10 = t_r43_c57_7 + t_r43_c57_8;
  assign t_r43_c57_11 = t_r43_c57_9 + t_r43_c57_10;
  assign t_r43_c57_12 = t_r43_c57_11 + p_44_58;
  assign out_43_57 = t_r43_c57_12 >> 4;

  assign t_r43_c58_0 = p_42_58 << 1;
  assign t_r43_c58_1 = p_43_57 << 1;
  assign t_r43_c58_2 = p_43_58 << 2;
  assign t_r43_c58_3 = p_43_59 << 1;
  assign t_r43_c58_4 = p_44_58 << 1;
  assign t_r43_c58_5 = t_r43_c58_0 + p_42_57;
  assign t_r43_c58_6 = t_r43_c58_1 + p_42_59;
  assign t_r43_c58_7 = t_r43_c58_2 + t_r43_c58_3;
  assign t_r43_c58_8 = t_r43_c58_4 + p_44_57;
  assign t_r43_c58_9 = t_r43_c58_5 + t_r43_c58_6;
  assign t_r43_c58_10 = t_r43_c58_7 + t_r43_c58_8;
  assign t_r43_c58_11 = t_r43_c58_9 + t_r43_c58_10;
  assign t_r43_c58_12 = t_r43_c58_11 + p_44_59;
  assign out_43_58 = t_r43_c58_12 >> 4;

  assign t_r43_c59_0 = p_42_59 << 1;
  assign t_r43_c59_1 = p_43_58 << 1;
  assign t_r43_c59_2 = p_43_59 << 2;
  assign t_r43_c59_3 = p_43_60 << 1;
  assign t_r43_c59_4 = p_44_59 << 1;
  assign t_r43_c59_5 = t_r43_c59_0 + p_42_58;
  assign t_r43_c59_6 = t_r43_c59_1 + p_42_60;
  assign t_r43_c59_7 = t_r43_c59_2 + t_r43_c59_3;
  assign t_r43_c59_8 = t_r43_c59_4 + p_44_58;
  assign t_r43_c59_9 = t_r43_c59_5 + t_r43_c59_6;
  assign t_r43_c59_10 = t_r43_c59_7 + t_r43_c59_8;
  assign t_r43_c59_11 = t_r43_c59_9 + t_r43_c59_10;
  assign t_r43_c59_12 = t_r43_c59_11 + p_44_60;
  assign out_43_59 = t_r43_c59_12 >> 4;

  assign t_r43_c60_0 = p_42_60 << 1;
  assign t_r43_c60_1 = p_43_59 << 1;
  assign t_r43_c60_2 = p_43_60 << 2;
  assign t_r43_c60_3 = p_43_61 << 1;
  assign t_r43_c60_4 = p_44_60 << 1;
  assign t_r43_c60_5 = t_r43_c60_0 + p_42_59;
  assign t_r43_c60_6 = t_r43_c60_1 + p_42_61;
  assign t_r43_c60_7 = t_r43_c60_2 + t_r43_c60_3;
  assign t_r43_c60_8 = t_r43_c60_4 + p_44_59;
  assign t_r43_c60_9 = t_r43_c60_5 + t_r43_c60_6;
  assign t_r43_c60_10 = t_r43_c60_7 + t_r43_c60_8;
  assign t_r43_c60_11 = t_r43_c60_9 + t_r43_c60_10;
  assign t_r43_c60_12 = t_r43_c60_11 + p_44_61;
  assign out_43_60 = t_r43_c60_12 >> 4;

  assign t_r43_c61_0 = p_42_61 << 1;
  assign t_r43_c61_1 = p_43_60 << 1;
  assign t_r43_c61_2 = p_43_61 << 2;
  assign t_r43_c61_3 = p_43_62 << 1;
  assign t_r43_c61_4 = p_44_61 << 1;
  assign t_r43_c61_5 = t_r43_c61_0 + p_42_60;
  assign t_r43_c61_6 = t_r43_c61_1 + p_42_62;
  assign t_r43_c61_7 = t_r43_c61_2 + t_r43_c61_3;
  assign t_r43_c61_8 = t_r43_c61_4 + p_44_60;
  assign t_r43_c61_9 = t_r43_c61_5 + t_r43_c61_6;
  assign t_r43_c61_10 = t_r43_c61_7 + t_r43_c61_8;
  assign t_r43_c61_11 = t_r43_c61_9 + t_r43_c61_10;
  assign t_r43_c61_12 = t_r43_c61_11 + p_44_62;
  assign out_43_61 = t_r43_c61_12 >> 4;

  assign t_r43_c62_0 = p_42_62 << 1;
  assign t_r43_c62_1 = p_43_61 << 1;
  assign t_r43_c62_2 = p_43_62 << 2;
  assign t_r43_c62_3 = p_43_63 << 1;
  assign t_r43_c62_4 = p_44_62 << 1;
  assign t_r43_c62_5 = t_r43_c62_0 + p_42_61;
  assign t_r43_c62_6 = t_r43_c62_1 + p_42_63;
  assign t_r43_c62_7 = t_r43_c62_2 + t_r43_c62_3;
  assign t_r43_c62_8 = t_r43_c62_4 + p_44_61;
  assign t_r43_c62_9 = t_r43_c62_5 + t_r43_c62_6;
  assign t_r43_c62_10 = t_r43_c62_7 + t_r43_c62_8;
  assign t_r43_c62_11 = t_r43_c62_9 + t_r43_c62_10;
  assign t_r43_c62_12 = t_r43_c62_11 + p_44_63;
  assign out_43_62 = t_r43_c62_12 >> 4;

  assign t_r43_c63_0 = p_42_63 << 1;
  assign t_r43_c63_1 = p_43_62 << 1;
  assign t_r43_c63_2 = p_43_63 << 2;
  assign t_r43_c63_3 = p_43_64 << 1;
  assign t_r43_c63_4 = p_44_63 << 1;
  assign t_r43_c63_5 = t_r43_c63_0 + p_42_62;
  assign t_r43_c63_6 = t_r43_c63_1 + p_42_64;
  assign t_r43_c63_7 = t_r43_c63_2 + t_r43_c63_3;
  assign t_r43_c63_8 = t_r43_c63_4 + p_44_62;
  assign t_r43_c63_9 = t_r43_c63_5 + t_r43_c63_6;
  assign t_r43_c63_10 = t_r43_c63_7 + t_r43_c63_8;
  assign t_r43_c63_11 = t_r43_c63_9 + t_r43_c63_10;
  assign t_r43_c63_12 = t_r43_c63_11 + p_44_64;
  assign out_43_63 = t_r43_c63_12 >> 4;

  assign t_r43_c64_0 = p_42_64 << 1;
  assign t_r43_c64_1 = p_43_63 << 1;
  assign t_r43_c64_2 = p_43_64 << 2;
  assign t_r43_c64_3 = p_43_65 << 1;
  assign t_r43_c64_4 = p_44_64 << 1;
  assign t_r43_c64_5 = t_r43_c64_0 + p_42_63;
  assign t_r43_c64_6 = t_r43_c64_1 + p_42_65;
  assign t_r43_c64_7 = t_r43_c64_2 + t_r43_c64_3;
  assign t_r43_c64_8 = t_r43_c64_4 + p_44_63;
  assign t_r43_c64_9 = t_r43_c64_5 + t_r43_c64_6;
  assign t_r43_c64_10 = t_r43_c64_7 + t_r43_c64_8;
  assign t_r43_c64_11 = t_r43_c64_9 + t_r43_c64_10;
  assign t_r43_c64_12 = t_r43_c64_11 + p_44_65;
  assign out_43_64 = t_r43_c64_12 >> 4;

endmodule
