module adder(G11,G12,G14);
input [1:0] G11,G12;
output [1:0] G14;
assign G14 = G11+G12;
endmodule
