module adder(G11, G12, G14);
  wire _00_, _01_, _02_, _03_, _04_, _05_, _06_, _07_, _08_, _09_, _10_, _11_, _12_, _13_, _14_, _15_, _16_, _17_, _18_, _19_, _20_, _21_, _22_, _23_, _24_, _25_;
  input [7:0] G11;
  input [7:0] G12;
  input G11[0], G11[1], G11[2], G11[3], G11[4], G11[5], G11[6], G11[7], G12[0], G12[1], G12[2], G12[3], G12[4], G12[5], G12[6], G12[7];
  output G14[0], G14[1], G14[2], G14[3], G14[4], G14[5], G14[6], G14[7];
  lut lut_gate1(0x6, _01_, _00_, G14[1]);
  lut lut_gate2(0x8, G11[0], G12[0], _00_);
  lut lut_gate3(0x6, G11[1], G12[1], _01_);
  lut lut_gate4(0x9, _05_, _02_, G14[2]);
  lut lut_gate5(0x1, _04_, _03_, _02_);
  lut lut_gate6(0x8, _01_, _00_, _03_);
  lut lut_gate7(0x8, G11[1], G12[1], _04_);
  lut lut_gate8(0x6, G11[2], G12[2], _05_);
  lut lut_gate9(0x9, _09_, _06_, G14[3]);
  lut lut_gate10(0x1, _08_, _07_, _06_);
  lut lut_gate11(0x4, _05_, _02_, _07_);
  lut lut_gate12(0x8, G11[2], G12[2], _08_);
  lut lut_gate13(0x6, G11[3], G12[3], _09_);
  lut lut_gate14(0x9, _13_, _10_, G14[4]);
  lut lut_gate15(0x1, _12_, _11_, _10_);
  lut lut_gate16(0x4, _09_, _06_, _11_);
  lut lut_gate17(0x8, G11[3], G12[3], _12_);
  lut lut_gate18(0x6, G11[4], G12[4], _13_);
  lut lut_gate19(0x6, G11[0], G12[0], G14[0]);
  lut lut_gate20(0x6, _25_, _14_, G14[7]);
  lut lut_gate21(0x1, _24_, _15_, _14_);
  lut lut_gate22(0x4, _23_, _16_, _15_);
  lut lut_gate23(0x1, _22_, _17_, _16_);
  lut lut_gate24(0x4, _21_, _18_, _17_);
  lut lut_gate25(0x1, _20_, _19_, _18_);
  lut lut_gate26(0x4, _13_, _10_, _19_);
  lut lut_gate27(0x8, G11[4], G12[4], _20_);
  lut lut_gate28(0x6, G11[5], G12[5], _21_);
  lut lut_gate29(0x8, G11[5], G12[5], _22_);
  lut lut_gate30(0x6, G11[6], G12[6], _23_);
  lut lut_gate31(0x8, G11[6], G12[6], _24_);
  lut lut_gate32(0x9, G11[7], G12[7], _25_);
  lut lut_gate33(0x9, _21_, _18_, G14[5]);
  lut lut_gate34(0x9, _23_, _16_, G14[6]);

endmodule
