module mmult (a_0_0, b_0_0, a_0_1, b_0_1, a_0_2, b_0_2, a_0_3, b_0_3, a_0_4, b_0_4, a_1_0, b_1_0, a_1_1, b_1_1, a_1_2, b_1_2, a_1_3, b_1_3, a_1_4, b_1_4, a_2_0, b_2_0, a_2_1, b_2_1, a_2_2, b_2_2, a_2_3, b_2_3, a_2_4, b_2_4, a_3_0, b_3_0, a_3_1, b_3_1, a_3_2, b_3_2, a_3_3, b_3_3, a_3_4, b_3_4, a_4_0, b_4_0, a_4_1, b_4_1, a_4_2, b_4_2, a_4_3, b_4_3, a_4_4, b_4_4, c_0_0, c_0_1, c_0_2, c_0_3, c_0_4, c_1_0, c_1_1, c_1_2, c_1_3, c_1_4, c_2_0, c_2_1, c_2_2, c_2_3, c_2_4, c_3_0, c_3_1, c_3_2, c_3_3, c_3_4, c_4_0, c_4_1, c_4_2, c_4_3, c_4_4);

  input [15:0] a_0_0;
  input [15:0] b_0_0;
  input [15:0] a_0_1;
  input [15:0] b_0_1;
  input [15:0] a_0_2;
  input [15:0] b_0_2;
  input [15:0] a_0_3;
  input [15:0] b_0_3;
  input [15:0] a_0_4;
  input [15:0] b_0_4;
  input [15:0] a_1_0;
  input [15:0] b_1_0;
  input [15:0] a_1_1;
  input [15:0] b_1_1;
  input [15:0] a_1_2;
  input [15:0] b_1_2;
  input [15:0] a_1_3;
  input [15:0] b_1_3;
  input [15:0] a_1_4;
  input [15:0] b_1_4;
  input [15:0] a_2_0;
  input [15:0] b_2_0;
  input [15:0] a_2_1;
  input [15:0] b_2_1;
  input [15:0] a_2_2;
  input [15:0] b_2_2;
  input [15:0] a_2_3;
  input [15:0] b_2_3;
  input [15:0] a_2_4;
  input [15:0] b_2_4;
  input [15:0] a_3_0;
  input [15:0] b_3_0;
  input [15:0] a_3_1;
  input [15:0] b_3_1;
  input [15:0] a_3_2;
  input [15:0] b_3_2;
  input [15:0] a_3_3;
  input [15:0] b_3_3;
  input [15:0] a_3_4;
  input [15:0] b_3_4;
  input [15:0] a_4_0;
  input [15:0] b_4_0;
  input [15:0] a_4_1;
  input [15:0] b_4_1;
  input [15:0] a_4_2;
  input [15:0] b_4_2;
  input [15:0] a_4_3;
  input [15:0] b_4_3;
  input [15:0] a_4_4;
  input [15:0] b_4_4;

  output [15:0] c_0_0;
  output [15:0] c_0_1;
  output [15:0] c_0_2;
  output [15:0] c_0_3;
  output [15:0] c_0_4;
  output [15:0] c_1_0;
  output [15:0] c_1_1;
  output [15:0] c_1_2;
  output [15:0] c_1_3;
  output [15:0] c_1_4;
  output [15:0] c_2_0;
  output [15:0] c_2_1;
  output [15:0] c_2_2;
  output [15:0] c_2_3;
  output [15:0] c_2_4;
  output [15:0] c_3_0;
  output [15:0] c_3_1;
  output [15:0] c_3_2;
  output [15:0] c_3_3;
  output [15:0] c_3_4;
  output [15:0] c_4_0;
  output [15:0] c_4_1;
  output [15:0] c_4_2;
  output [15:0] c_4_3;
  output [15:0] c_4_4;

  wire [15:0] t0_r0_c0_rr0;
  wire [15:0] t0_r0_c0_rr1;
  wire [15:0] t0_r0_c0_rr2;
  wire [15:0] t0_r0_c0_rr3;
  wire [15:0] t0_r0_c0_rr4;
  wire [15:0] t1_r0_c0_rr0;
  wire [15:0] t1_r0_c0_rr1;
  wire [15:0] t1_r0_c0_rr2;
  wire [15:0] t2_r0_c0_rr0;
  wire [15:0] t2_r0_c0_rr1;
  wire [15:0] t3_r0_c0_rr0;
  wire [15:0] t0_r0_c1_rr0;
  wire [15:0] t0_r0_c1_rr1;
  wire [15:0] t0_r0_c1_rr2;
  wire [15:0] t0_r0_c1_rr3;
  wire [15:0] t0_r0_c1_rr4;
  wire [15:0] t1_r0_c1_rr0;
  wire [15:0] t1_r0_c1_rr1;
  wire [15:0] t1_r0_c1_rr2;
  wire [15:0] t2_r0_c1_rr0;
  wire [15:0] t2_r0_c1_rr1;
  wire [15:0] t3_r0_c1_rr0;
  wire [15:0] t0_r0_c2_rr0;
  wire [15:0] t0_r0_c2_rr1;
  wire [15:0] t0_r0_c2_rr2;
  wire [15:0] t0_r0_c2_rr3;
  wire [15:0] t0_r0_c2_rr4;
  wire [15:0] t1_r0_c2_rr0;
  wire [15:0] t1_r0_c2_rr1;
  wire [15:0] t1_r0_c2_rr2;
  wire [15:0] t2_r0_c2_rr0;
  wire [15:0] t2_r0_c2_rr1;
  wire [15:0] t3_r0_c2_rr0;
  wire [15:0] t0_r0_c3_rr0;
  wire [15:0] t0_r0_c3_rr1;
  wire [15:0] t0_r0_c3_rr2;
  wire [15:0] t0_r0_c3_rr3;
  wire [15:0] t0_r0_c3_rr4;
  wire [15:0] t1_r0_c3_rr0;
  wire [15:0] t1_r0_c3_rr1;
  wire [15:0] t1_r0_c3_rr2;
  wire [15:0] t2_r0_c3_rr0;
  wire [15:0] t2_r0_c3_rr1;
  wire [15:0] t3_r0_c3_rr0;
  wire [15:0] t0_r0_c4_rr0;
  wire [15:0] t0_r0_c4_rr1;
  wire [15:0] t0_r0_c4_rr2;
  wire [15:0] t0_r0_c4_rr3;
  wire [15:0] t0_r0_c4_rr4;
  wire [15:0] t1_r0_c4_rr0;
  wire [15:0] t1_r0_c4_rr1;
  wire [15:0] t1_r0_c4_rr2;
  wire [15:0] t2_r0_c4_rr0;
  wire [15:0] t2_r0_c4_rr1;
  wire [15:0] t3_r0_c4_rr0;
  wire [15:0] t0_r1_c0_rr0;
  wire [15:0] t0_r1_c0_rr1;
  wire [15:0] t0_r1_c0_rr2;
  wire [15:0] t0_r1_c0_rr3;
  wire [15:0] t0_r1_c0_rr4;
  wire [15:0] t1_r1_c0_rr0;
  wire [15:0] t1_r1_c0_rr1;
  wire [15:0] t1_r1_c0_rr2;
  wire [15:0] t2_r1_c0_rr0;
  wire [15:0] t2_r1_c0_rr1;
  wire [15:0] t3_r1_c0_rr0;
  wire [15:0] t0_r1_c1_rr0;
  wire [15:0] t0_r1_c1_rr1;
  wire [15:0] t0_r1_c1_rr2;
  wire [15:0] t0_r1_c1_rr3;
  wire [15:0] t0_r1_c1_rr4;
  wire [15:0] t1_r1_c1_rr0;
  wire [15:0] t1_r1_c1_rr1;
  wire [15:0] t1_r1_c1_rr2;
  wire [15:0] t2_r1_c1_rr0;
  wire [15:0] t2_r1_c1_rr1;
  wire [15:0] t3_r1_c1_rr0;
  wire [15:0] t0_r1_c2_rr0;
  wire [15:0] t0_r1_c2_rr1;
  wire [15:0] t0_r1_c2_rr2;
  wire [15:0] t0_r1_c2_rr3;
  wire [15:0] t0_r1_c2_rr4;
  wire [15:0] t1_r1_c2_rr0;
  wire [15:0] t1_r1_c2_rr1;
  wire [15:0] t1_r1_c2_rr2;
  wire [15:0] t2_r1_c2_rr0;
  wire [15:0] t2_r1_c2_rr1;
  wire [15:0] t3_r1_c2_rr0;
  wire [15:0] t0_r1_c3_rr0;
  wire [15:0] t0_r1_c3_rr1;
  wire [15:0] t0_r1_c3_rr2;
  wire [15:0] t0_r1_c3_rr3;
  wire [15:0] t0_r1_c3_rr4;
  wire [15:0] t1_r1_c3_rr0;
  wire [15:0] t1_r1_c3_rr1;
  wire [15:0] t1_r1_c3_rr2;
  wire [15:0] t2_r1_c3_rr0;
  wire [15:0] t2_r1_c3_rr1;
  wire [15:0] t3_r1_c3_rr0;
  wire [15:0] t0_r1_c4_rr0;
  wire [15:0] t0_r1_c4_rr1;
  wire [15:0] t0_r1_c4_rr2;
  wire [15:0] t0_r1_c4_rr3;
  wire [15:0] t0_r1_c4_rr4;
  wire [15:0] t1_r1_c4_rr0;
  wire [15:0] t1_r1_c4_rr1;
  wire [15:0] t1_r1_c4_rr2;
  wire [15:0] t2_r1_c4_rr0;
  wire [15:0] t2_r1_c4_rr1;
  wire [15:0] t3_r1_c4_rr0;
  wire [15:0] t0_r2_c0_rr0;
  wire [15:0] t0_r2_c0_rr1;
  wire [15:0] t0_r2_c0_rr2;
  wire [15:0] t0_r2_c0_rr3;
  wire [15:0] t0_r2_c0_rr4;
  wire [15:0] t1_r2_c0_rr0;
  wire [15:0] t1_r2_c0_rr1;
  wire [15:0] t1_r2_c0_rr2;
  wire [15:0] t2_r2_c0_rr0;
  wire [15:0] t2_r2_c0_rr1;
  wire [15:0] t3_r2_c0_rr0;
  wire [15:0] t0_r2_c1_rr0;
  wire [15:0] t0_r2_c1_rr1;
  wire [15:0] t0_r2_c1_rr2;
  wire [15:0] t0_r2_c1_rr3;
  wire [15:0] t0_r2_c1_rr4;
  wire [15:0] t1_r2_c1_rr0;
  wire [15:0] t1_r2_c1_rr1;
  wire [15:0] t1_r2_c1_rr2;
  wire [15:0] t2_r2_c1_rr0;
  wire [15:0] t2_r2_c1_rr1;
  wire [15:0] t3_r2_c1_rr0;
  wire [15:0] t0_r2_c2_rr0;
  wire [15:0] t0_r2_c2_rr1;
  wire [15:0] t0_r2_c2_rr2;
  wire [15:0] t0_r2_c2_rr3;
  wire [15:0] t0_r2_c2_rr4;
  wire [15:0] t1_r2_c2_rr0;
  wire [15:0] t1_r2_c2_rr1;
  wire [15:0] t1_r2_c2_rr2;
  wire [15:0] t2_r2_c2_rr0;
  wire [15:0] t2_r2_c2_rr1;
  wire [15:0] t3_r2_c2_rr0;
  wire [15:0] t0_r2_c3_rr0;
  wire [15:0] t0_r2_c3_rr1;
  wire [15:0] t0_r2_c3_rr2;
  wire [15:0] t0_r2_c3_rr3;
  wire [15:0] t0_r2_c3_rr4;
  wire [15:0] t1_r2_c3_rr0;
  wire [15:0] t1_r2_c3_rr1;
  wire [15:0] t1_r2_c3_rr2;
  wire [15:0] t2_r2_c3_rr0;
  wire [15:0] t2_r2_c3_rr1;
  wire [15:0] t3_r2_c3_rr0;
  wire [15:0] t0_r2_c4_rr0;
  wire [15:0] t0_r2_c4_rr1;
  wire [15:0] t0_r2_c4_rr2;
  wire [15:0] t0_r2_c4_rr3;
  wire [15:0] t0_r2_c4_rr4;
  wire [15:0] t1_r2_c4_rr0;
  wire [15:0] t1_r2_c4_rr1;
  wire [15:0] t1_r2_c4_rr2;
  wire [15:0] t2_r2_c4_rr0;
  wire [15:0] t2_r2_c4_rr1;
  wire [15:0] t3_r2_c4_rr0;
  wire [15:0] t0_r3_c0_rr0;
  wire [15:0] t0_r3_c0_rr1;
  wire [15:0] t0_r3_c0_rr2;
  wire [15:0] t0_r3_c0_rr3;
  wire [15:0] t0_r3_c0_rr4;
  wire [15:0] t1_r3_c0_rr0;
  wire [15:0] t1_r3_c0_rr1;
  wire [15:0] t1_r3_c0_rr2;
  wire [15:0] t2_r3_c0_rr0;
  wire [15:0] t2_r3_c0_rr1;
  wire [15:0] t3_r3_c0_rr0;
  wire [15:0] t0_r3_c1_rr0;
  wire [15:0] t0_r3_c1_rr1;
  wire [15:0] t0_r3_c1_rr2;
  wire [15:0] t0_r3_c1_rr3;
  wire [15:0] t0_r3_c1_rr4;
  wire [15:0] t1_r3_c1_rr0;
  wire [15:0] t1_r3_c1_rr1;
  wire [15:0] t1_r3_c1_rr2;
  wire [15:0] t2_r3_c1_rr0;
  wire [15:0] t2_r3_c1_rr1;
  wire [15:0] t3_r3_c1_rr0;
  wire [15:0] t0_r3_c2_rr0;
  wire [15:0] t0_r3_c2_rr1;
  wire [15:0] t0_r3_c2_rr2;
  wire [15:0] t0_r3_c2_rr3;
  wire [15:0] t0_r3_c2_rr4;
  wire [15:0] t1_r3_c2_rr0;
  wire [15:0] t1_r3_c2_rr1;
  wire [15:0] t1_r3_c2_rr2;
  wire [15:0] t2_r3_c2_rr0;
  wire [15:0] t2_r3_c2_rr1;
  wire [15:0] t3_r3_c2_rr0;
  wire [15:0] t0_r3_c3_rr0;
  wire [15:0] t0_r3_c3_rr1;
  wire [15:0] t0_r3_c3_rr2;
  wire [15:0] t0_r3_c3_rr3;
  wire [15:0] t0_r3_c3_rr4;
  wire [15:0] t1_r3_c3_rr0;
  wire [15:0] t1_r3_c3_rr1;
  wire [15:0] t1_r3_c3_rr2;
  wire [15:0] t2_r3_c3_rr0;
  wire [15:0] t2_r3_c3_rr1;
  wire [15:0] t3_r3_c3_rr0;
  wire [15:0] t0_r3_c4_rr0;
  wire [15:0] t0_r3_c4_rr1;
  wire [15:0] t0_r3_c4_rr2;
  wire [15:0] t0_r3_c4_rr3;
  wire [15:0] t0_r3_c4_rr4;
  wire [15:0] t1_r3_c4_rr0;
  wire [15:0] t1_r3_c4_rr1;
  wire [15:0] t1_r3_c4_rr2;
  wire [15:0] t2_r3_c4_rr0;
  wire [15:0] t2_r3_c4_rr1;
  wire [15:0] t3_r3_c4_rr0;
  wire [15:0] t0_r4_c0_rr0;
  wire [15:0] t0_r4_c0_rr1;
  wire [15:0] t0_r4_c0_rr2;
  wire [15:0] t0_r4_c0_rr3;
  wire [15:0] t0_r4_c0_rr4;
  wire [15:0] t1_r4_c0_rr0;
  wire [15:0] t1_r4_c0_rr1;
  wire [15:0] t1_r4_c0_rr2;
  wire [15:0] t2_r4_c0_rr0;
  wire [15:0] t2_r4_c0_rr1;
  wire [15:0] t3_r4_c0_rr0;
  wire [15:0] t0_r4_c1_rr0;
  wire [15:0] t0_r4_c1_rr1;
  wire [15:0] t0_r4_c1_rr2;
  wire [15:0] t0_r4_c1_rr3;
  wire [15:0] t0_r4_c1_rr4;
  wire [15:0] t1_r4_c1_rr0;
  wire [15:0] t1_r4_c1_rr1;
  wire [15:0] t1_r4_c1_rr2;
  wire [15:0] t2_r4_c1_rr0;
  wire [15:0] t2_r4_c1_rr1;
  wire [15:0] t3_r4_c1_rr0;
  wire [15:0] t0_r4_c2_rr0;
  wire [15:0] t0_r4_c2_rr1;
  wire [15:0] t0_r4_c2_rr2;
  wire [15:0] t0_r4_c2_rr3;
  wire [15:0] t0_r4_c2_rr4;
  wire [15:0] t1_r4_c2_rr0;
  wire [15:0] t1_r4_c2_rr1;
  wire [15:0] t1_r4_c2_rr2;
  wire [15:0] t2_r4_c2_rr0;
  wire [15:0] t2_r4_c2_rr1;
  wire [15:0] t3_r4_c2_rr0;
  wire [15:0] t0_r4_c3_rr0;
  wire [15:0] t0_r4_c3_rr1;
  wire [15:0] t0_r4_c3_rr2;
  wire [15:0] t0_r4_c3_rr3;
  wire [15:0] t0_r4_c3_rr4;
  wire [15:0] t1_r4_c3_rr0;
  wire [15:0] t1_r4_c3_rr1;
  wire [15:0] t1_r4_c3_rr2;
  wire [15:0] t2_r4_c3_rr0;
  wire [15:0] t2_r4_c3_rr1;
  wire [15:0] t3_r4_c3_rr0;
  wire [15:0] t0_r4_c4_rr0;
  wire [15:0] t0_r4_c4_rr1;
  wire [15:0] t0_r4_c4_rr2;
  wire [15:0] t0_r4_c4_rr3;
  wire [15:0] t0_r4_c4_rr4;
  wire [15:0] t1_r4_c4_rr0;
  wire [15:0] t1_r4_c4_rr1;
  wire [15:0] t1_r4_c4_rr2;
  wire [15:0] t2_r4_c4_rr0;
  wire [15:0] t2_r4_c4_rr1;
  wire [15:0] t3_r4_c4_rr0;

  assign t0_r0_c0_rr0 = a_0_0 * b_0_0;
  assign t0_r0_c0_rr1 = a_0_1 * b_1_0;
  assign t0_r0_c0_rr2 = a_0_2 * b_2_0;
  assign t0_r0_c0_rr3 = a_0_3 * b_3_0;
  assign t0_r0_c0_rr4 = a_0_4 * b_4_0;
  assign t1_r0_c0_rr0 = t0_r0_c0_rr0 + t0_r0_c0_rr1;
  assign t1_r0_c0_rr1 = t0_r0_c0_rr2 + t0_r0_c0_rr3;
  assign t1_r0_c0_rr2 = t0_r0_c0_rr4;

  assign t2_r0_c0_rr0 = t1_r0_c0_rr0 + t1_r0_c0_rr1;
  assign t2_r0_c0_rr1 = t1_r0_c0_rr2;

  assign t3_r0_c0_rr0 = t2_r0_c0_rr0 + t2_r0_c0_rr1;

  assign c_0_0 = t3_r0_c0_rr0;
  assign t0_r0_c1_rr0 = a_0_0 * b_0_1;
  assign t0_r0_c1_rr1 = a_0_1 * b_1_1;
  assign t0_r0_c1_rr2 = a_0_2 * b_2_1;
  assign t0_r0_c1_rr3 = a_0_3 * b_3_1;
  assign t0_r0_c1_rr4 = a_0_4 * b_4_1;
  assign t1_r0_c1_rr0 = t0_r0_c1_rr0 + t0_r0_c1_rr1;
  assign t1_r0_c1_rr1 = t0_r0_c1_rr2 + t0_r0_c1_rr3;
  assign t1_r0_c1_rr2 = t0_r0_c1_rr4;

  assign t2_r0_c1_rr0 = t1_r0_c1_rr0 + t1_r0_c1_rr1;
  assign t2_r0_c1_rr1 = t1_r0_c1_rr2;

  assign t3_r0_c1_rr0 = t2_r0_c1_rr0 + t2_r0_c1_rr1;

  assign c_0_1 = t3_r0_c1_rr0;
  assign t0_r0_c2_rr0 = a_0_0 * b_0_2;
  assign t0_r0_c2_rr1 = a_0_1 * b_1_2;
  assign t0_r0_c2_rr2 = a_0_2 * b_2_2;
  assign t0_r0_c2_rr3 = a_0_3 * b_3_2;
  assign t0_r0_c2_rr4 = a_0_4 * b_4_2;
  assign t1_r0_c2_rr0 = t0_r0_c2_rr0 + t0_r0_c2_rr1;
  assign t1_r0_c2_rr1 = t0_r0_c2_rr2 + t0_r0_c2_rr3;
  assign t1_r0_c2_rr2 = t0_r0_c2_rr4;

  assign t2_r0_c2_rr0 = t1_r0_c2_rr0 + t1_r0_c2_rr1;
  assign t2_r0_c2_rr1 = t1_r0_c2_rr2;

  assign t3_r0_c2_rr0 = t2_r0_c2_rr0 + t2_r0_c2_rr1;

  assign c_0_2 = t3_r0_c2_rr0;
  assign t0_r0_c3_rr0 = a_0_0 * b_0_3;
  assign t0_r0_c3_rr1 = a_0_1 * b_1_3;
  assign t0_r0_c3_rr2 = a_0_2 * b_2_3;
  assign t0_r0_c3_rr3 = a_0_3 * b_3_3;
  assign t0_r0_c3_rr4 = a_0_4 * b_4_3;
  assign t1_r0_c3_rr0 = t0_r0_c3_rr0 + t0_r0_c3_rr1;
  assign t1_r0_c3_rr1 = t0_r0_c3_rr2 + t0_r0_c3_rr3;
  assign t1_r0_c3_rr2 = t0_r0_c3_rr4;

  assign t2_r0_c3_rr0 = t1_r0_c3_rr0 + t1_r0_c3_rr1;
  assign t2_r0_c3_rr1 = t1_r0_c3_rr2;

  assign t3_r0_c3_rr0 = t2_r0_c3_rr0 + t2_r0_c3_rr1;

  assign c_0_3 = t3_r0_c3_rr0;
  assign t0_r0_c4_rr0 = a_0_0 * b_0_4;
  assign t0_r0_c4_rr1 = a_0_1 * b_1_4;
  assign t0_r0_c4_rr2 = a_0_2 * b_2_4;
  assign t0_r0_c4_rr3 = a_0_3 * b_3_4;
  assign t0_r0_c4_rr4 = a_0_4 * b_4_4;
  assign t1_r0_c4_rr0 = t0_r0_c4_rr0 + t0_r0_c4_rr1;
  assign t1_r0_c4_rr1 = t0_r0_c4_rr2 + t0_r0_c4_rr3;
  assign t1_r0_c4_rr2 = t0_r0_c4_rr4;

  assign t2_r0_c4_rr0 = t1_r0_c4_rr0 + t1_r0_c4_rr1;
  assign t2_r0_c4_rr1 = t1_r0_c4_rr2;

  assign t3_r0_c4_rr0 = t2_r0_c4_rr0 + t2_r0_c4_rr1;

  assign c_0_4 = t3_r0_c4_rr0;
  assign t0_r1_c0_rr0 = a_1_0 * b_0_0;
  assign t0_r1_c0_rr1 = a_1_1 * b_1_0;
  assign t0_r1_c0_rr2 = a_1_2 * b_2_0;
  assign t0_r1_c0_rr3 = a_1_3 * b_3_0;
  assign t0_r1_c0_rr4 = a_1_4 * b_4_0;
  assign t1_r1_c0_rr0 = t0_r1_c0_rr0 + t0_r1_c0_rr1;
  assign t1_r1_c0_rr1 = t0_r1_c0_rr2 + t0_r1_c0_rr3;
  assign t1_r1_c0_rr2 = t0_r1_c0_rr4;

  assign t2_r1_c0_rr0 = t1_r1_c0_rr0 + t1_r1_c0_rr1;
  assign t2_r1_c0_rr1 = t1_r1_c0_rr2;

  assign t3_r1_c0_rr0 = t2_r1_c0_rr0 + t2_r1_c0_rr1;

  assign c_1_0 = t3_r1_c0_rr0;
  assign t0_r1_c1_rr0 = a_1_0 * b_0_1;
  assign t0_r1_c1_rr1 = a_1_1 * b_1_1;
  assign t0_r1_c1_rr2 = a_1_2 * b_2_1;
  assign t0_r1_c1_rr3 = a_1_3 * b_3_1;
  assign t0_r1_c1_rr4 = a_1_4 * b_4_1;
  assign t1_r1_c1_rr0 = t0_r1_c1_rr0 + t0_r1_c1_rr1;
  assign t1_r1_c1_rr1 = t0_r1_c1_rr2 + t0_r1_c1_rr3;
  assign t1_r1_c1_rr2 = t0_r1_c1_rr4;

  assign t2_r1_c1_rr0 = t1_r1_c1_rr0 + t1_r1_c1_rr1;
  assign t2_r1_c1_rr1 = t1_r1_c1_rr2;

  assign t3_r1_c1_rr0 = t2_r1_c1_rr0 + t2_r1_c1_rr1;

  assign c_1_1 = t3_r1_c1_rr0;
  assign t0_r1_c2_rr0 = a_1_0 * b_0_2;
  assign t0_r1_c2_rr1 = a_1_1 * b_1_2;
  assign t0_r1_c2_rr2 = a_1_2 * b_2_2;
  assign t0_r1_c2_rr3 = a_1_3 * b_3_2;
  assign t0_r1_c2_rr4 = a_1_4 * b_4_2;
  assign t1_r1_c2_rr0 = t0_r1_c2_rr0 + t0_r1_c2_rr1;
  assign t1_r1_c2_rr1 = t0_r1_c2_rr2 + t0_r1_c2_rr3;
  assign t1_r1_c2_rr2 = t0_r1_c2_rr4;

  assign t2_r1_c2_rr0 = t1_r1_c2_rr0 + t1_r1_c2_rr1;
  assign t2_r1_c2_rr1 = t1_r1_c2_rr2;

  assign t3_r1_c2_rr0 = t2_r1_c2_rr0 + t2_r1_c2_rr1;

  assign c_1_2 = t3_r1_c2_rr0;
  assign t0_r1_c3_rr0 = a_1_0 * b_0_3;
  assign t0_r1_c3_rr1 = a_1_1 * b_1_3;
  assign t0_r1_c3_rr2 = a_1_2 * b_2_3;
  assign t0_r1_c3_rr3 = a_1_3 * b_3_3;
  assign t0_r1_c3_rr4 = a_1_4 * b_4_3;
  assign t1_r1_c3_rr0 = t0_r1_c3_rr0 + t0_r1_c3_rr1;
  assign t1_r1_c3_rr1 = t0_r1_c3_rr2 + t0_r1_c3_rr3;
  assign t1_r1_c3_rr2 = t0_r1_c3_rr4;

  assign t2_r1_c3_rr0 = t1_r1_c3_rr0 + t1_r1_c3_rr1;
  assign t2_r1_c3_rr1 = t1_r1_c3_rr2;

  assign t3_r1_c3_rr0 = t2_r1_c3_rr0 + t2_r1_c3_rr1;

  assign c_1_3 = t3_r1_c3_rr0;
  assign t0_r1_c4_rr0 = a_1_0 * b_0_4;
  assign t0_r1_c4_rr1 = a_1_1 * b_1_4;
  assign t0_r1_c4_rr2 = a_1_2 * b_2_4;
  assign t0_r1_c4_rr3 = a_1_3 * b_3_4;
  assign t0_r1_c4_rr4 = a_1_4 * b_4_4;
  assign t1_r1_c4_rr0 = t0_r1_c4_rr0 + t0_r1_c4_rr1;
  assign t1_r1_c4_rr1 = t0_r1_c4_rr2 + t0_r1_c4_rr3;
  assign t1_r1_c4_rr2 = t0_r1_c4_rr4;

  assign t2_r1_c4_rr0 = t1_r1_c4_rr0 + t1_r1_c4_rr1;
  assign t2_r1_c4_rr1 = t1_r1_c4_rr2;

  assign t3_r1_c4_rr0 = t2_r1_c4_rr0 + t2_r1_c4_rr1;

  assign c_1_4 = t3_r1_c4_rr0;
  assign t0_r2_c0_rr0 = a_2_0 * b_0_0;
  assign t0_r2_c0_rr1 = a_2_1 * b_1_0;
  assign t0_r2_c0_rr2 = a_2_2 * b_2_0;
  assign t0_r2_c0_rr3 = a_2_3 * b_3_0;
  assign t0_r2_c0_rr4 = a_2_4 * b_4_0;
  assign t1_r2_c0_rr0 = t0_r2_c0_rr0 + t0_r2_c0_rr1;
  assign t1_r2_c0_rr1 = t0_r2_c0_rr2 + t0_r2_c0_rr3;
  assign t1_r2_c0_rr2 = t0_r2_c0_rr4;

  assign t2_r2_c0_rr0 = t1_r2_c0_rr0 + t1_r2_c0_rr1;
  assign t2_r2_c0_rr1 = t1_r2_c0_rr2;

  assign t3_r2_c0_rr0 = t2_r2_c0_rr0 + t2_r2_c0_rr1;

  assign c_2_0 = t3_r2_c0_rr0;
  assign t0_r2_c1_rr0 = a_2_0 * b_0_1;
  assign t0_r2_c1_rr1 = a_2_1 * b_1_1;
  assign t0_r2_c1_rr2 = a_2_2 * b_2_1;
  assign t0_r2_c1_rr3 = a_2_3 * b_3_1;
  assign t0_r2_c1_rr4 = a_2_4 * b_4_1;
  assign t1_r2_c1_rr0 = t0_r2_c1_rr0 + t0_r2_c1_rr1;
  assign t1_r2_c1_rr1 = t0_r2_c1_rr2 + t0_r2_c1_rr3;
  assign t1_r2_c1_rr2 = t0_r2_c1_rr4;

  assign t2_r2_c1_rr0 = t1_r2_c1_rr0 + t1_r2_c1_rr1;
  assign t2_r2_c1_rr1 = t1_r2_c1_rr2;

  assign t3_r2_c1_rr0 = t2_r2_c1_rr0 + t2_r2_c1_rr1;

  assign c_2_1 = t3_r2_c1_rr0;
  assign t0_r2_c2_rr0 = a_2_0 * b_0_2;
  assign t0_r2_c2_rr1 = a_2_1 * b_1_2;
  assign t0_r2_c2_rr2 = a_2_2 * b_2_2;
  assign t0_r2_c2_rr3 = a_2_3 * b_3_2;
  assign t0_r2_c2_rr4 = a_2_4 * b_4_2;
  assign t1_r2_c2_rr0 = t0_r2_c2_rr0 + t0_r2_c2_rr1;
  assign t1_r2_c2_rr1 = t0_r2_c2_rr2 + t0_r2_c2_rr3;
  assign t1_r2_c2_rr2 = t0_r2_c2_rr4;

  assign t2_r2_c2_rr0 = t1_r2_c2_rr0 + t1_r2_c2_rr1;
  assign t2_r2_c2_rr1 = t1_r2_c2_rr2;

  assign t3_r2_c2_rr0 = t2_r2_c2_rr0 + t2_r2_c2_rr1;

  assign c_2_2 = t3_r2_c2_rr0;
  assign t0_r2_c3_rr0 = a_2_0 * b_0_3;
  assign t0_r2_c3_rr1 = a_2_1 * b_1_3;
  assign t0_r2_c3_rr2 = a_2_2 * b_2_3;
  assign t0_r2_c3_rr3 = a_2_3 * b_3_3;
  assign t0_r2_c3_rr4 = a_2_4 * b_4_3;
  assign t1_r2_c3_rr0 = t0_r2_c3_rr0 + t0_r2_c3_rr1;
  assign t1_r2_c3_rr1 = t0_r2_c3_rr2 + t0_r2_c3_rr3;
  assign t1_r2_c3_rr2 = t0_r2_c3_rr4;

  assign t2_r2_c3_rr0 = t1_r2_c3_rr0 + t1_r2_c3_rr1;
  assign t2_r2_c3_rr1 = t1_r2_c3_rr2;

  assign t3_r2_c3_rr0 = t2_r2_c3_rr0 + t2_r2_c3_rr1;

  assign c_2_3 = t3_r2_c3_rr0;
  assign t0_r2_c4_rr0 = a_2_0 * b_0_4;
  assign t0_r2_c4_rr1 = a_2_1 * b_1_4;
  assign t0_r2_c4_rr2 = a_2_2 * b_2_4;
  assign t0_r2_c4_rr3 = a_2_3 * b_3_4;
  assign t0_r2_c4_rr4 = a_2_4 * b_4_4;
  assign t1_r2_c4_rr0 = t0_r2_c4_rr0 + t0_r2_c4_rr1;
  assign t1_r2_c4_rr1 = t0_r2_c4_rr2 + t0_r2_c4_rr3;
  assign t1_r2_c4_rr2 = t0_r2_c4_rr4;

  assign t2_r2_c4_rr0 = t1_r2_c4_rr0 + t1_r2_c4_rr1;
  assign t2_r2_c4_rr1 = t1_r2_c4_rr2;

  assign t3_r2_c4_rr0 = t2_r2_c4_rr0 + t2_r2_c4_rr1;

  assign c_2_4 = t3_r2_c4_rr0;
  assign t0_r3_c0_rr0 = a_3_0 * b_0_0;
  assign t0_r3_c0_rr1 = a_3_1 * b_1_0;
  assign t0_r3_c0_rr2 = a_3_2 * b_2_0;
  assign t0_r3_c0_rr3 = a_3_3 * b_3_0;
  assign t0_r3_c0_rr4 = a_3_4 * b_4_0;
  assign t1_r3_c0_rr0 = t0_r3_c0_rr0 + t0_r3_c0_rr1;
  assign t1_r3_c0_rr1 = t0_r3_c0_rr2 + t0_r3_c0_rr3;
  assign t1_r3_c0_rr2 = t0_r3_c0_rr4;

  assign t2_r3_c0_rr0 = t1_r3_c0_rr0 + t1_r3_c0_rr1;
  assign t2_r3_c0_rr1 = t1_r3_c0_rr2;

  assign t3_r3_c0_rr0 = t2_r3_c0_rr0 + t2_r3_c0_rr1;

  assign c_3_0 = t3_r3_c0_rr0;
  assign t0_r3_c1_rr0 = a_3_0 * b_0_1;
  assign t0_r3_c1_rr1 = a_3_1 * b_1_1;
  assign t0_r3_c1_rr2 = a_3_2 * b_2_1;
  assign t0_r3_c1_rr3 = a_3_3 * b_3_1;
  assign t0_r3_c1_rr4 = a_3_4 * b_4_1;
  assign t1_r3_c1_rr0 = t0_r3_c1_rr0 + t0_r3_c1_rr1;
  assign t1_r3_c1_rr1 = t0_r3_c1_rr2 + t0_r3_c1_rr3;
  assign t1_r3_c1_rr2 = t0_r3_c1_rr4;

  assign t2_r3_c1_rr0 = t1_r3_c1_rr0 + t1_r3_c1_rr1;
  assign t2_r3_c1_rr1 = t1_r3_c1_rr2;

  assign t3_r3_c1_rr0 = t2_r3_c1_rr0 + t2_r3_c1_rr1;

  assign c_3_1 = t3_r3_c1_rr0;
  assign t0_r3_c2_rr0 = a_3_0 * b_0_2;
  assign t0_r3_c2_rr1 = a_3_1 * b_1_2;
  assign t0_r3_c2_rr2 = a_3_2 * b_2_2;
  assign t0_r3_c2_rr3 = a_3_3 * b_3_2;
  assign t0_r3_c2_rr4 = a_3_4 * b_4_2;
  assign t1_r3_c2_rr0 = t0_r3_c2_rr0 + t0_r3_c2_rr1;
  assign t1_r3_c2_rr1 = t0_r3_c2_rr2 + t0_r3_c2_rr3;
  assign t1_r3_c2_rr2 = t0_r3_c2_rr4;

  assign t2_r3_c2_rr0 = t1_r3_c2_rr0 + t1_r3_c2_rr1;
  assign t2_r3_c2_rr1 = t1_r3_c2_rr2;

  assign t3_r3_c2_rr0 = t2_r3_c2_rr0 + t2_r3_c2_rr1;

  assign c_3_2 = t3_r3_c2_rr0;
  assign t0_r3_c3_rr0 = a_3_0 * b_0_3;
  assign t0_r3_c3_rr1 = a_3_1 * b_1_3;
  assign t0_r3_c3_rr2 = a_3_2 * b_2_3;
  assign t0_r3_c3_rr3 = a_3_3 * b_3_3;
  assign t0_r3_c3_rr4 = a_3_4 * b_4_3;
  assign t1_r3_c3_rr0 = t0_r3_c3_rr0 + t0_r3_c3_rr1;
  assign t1_r3_c3_rr1 = t0_r3_c3_rr2 + t0_r3_c3_rr3;
  assign t1_r3_c3_rr2 = t0_r3_c3_rr4;

  assign t2_r3_c3_rr0 = t1_r3_c3_rr0 + t1_r3_c3_rr1;
  assign t2_r3_c3_rr1 = t1_r3_c3_rr2;

  assign t3_r3_c3_rr0 = t2_r3_c3_rr0 + t2_r3_c3_rr1;

  assign c_3_3 = t3_r3_c3_rr0;
  assign t0_r3_c4_rr0 = a_3_0 * b_0_4;
  assign t0_r3_c4_rr1 = a_3_1 * b_1_4;
  assign t0_r3_c4_rr2 = a_3_2 * b_2_4;
  assign t0_r3_c4_rr3 = a_3_3 * b_3_4;
  assign t0_r3_c4_rr4 = a_3_4 * b_4_4;
  assign t1_r3_c4_rr0 = t0_r3_c4_rr0 + t0_r3_c4_rr1;
  assign t1_r3_c4_rr1 = t0_r3_c4_rr2 + t0_r3_c4_rr3;
  assign t1_r3_c4_rr2 = t0_r3_c4_rr4;

  assign t2_r3_c4_rr0 = t1_r3_c4_rr0 + t1_r3_c4_rr1;
  assign t2_r3_c4_rr1 = t1_r3_c4_rr2;

  assign t3_r3_c4_rr0 = t2_r3_c4_rr0 + t2_r3_c4_rr1;

  assign c_3_4 = t3_r3_c4_rr0;
  assign t0_r4_c0_rr0 = a_4_0 * b_0_0;
  assign t0_r4_c0_rr1 = a_4_1 * b_1_0;
  assign t0_r4_c0_rr2 = a_4_2 * b_2_0;
  assign t0_r4_c0_rr3 = a_4_3 * b_3_0;
  assign t0_r4_c0_rr4 = a_4_4 * b_4_0;
  assign t1_r4_c0_rr0 = t0_r4_c0_rr0 + t0_r4_c0_rr1;
  assign t1_r4_c0_rr1 = t0_r4_c0_rr2 + t0_r4_c0_rr3;
  assign t1_r4_c0_rr2 = t0_r4_c0_rr4;

  assign t2_r4_c0_rr0 = t1_r4_c0_rr0 + t1_r4_c0_rr1;
  assign t2_r4_c0_rr1 = t1_r4_c0_rr2;

  assign t3_r4_c0_rr0 = t2_r4_c0_rr0 + t2_r4_c0_rr1;

  assign c_4_0 = t3_r4_c0_rr0;
  assign t0_r4_c1_rr0 = a_4_0 * b_0_1;
  assign t0_r4_c1_rr1 = a_4_1 * b_1_1;
  assign t0_r4_c1_rr2 = a_4_2 * b_2_1;
  assign t0_r4_c1_rr3 = a_4_3 * b_3_1;
  assign t0_r4_c1_rr4 = a_4_4 * b_4_1;
  assign t1_r4_c1_rr0 = t0_r4_c1_rr0 + t0_r4_c1_rr1;
  assign t1_r4_c1_rr1 = t0_r4_c1_rr2 + t0_r4_c1_rr3;
  assign t1_r4_c1_rr2 = t0_r4_c1_rr4;

  assign t2_r4_c1_rr0 = t1_r4_c1_rr0 + t1_r4_c1_rr1;
  assign t2_r4_c1_rr1 = t1_r4_c1_rr2;

  assign t3_r4_c1_rr0 = t2_r4_c1_rr0 + t2_r4_c1_rr1;

  assign c_4_1 = t3_r4_c1_rr0;
  assign t0_r4_c2_rr0 = a_4_0 * b_0_2;
  assign t0_r4_c2_rr1 = a_4_1 * b_1_2;
  assign t0_r4_c2_rr2 = a_4_2 * b_2_2;
  assign t0_r4_c2_rr3 = a_4_3 * b_3_2;
  assign t0_r4_c2_rr4 = a_4_4 * b_4_2;
  assign t1_r4_c2_rr0 = t0_r4_c2_rr0 + t0_r4_c2_rr1;
  assign t1_r4_c2_rr1 = t0_r4_c2_rr2 + t0_r4_c2_rr3;
  assign t1_r4_c2_rr2 = t0_r4_c2_rr4;

  assign t2_r4_c2_rr0 = t1_r4_c2_rr0 + t1_r4_c2_rr1;
  assign t2_r4_c2_rr1 = t1_r4_c2_rr2;

  assign t3_r4_c2_rr0 = t2_r4_c2_rr0 + t2_r4_c2_rr1;

  assign c_4_2 = t3_r4_c2_rr0;
  assign t0_r4_c3_rr0 = a_4_0 * b_0_3;
  assign t0_r4_c3_rr1 = a_4_1 * b_1_3;
  assign t0_r4_c3_rr2 = a_4_2 * b_2_3;
  assign t0_r4_c3_rr3 = a_4_3 * b_3_3;
  assign t0_r4_c3_rr4 = a_4_4 * b_4_3;
  assign t1_r4_c3_rr0 = t0_r4_c3_rr0 + t0_r4_c3_rr1;
  assign t1_r4_c3_rr1 = t0_r4_c3_rr2 + t0_r4_c3_rr3;
  assign t1_r4_c3_rr2 = t0_r4_c3_rr4;

  assign t2_r4_c3_rr0 = t1_r4_c3_rr0 + t1_r4_c3_rr1;
  assign t2_r4_c3_rr1 = t1_r4_c3_rr2;

  assign t3_r4_c3_rr0 = t2_r4_c3_rr0 + t2_r4_c3_rr1;

  assign c_4_3 = t3_r4_c3_rr0;
  assign t0_r4_c4_rr0 = a_4_0 * b_0_4;
  assign t0_r4_c4_rr1 = a_4_1 * b_1_4;
  assign t0_r4_c4_rr2 = a_4_2 * b_2_4;
  assign t0_r4_c4_rr3 = a_4_3 * b_3_4;
  assign t0_r4_c4_rr4 = a_4_4 * b_4_4;
  assign t1_r4_c4_rr0 = t0_r4_c4_rr0 + t0_r4_c4_rr1;
  assign t1_r4_c4_rr1 = t0_r4_c4_rr2 + t0_r4_c4_rr3;
  assign t1_r4_c4_rr2 = t0_r4_c4_rr4;

  assign t2_r4_c4_rr0 = t1_r4_c4_rr0 + t1_r4_c4_rr1;
  assign t2_r4_c4_rr1 = t1_r4_c4_rr2;

  assign t3_r4_c4_rr0 = t2_r4_c4_rr0 + t2_r4_c4_rr1;

  assign c_4_4 = t3_r4_c4_rr0;
endmodule
