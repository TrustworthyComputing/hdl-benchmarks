module mmult (a_0_0, b_0_0, a_0_1, b_0_1, a_0_2, b_0_2, a_0_3, b_0_3, a_0_4, b_0_4, a_1_0, b_1_0, a_1_1, b_1_1, a_1_2, b_1_2, a_1_3, b_1_3, a_1_4, b_1_4, a_2_0, b_2_0, a_2_1, b_2_1, a_2_2, b_2_2, a_2_3, b_2_3, a_2_4, b_2_4, a_3_0, b_3_0, a_3_1, b_3_1, a_3_2, b_3_2, a_3_3, b_3_3, a_3_4, b_3_4, a_4_0, b_4_0, a_4_1, b_4_1, a_4_2, b_4_2, a_4_3, b_4_3, a_4_4, b_4_4, c_0_0, c_0_1, c_0_2, c_0_3, c_0_4, c_1_0, c_1_1, c_1_2, c_1_3, c_1_4, c_2_0, c_2_1, c_2_2, c_2_3, c_2_4, c_3_0, c_3_1, c_3_2, c_3_3, c_3_4, c_4_0, c_4_1, c_4_2, c_4_3, c_4_4);
  wire t0_r0_c0_rr0, t0_r0_c0_rr1, t0_r0_c0_rr2, t0_r0_c0_rr3, t0_r0_c0_rr4, t1_r0_c0_rr0, t1_r0_c0_rr1, t1_r0_c0_rr2, t2_r0_c0_rr0, t2_r0_c0_rr1, t3_r0_c0_rr0, t0_r0_c1_rr0, t0_r0_c1_rr1, t0_r0_c1_rr2, t0_r0_c1_rr3, t0_r0_c1_rr4, t1_r0_c1_rr0, t1_r0_c1_rr1, t1_r0_c1_rr2, t2_r0_c1_rr0, t2_r0_c1_rr1, t3_r0_c1_rr0, t0_r0_c2_rr0, t0_r0_c2_rr1, t0_r0_c2_rr2, t0_r0_c2_rr3, t0_r0_c2_rr4, t1_r0_c2_rr0, t1_r0_c2_rr1, t1_r0_c2_rr2, t2_r0_c2_rr0, t2_r0_c2_rr1, t3_r0_c2_rr0, t0_r0_c3_rr0, t0_r0_c3_rr1, t0_r0_c3_rr2, t0_r0_c3_rr3, t0_r0_c3_rr4, t1_r0_c3_rr0, t1_r0_c3_rr1, t1_r0_c3_rr2, t2_r0_c3_rr0, t2_r0_c3_rr1, t3_r0_c3_rr0, t0_r0_c4_rr0, t0_r0_c4_rr1, t0_r0_c4_rr2, t0_r0_c4_rr3, t0_r0_c4_rr4, t1_r0_c4_rr0, t1_r0_c4_rr1, t1_r0_c4_rr2, t2_r0_c4_rr0, t2_r0_c4_rr1, t3_r0_c4_rr0, t0_r1_c0_rr0, t0_r1_c0_rr1, t0_r1_c0_rr2, t0_r1_c0_rr3, t0_r1_c0_rr4, t1_r1_c0_rr0, t1_r1_c0_rr1, t1_r1_c0_rr2, t2_r1_c0_rr0, t2_r1_c0_rr1, t3_r1_c0_rr0, t0_r1_c1_rr0, t0_r1_c1_rr1, t0_r1_c1_rr2, t0_r1_c1_rr3, t0_r1_c1_rr4, t1_r1_c1_rr0, t1_r1_c1_rr1, t1_r1_c1_rr2, t2_r1_c1_rr0, t2_r1_c1_rr1, t3_r1_c1_rr0, t0_r1_c2_rr0, t0_r1_c2_rr1, t0_r1_c2_rr2, t0_r1_c2_rr3, t0_r1_c2_rr4, t1_r1_c2_rr0, t1_r1_c2_rr1, t1_r1_c2_rr2, t2_r1_c2_rr0, t2_r1_c2_rr1, t3_r1_c2_rr0, t0_r1_c3_rr0, t0_r1_c3_rr1, t0_r1_c3_rr2, t0_r1_c3_rr3, t0_r1_c3_rr4, t1_r1_c3_rr0, t1_r1_c3_rr1, t1_r1_c3_rr2, t2_r1_c3_rr0, t2_r1_c3_rr1, t3_r1_c3_rr0, t0_r1_c4_rr0, t0_r1_c4_rr1, t0_r1_c4_rr2, t0_r1_c4_rr3, t0_r1_c4_rr4, t1_r1_c4_rr0, t1_r1_c4_rr1, t1_r1_c4_rr2, t2_r1_c4_rr0, t2_r1_c4_rr1, t3_r1_c4_rr0, t0_r2_c0_rr0, t0_r2_c0_rr1, t0_r2_c0_rr2, t0_r2_c0_rr3, t0_r2_c0_rr4, t1_r2_c0_rr0, t1_r2_c0_rr1, t1_r2_c0_rr2, t2_r2_c0_rr0, t2_r2_c0_rr1, t3_r2_c0_rr0, t0_r2_c1_rr0, t0_r2_c1_rr1, t0_r2_c1_rr2, t0_r2_c1_rr3, t0_r2_c1_rr4, t1_r2_c1_rr0, t1_r2_c1_rr1, t1_r2_c1_rr2, t2_r2_c1_rr0, t2_r2_c1_rr1, t3_r2_c1_rr0, t0_r2_c2_rr0, t0_r2_c2_rr1, t0_r2_c2_rr2, t0_r2_c2_rr3, t0_r2_c2_rr4, t1_r2_c2_rr0, t1_r2_c2_rr1, t1_r2_c2_rr2, t2_r2_c2_rr0, t2_r2_c2_rr1, t3_r2_c2_rr0, t0_r2_c3_rr0, t0_r2_c3_rr1, t0_r2_c3_rr2, t0_r2_c3_rr3, t0_r2_c3_rr4, t1_r2_c3_rr0, t1_r2_c3_rr1, t1_r2_c3_rr2, t2_r2_c3_rr0, t2_r2_c3_rr1, t3_r2_c3_rr0, t0_r2_c4_rr0, t0_r2_c4_rr1, t0_r2_c4_rr2, t0_r2_c4_rr3, t0_r2_c4_rr4, t1_r2_c4_rr0, t1_r2_c4_rr1, t1_r2_c4_rr2, t2_r2_c4_rr0, t2_r2_c4_rr1, t3_r2_c4_rr0, t0_r3_c0_rr0, t0_r3_c0_rr1, t0_r3_c0_rr2, t0_r3_c0_rr3, t0_r3_c0_rr4, t1_r3_c0_rr0, t1_r3_c0_rr1, t1_r3_c0_rr2, t2_r3_c0_rr0, t2_r3_c0_rr1, t3_r3_c0_rr0, t0_r3_c1_rr0, t0_r3_c1_rr1, t0_r3_c1_rr2, t0_r3_c1_rr3, t0_r3_c1_rr4, t1_r3_c1_rr0, t1_r3_c1_rr1, t1_r3_c1_rr2, t2_r3_c1_rr0, t2_r3_c1_rr1, t3_r3_c1_rr0, t0_r3_c2_rr0, t0_r3_c2_rr1, t0_r3_c2_rr2, t0_r3_c2_rr3, t0_r3_c2_rr4, t1_r3_c2_rr0, t1_r3_c2_rr1, t1_r3_c2_rr2, t2_r3_c2_rr0, t2_r3_c2_rr1, t3_r3_c2_rr0, t0_r3_c3_rr0, t0_r3_c3_rr1, t0_r3_c3_rr2, t0_r3_c3_rr3, t0_r3_c3_rr4, t1_r3_c3_rr0, t1_r3_c3_rr1, t1_r3_c3_rr2, t2_r3_c3_rr0, t2_r3_c3_rr1, t3_r3_c3_rr0, t0_r3_c4_rr0, t0_r3_c4_rr1, t0_r3_c4_rr2, t0_r3_c4_rr3, t0_r3_c4_rr4, t1_r3_c4_rr0, t1_r3_c4_rr1, t1_r3_c4_rr2, t2_r3_c4_rr0, t2_r3_c4_rr1, t3_r3_c4_rr0, t0_r4_c0_rr0, t0_r4_c0_rr1, t0_r4_c0_rr2, t0_r4_c0_rr3, t0_r4_c0_rr4, t1_r4_c0_rr0, t1_r4_c0_rr1, t1_r4_c0_rr2, t2_r4_c0_rr0, t2_r4_c0_rr1, t3_r4_c0_rr0, t0_r4_c1_rr0, t0_r4_c1_rr1, t0_r4_c1_rr2, t0_r4_c1_rr3, t0_r4_c1_rr4, t1_r4_c1_rr0, t1_r4_c1_rr1, t1_r4_c1_rr2, t2_r4_c1_rr0, t2_r4_c1_rr1, t3_r4_c1_rr0, t0_r4_c2_rr0, t0_r4_c2_rr1, t0_r4_c2_rr2, t0_r4_c2_rr3, t0_r4_c2_rr4, t1_r4_c2_rr0, t1_r4_c2_rr1, t1_r4_c2_rr2, t2_r4_c2_rr0, t2_r4_c2_rr1, t3_r4_c2_rr0, t0_r4_c3_rr0, t0_r4_c3_rr1, t0_r4_c3_rr2, t0_r4_c3_rr3, t0_r4_c3_rr4, t1_r4_c3_rr0, t1_r4_c3_rr1, t1_r4_c3_rr2, t2_r4_c3_rr0, t2_r4_c3_rr1, t3_r4_c3_rr0, t0_r4_c4_rr0, t0_r4_c4_rr1, t0_r4_c4_rr2, t0_r4_c4_rr3, t0_r4_c4_rr4, t1_r4_c4_rr0, t1_r4_c4_rr1, t1_r4_c4_rr2, t2_r4_c4_rr0, t2_r4_c4_rr1, t3_r4_c4_rr0;
  input [15:0] a_0_0;
  input [15:0] b_0_0;
  input [15:0] a_0_1;
  input [15:0] b_0_1;
  input [15:0] a_0_2;
  input [15:0] b_0_2;
  input [15:0] a_0_3;
  input [15:0] b_0_3;
  input [15:0] a_0_4;
  input [15:0] b_0_4;
  input [15:0] a_1_0;
  input [15:0] b_1_0;
  input [15:0] a_1_1;
  input [15:0] b_1_1;
  input [15:0] a_1_2;
  input [15:0] b_1_2;
  input [15:0] a_1_3;
  input [15:0] b_1_3;
  input [15:0] a_1_4;
  input [15:0] b_1_4;
  input [15:0] a_2_0;
  input [15:0] b_2_0;
  input [15:0] a_2_1;
  input [15:0] b_2_1;
  input [15:0] a_2_2;
  input [15:0] b_2_2;
  input [15:0] a_2_3;
  input [15:0] b_2_3;
  input [15:0] a_2_4;
  input [15:0] b_2_4;
  input [15:0] a_3_0;
  input [15:0] b_3_0;
  input [15:0] a_3_1;
  input [15:0] b_3_1;
  input [15:0] a_3_2;
  input [15:0] b_3_2;
  input [15:0] a_3_3;
  input [15:0] b_3_3;
  input [15:0] a_3_4;
  input [15:0] b_3_4;
  input [15:0] a_4_0;
  input [15:0] b_4_0;
  input [15:0] a_4_1;
  input [15:0] b_4_1;
  input [15:0] a_4_2;
  input [15:0] b_4_2;
  input [15:0] a_4_3;
  input [15:0] b_4_3;
  input [15:0] a_4_4;
  input [15:0] b_4_4;
  output [15:0] c_0_0;
  output [15:0] c_0_1;
  output [15:0] c_0_2;
  output [15:0] c_0_3;
  output [15:0] c_0_4;
  output [15:0] c_1_0;
  output [15:0] c_1_1;
  output [15:0] c_1_2;
  output [15:0] c_1_3;
  output [15:0] c_1_4;
  output [15:0] c_2_0;
  output [15:0] c_2_1;
  output [15:0] c_2_2;
  output [15:0] c_2_3;
  output [15:0] c_2_4;
  output [15:0] c_3_0;
  output [15:0] c_3_1;
  output [15:0] c_3_2;
  output [15:0] c_3_3;
  output [15:0] c_3_4;
  output [15:0] c_4_0;
  output [15:0] c_4_1;
  output [15:0] c_4_2;
  output [15:0] c_4_3;
  output [15:0] c_4_4;
  mult m1(a_0_0, b_0_0, t0_r0_c0_rr0);
  mult m2(a_0_1, b_1_0, t0_r0_c0_rr1);
  mult m3(a_0_2, b_2_0, t0_r0_c0_rr2);
  mult m4(a_0_3, b_3_0, t0_r0_c0_rr3);
  mult m5(a_0_4, b_4_0, t0_r0_c0_rr4);
  add a6(t0_r0_c0_rr0, t0_r0_c0_rr1, t1_r0_c0_rr0);
  add a7(t0_r0_c0_rr2, t0_r0_c0_rr3, t1_r0_c0_rr1);
  copy c8(t0_r0_c0_rr4, t1_r0_c0_rr2);
  add a9(t1_r0_c0_rr0, t1_r0_c0_rr1, t2_r0_c0_rr0);
  copy c10(t1_r0_c0_rr2, t2_r0_c0_rr1);
  add a11(t2_r0_c0_rr0, t2_r0_c0_rr1, t3_r0_c0_rr0);
  copy c12(t3_r0_c0_rr0, c_0_0);
  mult m13(a_0_0, b_0_1, t0_r0_c1_rr0);
  mult m14(a_0_1, b_1_1, t0_r0_c1_rr1);
  mult m15(a_0_2, b_2_1, t0_r0_c1_rr2);
  mult m16(a_0_3, b_3_1, t0_r0_c1_rr3);
  mult m17(a_0_4, b_4_1, t0_r0_c1_rr4);
  add a18(t0_r0_c1_rr0, t0_r0_c1_rr1, t1_r0_c1_rr0);
  add a19(t0_r0_c1_rr2, t0_r0_c1_rr3, t1_r0_c1_rr1);
  copy c20(t0_r0_c1_rr4, t1_r0_c1_rr2);
  add a21(t1_r0_c1_rr0, t1_r0_c1_rr1, t2_r0_c1_rr0);
  copy c22(t1_r0_c1_rr2, t2_r0_c1_rr1);
  add a23(t2_r0_c1_rr0, t2_r0_c1_rr1, t3_r0_c1_rr0);
  copy c24(t3_r0_c1_rr0, c_0_1);
  mult m25(a_0_0, b_0_2, t0_r0_c2_rr0);
  mult m26(a_0_1, b_1_2, t0_r0_c2_rr1);
  mult m27(a_0_2, b_2_2, t0_r0_c2_rr2);
  mult m28(a_0_3, b_3_2, t0_r0_c2_rr3);
  mult m29(a_0_4, b_4_2, t0_r0_c2_rr4);
  add a30(t0_r0_c2_rr0, t0_r0_c2_rr1, t1_r0_c2_rr0);
  add a31(t0_r0_c2_rr2, t0_r0_c2_rr3, t1_r0_c2_rr1);
  copy c32(t0_r0_c2_rr4, t1_r0_c2_rr2);
  add a33(t1_r0_c2_rr0, t1_r0_c2_rr1, t2_r0_c2_rr0);
  copy c34(t1_r0_c2_rr2, t2_r0_c2_rr1);
  add a35(t2_r0_c2_rr0, t2_r0_c2_rr1, t3_r0_c2_rr0);
  copy c36(t3_r0_c2_rr0, c_0_2);
  mult m37(a_0_0, b_0_3, t0_r0_c3_rr0);
  mult m38(a_0_1, b_1_3, t0_r0_c3_rr1);
  mult m39(a_0_2, b_2_3, t0_r0_c3_rr2);
  mult m40(a_0_3, b_3_3, t0_r0_c3_rr3);
  mult m41(a_0_4, b_4_3, t0_r0_c3_rr4);
  add a42(t0_r0_c3_rr0, t0_r0_c3_rr1, t1_r0_c3_rr0);
  add a43(t0_r0_c3_rr2, t0_r0_c3_rr3, t1_r0_c3_rr1);
  copy c44(t0_r0_c3_rr4, t1_r0_c3_rr2);
  add a45(t1_r0_c3_rr0, t1_r0_c3_rr1, t2_r0_c3_rr0);
  copy c46(t1_r0_c3_rr2, t2_r0_c3_rr1);
  add a47(t2_r0_c3_rr0, t2_r0_c3_rr1, t3_r0_c3_rr0);
  copy c48(t3_r0_c3_rr0, c_0_3);
  mult m49(a_0_0, b_0_4, t0_r0_c4_rr0);
  mult m50(a_0_1, b_1_4, t0_r0_c4_rr1);
  mult m51(a_0_2, b_2_4, t0_r0_c4_rr2);
  mult m52(a_0_3, b_3_4, t0_r0_c4_rr3);
  mult m53(a_0_4, b_4_4, t0_r0_c4_rr4);
  add a54(t0_r0_c4_rr0, t0_r0_c4_rr1, t1_r0_c4_rr0);
  add a55(t0_r0_c4_rr2, t0_r0_c4_rr3, t1_r0_c4_rr1);
  copy c56(t0_r0_c4_rr4, t1_r0_c4_rr2);
  add a57(t1_r0_c4_rr0, t1_r0_c4_rr1, t2_r0_c4_rr0);
  copy c58(t1_r0_c4_rr2, t2_r0_c4_rr1);
  add a59(t2_r0_c4_rr0, t2_r0_c4_rr1, t3_r0_c4_rr0);
  copy c60(t3_r0_c4_rr0, c_0_4);
  mult m61(a_1_0, b_0_0, t0_r1_c0_rr0);
  mult m62(a_1_1, b_1_0, t0_r1_c0_rr1);
  mult m63(a_1_2, b_2_0, t0_r1_c0_rr2);
  mult m64(a_1_3, b_3_0, t0_r1_c0_rr3);
  mult m65(a_1_4, b_4_0, t0_r1_c0_rr4);
  add a66(t0_r1_c0_rr0, t0_r1_c0_rr1, t1_r1_c0_rr0);
  add a67(t0_r1_c0_rr2, t0_r1_c0_rr3, t1_r1_c0_rr1);
  copy c68(t0_r1_c0_rr4, t1_r1_c0_rr2);
  add a69(t1_r1_c0_rr0, t1_r1_c0_rr1, t2_r1_c0_rr0);
  copy c70(t1_r1_c0_rr2, t2_r1_c0_rr1);
  add a71(t2_r1_c0_rr0, t2_r1_c0_rr1, t3_r1_c0_rr0);
  copy c72(t3_r1_c0_rr0, c_1_0);
  mult m73(a_1_0, b_0_1, t0_r1_c1_rr0);
  mult m74(a_1_1, b_1_1, t0_r1_c1_rr1);
  mult m75(a_1_2, b_2_1, t0_r1_c1_rr2);
  mult m76(a_1_3, b_3_1, t0_r1_c1_rr3);
  mult m77(a_1_4, b_4_1, t0_r1_c1_rr4);
  add a78(t0_r1_c1_rr0, t0_r1_c1_rr1, t1_r1_c1_rr0);
  add a79(t0_r1_c1_rr2, t0_r1_c1_rr3, t1_r1_c1_rr1);
  copy c80(t0_r1_c1_rr4, t1_r1_c1_rr2);
  add a81(t1_r1_c1_rr0, t1_r1_c1_rr1, t2_r1_c1_rr0);
  copy c82(t1_r1_c1_rr2, t2_r1_c1_rr1);
  add a83(t2_r1_c1_rr0, t2_r1_c1_rr1, t3_r1_c1_rr0);
  copy c84(t3_r1_c1_rr0, c_1_1);
  mult m85(a_1_0, b_0_2, t0_r1_c2_rr0);
  mult m86(a_1_1, b_1_2, t0_r1_c2_rr1);
  mult m87(a_1_2, b_2_2, t0_r1_c2_rr2);
  mult m88(a_1_3, b_3_2, t0_r1_c2_rr3);
  mult m89(a_1_4, b_4_2, t0_r1_c2_rr4);
  add a90(t0_r1_c2_rr0, t0_r1_c2_rr1, t1_r1_c2_rr0);
  add a91(t0_r1_c2_rr2, t0_r1_c2_rr3, t1_r1_c2_rr1);
  copy c92(t0_r1_c2_rr4, t1_r1_c2_rr2);
  add a93(t1_r1_c2_rr0, t1_r1_c2_rr1, t2_r1_c2_rr0);
  copy c94(t1_r1_c2_rr2, t2_r1_c2_rr1);
  add a95(t2_r1_c2_rr0, t2_r1_c2_rr1, t3_r1_c2_rr0);
  copy c96(t3_r1_c2_rr0, c_1_2);
  mult m97(a_1_0, b_0_3, t0_r1_c3_rr0);
  mult m98(a_1_1, b_1_3, t0_r1_c3_rr1);
  mult m99(a_1_2, b_2_3, t0_r1_c3_rr2);
  mult m100(a_1_3, b_3_3, t0_r1_c3_rr3);
  mult m101(a_1_4, b_4_3, t0_r1_c3_rr4);
  add a102(t0_r1_c3_rr0, t0_r1_c3_rr1, t1_r1_c3_rr0);
  add a103(t0_r1_c3_rr2, t0_r1_c3_rr3, t1_r1_c3_rr1);
  copy c104(t0_r1_c3_rr4, t1_r1_c3_rr2);
  add a105(t1_r1_c3_rr0, t1_r1_c3_rr1, t2_r1_c3_rr0);
  copy c106(t1_r1_c3_rr2, t2_r1_c3_rr1);
  add a107(t2_r1_c3_rr0, t2_r1_c3_rr1, t3_r1_c3_rr0);
  copy c108(t3_r1_c3_rr0, c_1_3);
  mult m109(a_1_0, b_0_4, t0_r1_c4_rr0);
  mult m110(a_1_1, b_1_4, t0_r1_c4_rr1);
  mult m111(a_1_2, b_2_4, t0_r1_c4_rr2);
  mult m112(a_1_3, b_3_4, t0_r1_c4_rr3);
  mult m113(a_1_4, b_4_4, t0_r1_c4_rr4);
  add a114(t0_r1_c4_rr0, t0_r1_c4_rr1, t1_r1_c4_rr0);
  add a115(t0_r1_c4_rr2, t0_r1_c4_rr3, t1_r1_c4_rr1);
  copy c116(t0_r1_c4_rr4, t1_r1_c4_rr2);
  add a117(t1_r1_c4_rr0, t1_r1_c4_rr1, t2_r1_c4_rr0);
  copy c118(t1_r1_c4_rr2, t2_r1_c4_rr1);
  add a119(t2_r1_c4_rr0, t2_r1_c4_rr1, t3_r1_c4_rr0);
  copy c120(t3_r1_c4_rr0, c_1_4);
  mult m121(a_2_0, b_0_0, t0_r2_c0_rr0);
  mult m122(a_2_1, b_1_0, t0_r2_c0_rr1);
  mult m123(a_2_2, b_2_0, t0_r2_c0_rr2);
  mult m124(a_2_3, b_3_0, t0_r2_c0_rr3);
  mult m125(a_2_4, b_4_0, t0_r2_c0_rr4);
  add a126(t0_r2_c0_rr0, t0_r2_c0_rr1, t1_r2_c0_rr0);
  add a127(t0_r2_c0_rr2, t0_r2_c0_rr3, t1_r2_c0_rr1);
  copy c128(t0_r2_c0_rr4, t1_r2_c0_rr2);
  add a129(t1_r2_c0_rr0, t1_r2_c0_rr1, t2_r2_c0_rr0);
  copy c130(t1_r2_c0_rr2, t2_r2_c0_rr1);
  add a131(t2_r2_c0_rr0, t2_r2_c0_rr1, t3_r2_c0_rr0);
  copy c132(t3_r2_c0_rr0, c_2_0);
  mult m133(a_2_0, b_0_1, t0_r2_c1_rr0);
  mult m134(a_2_1, b_1_1, t0_r2_c1_rr1);
  mult m135(a_2_2, b_2_1, t0_r2_c1_rr2);
  mult m136(a_2_3, b_3_1, t0_r2_c1_rr3);
  mult m137(a_2_4, b_4_1, t0_r2_c1_rr4);
  add a138(t0_r2_c1_rr0, t0_r2_c1_rr1, t1_r2_c1_rr0);
  add a139(t0_r2_c1_rr2, t0_r2_c1_rr3, t1_r2_c1_rr1);
  copy c140(t0_r2_c1_rr4, t1_r2_c1_rr2);
  add a141(t1_r2_c1_rr0, t1_r2_c1_rr1, t2_r2_c1_rr0);
  copy c142(t1_r2_c1_rr2, t2_r2_c1_rr1);
  add a143(t2_r2_c1_rr0, t2_r2_c1_rr1, t3_r2_c1_rr0);
  copy c144(t3_r2_c1_rr0, c_2_1);
  mult m145(a_2_0, b_0_2, t0_r2_c2_rr0);
  mult m146(a_2_1, b_1_2, t0_r2_c2_rr1);
  mult m147(a_2_2, b_2_2, t0_r2_c2_rr2);
  mult m148(a_2_3, b_3_2, t0_r2_c2_rr3);
  mult m149(a_2_4, b_4_2, t0_r2_c2_rr4);
  add a150(t0_r2_c2_rr0, t0_r2_c2_rr1, t1_r2_c2_rr0);
  add a151(t0_r2_c2_rr2, t0_r2_c2_rr3, t1_r2_c2_rr1);
  copy c152(t0_r2_c2_rr4, t1_r2_c2_rr2);
  add a153(t1_r2_c2_rr0, t1_r2_c2_rr1, t2_r2_c2_rr0);
  copy c154(t1_r2_c2_rr2, t2_r2_c2_rr1);
  add a155(t2_r2_c2_rr0, t2_r2_c2_rr1, t3_r2_c2_rr0);
  copy c156(t3_r2_c2_rr0, c_2_2);
  mult m157(a_2_0, b_0_3, t0_r2_c3_rr0);
  mult m158(a_2_1, b_1_3, t0_r2_c3_rr1);
  mult m159(a_2_2, b_2_3, t0_r2_c3_rr2);
  mult m160(a_2_3, b_3_3, t0_r2_c3_rr3);
  mult m161(a_2_4, b_4_3, t0_r2_c3_rr4);
  add a162(t0_r2_c3_rr0, t0_r2_c3_rr1, t1_r2_c3_rr0);
  add a163(t0_r2_c3_rr2, t0_r2_c3_rr3, t1_r2_c3_rr1);
  copy c164(t0_r2_c3_rr4, t1_r2_c3_rr2);
  add a165(t1_r2_c3_rr0, t1_r2_c3_rr1, t2_r2_c3_rr0);
  copy c166(t1_r2_c3_rr2, t2_r2_c3_rr1);
  add a167(t2_r2_c3_rr0, t2_r2_c3_rr1, t3_r2_c3_rr0);
  copy c168(t3_r2_c3_rr0, c_2_3);
  mult m169(a_2_0, b_0_4, t0_r2_c4_rr0);
  mult m170(a_2_1, b_1_4, t0_r2_c4_rr1);
  mult m171(a_2_2, b_2_4, t0_r2_c4_rr2);
  mult m172(a_2_3, b_3_4, t0_r2_c4_rr3);
  mult m173(a_2_4, b_4_4, t0_r2_c4_rr4);
  add a174(t0_r2_c4_rr0, t0_r2_c4_rr1, t1_r2_c4_rr0);
  add a175(t0_r2_c4_rr2, t0_r2_c4_rr3, t1_r2_c4_rr1);
  copy c176(t0_r2_c4_rr4, t1_r2_c4_rr2);
  add a177(t1_r2_c4_rr0, t1_r2_c4_rr1, t2_r2_c4_rr0);
  copy c178(t1_r2_c4_rr2, t2_r2_c4_rr1);
  add a179(t2_r2_c4_rr0, t2_r2_c4_rr1, t3_r2_c4_rr0);
  copy c180(t3_r2_c4_rr0, c_2_4);
  mult m181(a_3_0, b_0_0, t0_r3_c0_rr0);
  mult m182(a_3_1, b_1_0, t0_r3_c0_rr1);
  mult m183(a_3_2, b_2_0, t0_r3_c0_rr2);
  mult m184(a_3_3, b_3_0, t0_r3_c0_rr3);
  mult m185(a_3_4, b_4_0, t0_r3_c0_rr4);
  add a186(t0_r3_c0_rr0, t0_r3_c0_rr1, t1_r3_c0_rr0);
  add a187(t0_r3_c0_rr2, t0_r3_c0_rr3, t1_r3_c0_rr1);
  copy c188(t0_r3_c0_rr4, t1_r3_c0_rr2);
  add a189(t1_r3_c0_rr0, t1_r3_c0_rr1, t2_r3_c0_rr0);
  copy c190(t1_r3_c0_rr2, t2_r3_c0_rr1);
  add a191(t2_r3_c0_rr0, t2_r3_c0_rr1, t3_r3_c0_rr0);
  copy c192(t3_r3_c0_rr0, c_3_0);
  mult m193(a_3_0, b_0_1, t0_r3_c1_rr0);
  mult m194(a_3_1, b_1_1, t0_r3_c1_rr1);
  mult m195(a_3_2, b_2_1, t0_r3_c1_rr2);
  mult m196(a_3_3, b_3_1, t0_r3_c1_rr3);
  mult m197(a_3_4, b_4_1, t0_r3_c1_rr4);
  add a198(t0_r3_c1_rr0, t0_r3_c1_rr1, t1_r3_c1_rr0);
  add a199(t0_r3_c1_rr2, t0_r3_c1_rr3, t1_r3_c1_rr1);
  copy c200(t0_r3_c1_rr4, t1_r3_c1_rr2);
  add a201(t1_r3_c1_rr0, t1_r3_c1_rr1, t2_r3_c1_rr0);
  copy c202(t1_r3_c1_rr2, t2_r3_c1_rr1);
  add a203(t2_r3_c1_rr0, t2_r3_c1_rr1, t3_r3_c1_rr0);
  copy c204(t3_r3_c1_rr0, c_3_1);
  mult m205(a_3_0, b_0_2, t0_r3_c2_rr0);
  mult m206(a_3_1, b_1_2, t0_r3_c2_rr1);
  mult m207(a_3_2, b_2_2, t0_r3_c2_rr2);
  mult m208(a_3_3, b_3_2, t0_r3_c2_rr3);
  mult m209(a_3_4, b_4_2, t0_r3_c2_rr4);
  add a210(t0_r3_c2_rr0, t0_r3_c2_rr1, t1_r3_c2_rr0);
  add a211(t0_r3_c2_rr2, t0_r3_c2_rr3, t1_r3_c2_rr1);
  copy c212(t0_r3_c2_rr4, t1_r3_c2_rr2);
  add a213(t1_r3_c2_rr0, t1_r3_c2_rr1, t2_r3_c2_rr0);
  copy c214(t1_r3_c2_rr2, t2_r3_c2_rr1);
  add a215(t2_r3_c2_rr0, t2_r3_c2_rr1, t3_r3_c2_rr0);
  copy c216(t3_r3_c2_rr0, c_3_2);
  mult m217(a_3_0, b_0_3, t0_r3_c3_rr0);
  mult m218(a_3_1, b_1_3, t0_r3_c3_rr1);
  mult m219(a_3_2, b_2_3, t0_r3_c3_rr2);
  mult m220(a_3_3, b_3_3, t0_r3_c3_rr3);
  mult m221(a_3_4, b_4_3, t0_r3_c3_rr4);
  add a222(t0_r3_c3_rr0, t0_r3_c3_rr1, t1_r3_c3_rr0);
  add a223(t0_r3_c3_rr2, t0_r3_c3_rr3, t1_r3_c3_rr1);
  copy c224(t0_r3_c3_rr4, t1_r3_c3_rr2);
  add a225(t1_r3_c3_rr0, t1_r3_c3_rr1, t2_r3_c3_rr0);
  copy c226(t1_r3_c3_rr2, t2_r3_c3_rr1);
  add a227(t2_r3_c3_rr0, t2_r3_c3_rr1, t3_r3_c3_rr0);
  copy c228(t3_r3_c3_rr0, c_3_3);
  mult m229(a_3_0, b_0_4, t0_r3_c4_rr0);
  mult m230(a_3_1, b_1_4, t0_r3_c4_rr1);
  mult m231(a_3_2, b_2_4, t0_r3_c4_rr2);
  mult m232(a_3_3, b_3_4, t0_r3_c4_rr3);
  mult m233(a_3_4, b_4_4, t0_r3_c4_rr4);
  add a234(t0_r3_c4_rr0, t0_r3_c4_rr1, t1_r3_c4_rr0);
  add a235(t0_r3_c4_rr2, t0_r3_c4_rr3, t1_r3_c4_rr1);
  copy c236(t0_r3_c4_rr4, t1_r3_c4_rr2);
  add a237(t1_r3_c4_rr0, t1_r3_c4_rr1, t2_r3_c4_rr0);
  copy c238(t1_r3_c4_rr2, t2_r3_c4_rr1);
  add a239(t2_r3_c4_rr0, t2_r3_c4_rr1, t3_r3_c4_rr0);
  copy c240(t3_r3_c4_rr0, c_3_4);
  mult m241(a_4_0, b_0_0, t0_r4_c0_rr0);
  mult m242(a_4_1, b_1_0, t0_r4_c0_rr1);
  mult m243(a_4_2, b_2_0, t0_r4_c0_rr2);
  mult m244(a_4_3, b_3_0, t0_r4_c0_rr3);
  mult m245(a_4_4, b_4_0, t0_r4_c0_rr4);
  add a246(t0_r4_c0_rr0, t0_r4_c0_rr1, t1_r4_c0_rr0);
  add a247(t0_r4_c0_rr2, t0_r4_c0_rr3, t1_r4_c0_rr1);
  copy c248(t0_r4_c0_rr4, t1_r4_c0_rr2);
  add a249(t1_r4_c0_rr0, t1_r4_c0_rr1, t2_r4_c0_rr0);
  copy c250(t1_r4_c0_rr2, t2_r4_c0_rr1);
  add a251(t2_r4_c0_rr0, t2_r4_c0_rr1, t3_r4_c0_rr0);
  copy c252(t3_r4_c0_rr0, c_4_0);
  mult m253(a_4_0, b_0_1, t0_r4_c1_rr0);
  mult m254(a_4_1, b_1_1, t0_r4_c1_rr1);
  mult m255(a_4_2, b_2_1, t0_r4_c1_rr2);
  mult m256(a_4_3, b_3_1, t0_r4_c1_rr3);
  mult m257(a_4_4, b_4_1, t0_r4_c1_rr4);
  add a258(t0_r4_c1_rr0, t0_r4_c1_rr1, t1_r4_c1_rr0);
  add a259(t0_r4_c1_rr2, t0_r4_c1_rr3, t1_r4_c1_rr1);
  copy c260(t0_r4_c1_rr4, t1_r4_c1_rr2);
  add a261(t1_r4_c1_rr0, t1_r4_c1_rr1, t2_r4_c1_rr0);
  copy c262(t1_r4_c1_rr2, t2_r4_c1_rr1);
  add a263(t2_r4_c1_rr0, t2_r4_c1_rr1, t3_r4_c1_rr0);
  copy c264(t3_r4_c1_rr0, c_4_1);
  mult m265(a_4_0, b_0_2, t0_r4_c2_rr0);
  mult m266(a_4_1, b_1_2, t0_r4_c2_rr1);
  mult m267(a_4_2, b_2_2, t0_r4_c2_rr2);
  mult m268(a_4_3, b_3_2, t0_r4_c2_rr3);
  mult m269(a_4_4, b_4_2, t0_r4_c2_rr4);
  add a270(t0_r4_c2_rr0, t0_r4_c2_rr1, t1_r4_c2_rr0);
  add a271(t0_r4_c2_rr2, t0_r4_c2_rr3, t1_r4_c2_rr1);
  copy c272(t0_r4_c2_rr4, t1_r4_c2_rr2);
  add a273(t1_r4_c2_rr0, t1_r4_c2_rr1, t2_r4_c2_rr0);
  copy c274(t1_r4_c2_rr2, t2_r4_c2_rr1);
  add a275(t2_r4_c2_rr0, t2_r4_c2_rr1, t3_r4_c2_rr0);
  copy c276(t3_r4_c2_rr0, c_4_2);
  mult m277(a_4_0, b_0_3, t0_r4_c3_rr0);
  mult m278(a_4_1, b_1_3, t0_r4_c3_rr1);
  mult m279(a_4_2, b_2_3, t0_r4_c3_rr2);
  mult m280(a_4_3, b_3_3, t0_r4_c3_rr3);
  mult m281(a_4_4, b_4_3, t0_r4_c3_rr4);
  add a282(t0_r4_c3_rr0, t0_r4_c3_rr1, t1_r4_c3_rr0);
  add a283(t0_r4_c3_rr2, t0_r4_c3_rr3, t1_r4_c3_rr1);
  copy c284(t0_r4_c3_rr4, t1_r4_c3_rr2);
  add a285(t1_r4_c3_rr0, t1_r4_c3_rr1, t2_r4_c3_rr0);
  copy c286(t1_r4_c3_rr2, t2_r4_c3_rr1);
  add a287(t2_r4_c3_rr0, t2_r4_c3_rr1, t3_r4_c3_rr0);
  copy c288(t3_r4_c3_rr0, c_4_3);
  mult m289(a_4_0, b_0_4, t0_r4_c4_rr0);
  mult m290(a_4_1, b_1_4, t0_r4_c4_rr1);
  mult m291(a_4_2, b_2_4, t0_r4_c4_rr2);
  mult m292(a_4_3, b_3_4, t0_r4_c4_rr3);
  mult m293(a_4_4, b_4_4, t0_r4_c4_rr4);
  add a294(t0_r4_c4_rr0, t0_r4_c4_rr1, t1_r4_c4_rr0);
  add a295(t0_r4_c4_rr2, t0_r4_c4_rr3, t1_r4_c4_rr1);
  copy c296(t0_r4_c4_rr4, t1_r4_c4_rr2);
  add a297(t1_r4_c4_rr0, t1_r4_c4_rr1, t2_r4_c4_rr0);
  copy c298(t1_r4_c4_rr2, t2_r4_c4_rr1);
  add a299(t2_r4_c4_rr0, t2_r4_c4_rr1, t3_r4_c4_rr0);
  copy c300(t3_r4_c4_rr0, c_4_4);

endmodule
