module c3540(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9);
  wire 0000, 0001, 0002, 0003, 0004, 0005, 0006, 0007, 0008, 0009, 0010, 0011, 0012, 0013, 0014, 0015, 0016, 0017, 0018, 0019, 0020, 0021, 0022, 0023, 0024, 0025, 0026, 0027, 0028, 0029, 0030, 0031, 0032, 0033, 0034, 0035, 0036, 0037, 0038, 0039, 0040, 0041, 0042, 0043, 0044, 0045, 0046, 0047, 0048, 0049, 0050, 0051, 0052, 0053, 0054, 0055, 0056, 0057, 0058, 0059, 0060, 0061, 0062, 0063, 0064, 0065, 0066, 0067, 0068, 0069, 0070, 0071, 0072, 0073, 0074, 0075, 0076, 0077, 0078, 0079, 0080, 0081, 0082, 0083, 0084, 0085, 0086, 0087, 0088, 0089, 0090, 0091, 0092, 0093, 0094, 0095, 0096, 0097, 0098, 0099, 0100, 0101, 0102, 0103, 0104, 0105, 0106, 0107, 0108, 0109, 0110, 0111, 0112, 0113, 0114, 0115, 0116, 0117, 0118, 0119, 0120, 0121, 0122, 0123, 0124, 0125, 0126, 0127, 0128, 0129, 0130, 0131, 0132, 0133, 0134, 0135, 0136, 0137, 0138, 0139, 0140, 0141, 0142, 0143, 0144, 0145, 0146, 0147, 0148, 0149, 0150, 0151, 0152, 0153, 0154, 0155, 0156, 0157, 0158, 0159, 0160, 0161, 0162, 0163, 0164, 0165, 0166, 0167, 0168, 0169, 0170, 0171, 0172, 0173, 0174, 0175, 0176, 0177, 0178, 0179, 0180, 0181, 0182, 0183, 0184, 0185, 0186, 0187, 0188, 0189, 0190, 0191, 0192, 0193, 0194, 0195, 0196, 0197, 0198, 0199, 0200, 0201, 0202, 0203, 0204, 0205, 0206, 0207, 0208, 0209, 0210, 0211, 0212, 0213, 0214, 0215, 0216, 0217, 0218, 0219, 0220, 0221, 0222, 0223, 0224, 0225, 0226, 0227, 0228, 0229, 0230, 0231, 0232, 0233, 0234, 0235, 0236, 0237, 0238, 0239, 0240, 0241, 0242, 0243, 0244, 0245, 0246, 0247, 0248, 0249, 0250, 0251, 0252, 0253, 0254, 0255, 0256, 0257, 0258, 0259, 0260, 0261, 0262, 0263, 0264, 0265, 0266, 0267, 0268, 0269, 0270, 0271, 0272, 0273, 0274, 0275, 0276, 0277, 0278, 0279, 0280, 0281, 0282, 0283, 0284, 0285, 0286, 0287, 0288, 0289, 0290, 0291, 0292, 0293, 0294, 0295, 0296, 0297, 0298, 0299, 0300, 0301, 0302, 0303, 0304, 0305, 0306, 0307, 0308, 0309, 0310, 0311, 0312, 0313, 0314, 0315, 0316, 0317, 0318, 0319, 0320, 0321, 0322, 0323, 0324, 0325, 0326, 0327, 0328, 0329, 0330, 0331, 0332, 0333, 0334, 0335, 0336, 0337, 0338, 0339, 0340, 0341, 0342, 0343, 0344, 0345, 0346, 0347, 0348, 0349, 0350, 0351, 0352, 0353, 0354, 0355, 0356, 0357, 0358, 0359, 0360, 0361, 0362, 0363, 0364, 0365, 0366, 0367, 0368, 0369, 0370, 0371, 0372, 0373, 0374, 0375, 0376, 0377, 0378, 0379, 0380, 0381, 0382, 0383, 0384, 0385, 0386, 0387, 0388, 0389, 0390, 0391, 0392, 0393, 0394, 0395, 0396, 0397, 0398, 0399, 0400, 0401, 0402, 0403, 0404, 0405, 0406, 0407, 0408, 0409, 0410, 0411, 0412, 0413, 0414, 0415, 0416, 0417, 0418, 0419, 0420, 0421, 0422, 0423, 0424, 0425, 0426, 0427, 0428, 0429, 0430, 0431, 0432, 0433, 0434, 0435, 0436, 0437, 0438, 0439, 0440, 0441, 0442, 0443, 0444, 0445, 0446, 0447, 0448, 0449, 0450, 0451, 0452, 0453, 0454, 0455, 0456, 0457, 0458, 0459, 0460, 0461, 0462, 0463, 0464, 0465, 0466, 0467, 0468, 0469, 0470, 0471, 0472, 0473, 0474, 0475, 0476, 0477, 0478, 0479, 0480, 0481, 0482, 0483, 0484, 0485, 0486, 0487, 0488, 0489, 0490, 0491, 0492, 0493, 0494, 0495, 0496, 0497, 0498, 0499, 0500, 0501, 0502, 0503, 0504, 0505, 0506, 0507, 0508, 0509, 0510, 0511, 0512, 0513, 0514, 0515, 0516, 0517, 0518, 0519, 0520, 0521, 0522, 0523, 0524, 0525, 0526, 0527, 0528, 0529, 0530, 0531, 0532, 0533, 0534, 0535, 0536, 0537, 0538, 0539, 0540, 0541, 0542, 0543, 0544, 0545, 0546, 0547, 0548, 0549, 0550, 0551, 0552, 0553, 0554, 0555, 0556, 0557, 0558, 0559, 0560, 0561, 0562, 0563, 0564, 0565, 0566, 0567, 0568, 0569, 0570, 0571, 0572, 0573, 0574, 0575, 0576, 0577, 0578, 0579, 0580, 0581, 0582, 0583, 0584, 0585, 0586, 0587, 0588, 0589, 0590, 0591, 0592, 0593, 0594, 0595, 0596, 0597, 0598, 0599, 0600, 0601, 0602, 0603, 0604, 0605, 0606, 0607, 0608, 0609, 0610, 0611, 0612, 0613, 0614, 0615, 0616, 0617, 0618, 0619, 0620, 0621, 0622, 0623, 0624, 0625, 0626, 0627, 0628, 0629, 0630, 0631, 0632, 0633, 0634, 0635, 0636, 0637, 0638, 0639, 0640, 0641, 0642, 0643, 0644, 0645, 0646, 0647, 0648, 0649, 0650, 0651, 0652, 0653, 0654, 0655, 0656, 0657, 0658, 0659, 0660, 0661, 0662, 0663, 0664, 0665, 0666, 0667, 0668, 0669, 0670, 0671, 0672, 0673, 0674, 0675, 0676, 0677, 0678, 0679, 0680, 0681, 0682, 0683, 0684, 0685, 0686, 0687, 0688, 0689, 0690, 0691, 0692, 0693, 0694, 0695, 0696, 0697, 0698, 0699, 0700, 0701, 0702, 0703, 0704, 0705, 0706, 0707, 0708, 0709, 0710, 0711, 0712, 0713, 0714, 0715, 0716, 0717, 0718, 0719, 0720, 0721, 0722, 0723, 0724, 0725, 0726, 0727, 0728, 0729, 0730, 0731, 0732, 0733, 0734, 0735, 0736, 0737, 0738, 0739, 0740, 0741, 0742, 0743, 0744, 0745, 0746, 0747, 0748, 0749, 0750, 0751, 0752, 0753, 0754, 0755, 0756, 0757, 0758, 0759, 0760, 0761, 0762, 0763, 0764, 0765, 0766, 0767, 0768, 0769, 0770, 0771, 0772, 0773, 0774, 0775, 0776, 0777, 0778, 0779, 0780, 0781, 0782, 0783, 0784, 0785, 0786, 0787, 0788, 0789, 0790, 0791, 0792, 0793, 0794, 0795, 0796, 0797, 0798, 0799, 0800, 0801, 0802, 0803, 0804, 0805, 0806, 0807, 0808, 0809, 0810, 0811, 0812, 0813, 0814, 0815, 0816, 0817, 0818, 0819, 0820, 0821, 0822, 0823, 0824, 0825, 0826, 0827, 0828, 0829, 0830, 0831, 0832, 0833, 0834, 0835, 0836, 0837, 0838, 0839, 0840, 0841, 0842, 0843, 0844, 0845, 0846, 0847, 0848, 0849, 0850, 0851, 0852, 0853, 0854, 0855, 0856, 0857, 0858, 0859, 0860, 0861, 0862, 0863, 0864, 0865, 0866, 0867, 0868, 0869, 0870, 0871, 0872, 0873, 0874, 0875, 0876, 0877, 0878, 0879, 0880, 0881, 0882, 0883, 0884, 0885, 0886, 0887, 0888, 0889, 0890, 0891, 0892, 0893, 0894, 0895, 0896, 0897, 0898, 0899, 0900, 0901, 0902, 0903, 0904, 0905, 0906, 0907, 0908, 0909, 0910, 0911, 0912, 0913, 0914, 0915, 0916, 0917, 0918, 0919, 0920, 0921, 0922, 0923, 0924, 0925, 0926, 0927, 0928, 0929, 0930, 0931, 0932, 0933, 0934, 0935, 0936, 0937, 0938, 0939, 0940, 0941, 0942, 0943, 0944, 0945, 0946, 0947, 0948, 0949, 0950, 0951, 0952, 0953, 0954, 0955, 0956, 0957, 0958, 0959, 0960, 0961, 0962, 0963, 0964, 0965, 0966, 0967, 0968, 0969, 0970, 0971, 0972, 0973, 0974, 0975, 0976, 0977, 0978, 0979, 0980, 0981, 0982, 0983, 0984, 0985, 0986, 0987, 0988, 0989, 0990, 0991, 0992, 0993, 0994, 0995, 0996, 0997, 0998, 0999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, G1022, G2943, G2974, G2985, G3005, G3030, G3100, G3135, G3195, G3202, G3226, G3257, G3265, G3266, G3267, G3275, G3281, G3294, G3300, G3301, G3311, G3312, G3320, G3332, G3341, G3342, G3343, G3345, G3373, G3376, G3379, G3394, G3515, G3516, G722, G723, G724, G725, G731, G734, G735, G736, G739, G742, G745, G749, G781, G786, G791, G792, G793, G794, G795, G796, G797, G798, G799, G816, G831, G882, G883, G890, G891, G892, G893, G894, G897, G898, G901, G904, G907, G910, G913, G916, G919, G922, G925;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540;
  lut lut_gate1(0x07, 1067, 1050, 1062, 1049);
  lut lut_gate2(0x40, 1061, 1051, 1059, 1050);
  lut lut_gate3(0xe0, 1052, 1058, G10, 1051);
  lut lut_gate4(0x0e, 1053, 1057, G7, 1052);
  lut lut_gate5(0x1, G12, 1054, 1053);
  lut lut_gate6(0x4, 1056, 1055, 1054);
  lut lut_gate7(0x8, G26, G3, 1055);
  lut lut_gate8(0x1f, G3, G25, G24, 1056);
  lut lut_gate9(0x8, G26, 1056, 1057);
  lut lut_gate10(0x01, 1056, G26, G24, 1058);
  lut lut_gate11(0x1, G13, 1060, 1059);
  lut lut_gate12(0x40, G25, 1055, G24, 1060);
  lut lut_gate13(0x0, G4, 1058, G22, 1061);
  lut lut_gate14(0xe0, 1063, 1066, G8, 1062);
  lut lut_gate15(0x0e, 1064, 1065, G11, 1063);
  lut lut_gate16(0x1, G9, 1060, 1064);
  lut lut_gate17(0x10, 1055, G25, G24, 1065);
  lut lut_gate18(0x4, 1056, G26, 1066);
  lut lut_gate19(0x80, 0687, 1071, 1068, 1067);
  lut lut_gate20(0x10, G4, 1070, 1069, 1068);
  lut lut_gate21(0x4, G44, 1066, 1069);
  lut lut_gate22(0x0e, 1058, G42, G46, 1070);
  lut lut_gate23(0x0, 0686, 1065, G41, 1071);
  lut lut_gate24(0x4, G40, 1054, 0686);
  lut lut_gate25(0x0, 0688, 1057, G45, 0687);
  lut lut_gate26(0x0e, 1060, G39, G43, 0688);
  lut lut_gate27(0x4, 0690, G6, 0689);
  lut lut_gate28(0x8, G5, 0691, 0690);
  lut lut_gate29(0x01, G3, G1, G2, 0691);
  lut lut_gate30(0x4, G2, G1, 0692);
  lut lut_gate31(0x4b, 0694, 0718, 0695, 0693);
  lut lut_gate32(0xc5, 0695, 0716, 0705, 0694);
  lut lut_gate33(0x0, 0702, 0696, G14, 0695);
  lut lut_gate34(0x35, 0697, 0700, G3, 0696);
  lut lut_gate35(0x1, 0699, 0698, 0697);
  lut lut_gate36(0x8, G1, G2, 0698);
  lut lut_gate37(0x80, G4, G3, G1, 0699);
  lut lut_gate38(0x0, 0701, G1, G4, 0700);
  lut lut_gate39(0x40, G3, G2, G1, 0701);
  lut lut_gate40(0x0b, 0703, 0701, G14, 0702);
  lut lut_gate41(0x40, 0698, 0704, G3, 0703);
  lut lut_gate42(0xc5, G4, G39, G12, 0704);
  lut lut_gate43(0x01, 0715, 0710, 0706, 0705);
  lut lut_gate44(0x8, G38, 0709, 0706);
  lut lut_gate45(0x4, 0698, 0708, 0707);
  lut lut_gate46(0x8, G5, G4, 0708);
  lut lut_gate47(0x01, G6, G5, G1, 0709);
  lut lut_gate48(0x0, 0707, 0711, 0713, 0710);
  lut lut_gate49(0x8, G35, 0712, 0711);
  lut lut_gate50(0x1, G49, G4, 0712);
  lut lut_gate51(0x0, 0714, 0709, G37, 0713);
  lut lut_gate52(0xca, G4, G36, G41, 0714);
  lut lut_gate53(0x1, G24, G23, 0715);
  lut lut_gate54(0x01, 0717, 0710, 0706, 0716);
  lut lut_gate55(0x1, G26, G25, 0717);
  lut lut_gate56(0x8, 0719, 0691, 0718);
  lut lut_gate57(0x8, G48, G27, 0719);
  lut lut_gate58(0x4, 0721, G2, 0720);
  lut lut_gate59(0x4, G4, G3, 0721);
  lut lut_gate60(0xf4, 0722, 0783, 0781, G3529);
  lut lut_gate61(0x41, 0723, 0766, 0689, 0722);
  lut lut_gate62(0x4, G47, 0724, 0723);
  lut lut_gate63(0x1, 0740, 1045, 0724);
  lut lut_gate64(0x1, 0710, 0706, 0725);
  lut lut_gate65(0x07, 0707, 0727, 0730, 0726);
  lut lut_gate66(0x0, 0729, 0728, G34, 0727);
  lut lut_gate67(0x1, G6, G1, 0728);
  lut lut_gate68(0x53, G4, G14, G33, 0729);
  lut lut_gate69(0x07, 0731, 0712, G32, 0730);
  lut lut_gate70(0x10, G38, G6, G1, 0731);
  lut lut_gate71(0x0, 0707, 0733, 0734, 0732);
  lut lut_gate72(0x4, G36, 0709, 0733);
  lut lut_gate73(0x70, 0735, 0712, G34, 0734);
  lut lut_gate74(0x35, G4, G35, G40, 0735);
  lut lut_gate75(0x0, 0707, 0737, 0738, 0736);
  lut lut_gate76(0x8, G33, 0712, 0737);
  lut lut_gate77(0x0, 0739, 0709, G35, 0738);
  lut lut_gate78(0xca, G4, G34, G39, 0739);
  lut lut_gate79(0x80, 0718, 0694, 0741, 0740);
  lut lut_gate80(0x80, 0761, 0751, 0742, 0741);
  lut lut_gate81(0xc5, 0743, 0750, 0749, 0742);
  lut lut_gate82(0x01, 0747, 0745, 0744, 0743);
  lut lut_gate83(0x80, G13, 0700, 0697, 0744);
  lut lut_gate84(0x10, G3, G13, 0746, 0745);
  lut lut_gate85(0x1, G2, 0699, 0746);
  lut lut_gate86(0x40, 0698, 0748, G3, 0747);
  lut lut_gate87(0xc5, G4, G14, G11, 0748);
  lut lut_gate88(0x01, 0715, 0732, 0706, 0749);
  lut lut_gate89(0x01, 0717, 0732, 0706, 0750);
  lut lut_gate90(0xc5, 0752, 0760, 0759, 0751);
  lut lut_gate91(0x01, 0758, 0757, 0753, 0752);
  lut lut_gate92(0x10, 0754, 0756, 0697, 0753);
  lut lut_gate93(0x0b, 0755, 0721, G13, 0754);
  lut lut_gate94(0x90, G3, G13, G12, 0755);
  lut lut_gate95(0x01, G10, G4, G3, 0756);
  lut lut_gate96(0x80, G12, 0700, 0697, 0757);
  lut lut_gate97(0x4, 0701, G12, 0758);
  lut lut_gate98(0x01, 0715, 0736, 0706, 0759);
  lut lut_gate99(0x01, 0717, 0736, 0706, 0760);
  lut lut_gate100(0xc5, 1009, 0765, 0764, 0761);
  lut lut_gate101(0x01, G13, G11, G12, 0762);
  lut lut_gate102(0x4, 0701, G11, 0763);
  lut lut_gate103(0x1, 0715, 0726, 0764);
  lut lut_gate104(0x1, 0717, 0726, 0765);
  lut lut_gate105(0xe1, 0771, 0780, 0767, 0766);
  lut lut_gate106(0x0, 0718, 0768, 1011, 0767);
  lut lut_gate107(0x40, 0705, 0741, 0695, 0768);
  lut lut_gate108(0x4, 0759, 0752, 0769);
  lut lut_gate109(0x4, 0749, 0743, 0770);
  lut lut_gate110(0xc5, 1016, 0779, 0772, 0771);
  lut lut_gate111(0x4, 0773, 0715, 0772);
  lut lut_gate112(0x0e, 0774, 0776, 0707, 0773);
  lut lut_gate113(0x8, G38, 0775, 0774);
  lut lut_gate114(0x0e, G1, G5, G6, 0775);
  lut lut_gate115(0x0, 0777, 0775, G33, 0776);
  lut lut_gate116(0x07, 0778, 0712, G31, 0777);
  lut lut_gate117(0xca, G4, G32, G13, 0778);
  lut lut_gate118(0x4, 0773, 0717, 0779);
  lut lut_gate119(0x4, 0718, 1016, 0780);
  lut lut_gate120(0x10, G4, G2, 0782, 0781);
  lut lut_gate121(0x9, 0780, 0771, 0782);
  lut lut_gate122(0x8, 0689, 1019, 0783);
  lut lut_gate123(0x4, G20, 1066, 0784);
  lut lut_gate124(0x1, G7, 1065, 0785);
  lut lut_gate125(0x10, 0789, 0788, 0787, 0786);
  lut lut_gate126(0x0b, 1058, G14, G42, 0787);
  lut lut_gate127(0x0, 1060, G39, G11, 0788);
  lut lut_gate128(0x0, G4, 1066, G40, 0789);
  lut lut_gate129(0x0, 0803, 0791, 0800, 0790);
  lut lut_gate130(0x4, 0767, 0792, 0791);
  lut lut_gate131(0x6, 0795, G3526, 0792);
  lut lut_gate132(0x40, G47, 0793, 0693, G3526);
  lut lut_gate133(0x9, 0794, 0742, 0793);
  lut lut_gate134(0x4, 0718, 0743, 0794);
  lut lut_gate135(0x1e, 0799, 0797, 0796, 0795);
  lut lut_gate136(0x4, 0770, 0718, 0796);
  lut lut_gate137(0x41, 0742, 0794, 0798, 0797);
  lut lut_gate138(0x10, 0705, 0718, 0695, 0798);
  lut lut_gate139(0x4b, 0751, 0718, 0752, 0799);
  lut lut_gate140(0x0b, 0690, 0767, 0801, 0800);
  lut lut_gate141(0x87, 0802, G47, 0693, 0801);
  lut lut_gate142(0x1e, 0742, 0798, 0794, 0802);
  lut lut_gate143(0x01, 0728, 0804, 0692, 0803);
  lut lut_gate144(0x4, G3, G1, 0804);
  lut lut_gate145(0xb4, 0761, 0718, 1009, 0805);
  lut lut_gate146(0x70, 0807, 0805, 0720, 0806);
  lut lut_gate147(0x8, 0689, 0808, 0807);
  lut lut_gate148(0x07, 0813, 0809, 0821, 0808);
  lut lut_gate149(0x40, G8, 0810, 0812, 0809);
  lut lut_gate150(0x0, 0811, 1057, G20, 0810);
  lut lut_gate151(0x4, G21, 1066, 0811);
  lut lut_gate152(0x0, 1060, G22, G10, 0812);
  lut lut_gate153(0x80, 0819, 0817, 0814, 0813);
  lut lut_gate154(0x10, G4, 0816, 0815, 0814);
  lut lut_gate155(0x0b, 1060, G12, G40, 0815);
  lut lut_gate156(0x0e, 1058, G39, G43, 0816);
  lut lut_gate157(0x0, 0818, 1066, G41, 0817);
  lut lut_gate158(0x1, G13, 1054, 0818);
  lut lut_gate159(0x0, 0820, 1057, G42, 0819);
  lut lut_gate160(0x1, G14, 1065, 0820);
  lut lut_gate161(0x01, G4, 0823, 0822, 0821);
  lut lut_gate162(0x1, G9, 1054, 0822);
  lut lut_gate163(0x0b, 1058, G7, G19, 0823);
  lut lut_gate164(0x4f, 0825, 0800, 0824, G3532);
  lut lut_gate165(0x4, 0801, 0767, 0824);
  lut lut_gate166(0x07, 0826, 0801, 0803, 0825);
  lut lut_gate167(0x0, 0827, 0793, 0720, 0826);
  lut lut_gate168(0x8, 0689, 0828, 0827);
  lut lut_gate169(0x07, 0835, 0829, 1023, 0828);
  lut lut_gate170(0x8, 0832, 0830, 0829);
  lut lut_gate171(0x0e, 0831, 1066, G7, 0830);
  lut lut_gate172(0x1, G11, 1054, 0831);
  lut lut_gate173(0x0, 0833, 1057, G22, 0832);
  lut lut_gate174(0x0b, 1058, G9, G21, 0833);
  lut lut_gate175(0x1, G10, 1065, 0834);
  lut lut_gate176(0x40, 0836, 0839, 0787, 0835);
  lut lut_gate177(0x10, G4, 0838, 0837, 0836);
  lut lut_gate178(0x4, G40, 1065, 0837);
  lut lut_gate179(0x0e, 1058, G41, G45, 0838);
  lut lut_gate180(0x0, 0840, 1057, G44, 0839);
  lut lut_gate181(0x4, G43, 1066, 0840);
  lut lut_gate182(0xb, 0842, 0841, G3533);
  lut lut_gate183(0x41, 0824, 0792, 0690, 0841);
  lut lut_gate184(0x07, 0843, 0792, 0803, 0842);
  lut lut_gate185(0x0, 0844, 0799, 0720, 0843);
  lut lut_gate186(0x8, 0689, 0845, 0844);
  lut lut_gate187(0x07, 0846, 0854, 0859, 0845);
  lut lut_gate188(0x40, 0847, 0852, G4, 0846);
  lut lut_gate189(0x10, 0848, 0851, 0850, 0847);
  lut lut_gate190(0x0e, 0849, 1065, G9, 0848);
  lut lut_gate191(0x1, G10, 1054, 0849);
  lut lut_gate192(0x0b, 1058, G8, G20, 0850);
  lut lut_gate193(0x07, 1060, G7, G11, 0851);
  lut lut_gate194(0x0, 0853, 1066, G22, 0852);
  lut lut_gate195(0x4, G21, 1057, 0853);
  lut lut_gate196(0x10, 0855, 0858, 0857, 0854);
  lut lut_gate197(0x0, 0856, 1066, G42, 0855);
  lut lut_gate198(0x0, 1060, G41, G13, 0856);
  lut lut_gate199(0x1, G14, 1054, 0857);
  lut lut_gate200(0x4, G43, 1057, 0858);
  lut lut_gate201(0x10, G4, 0861, 0860, 0859);
  lut lut_gate202(0x4, G39, 1065, 0860);
  lut lut_gate203(0x0e, 1058, G40, G44, 0861);
  lut lut_gate204(0x0e, 0910, 0863, 0803, 0862);
  lut lut_gate205(0x01, 0690, 0904, 0864, 0863);
  lut lut_gate206(0x40, G47, 0903, 0865, 0864);
  lut lut_gate207(0xe0, 0866, 0767, 0902, 0865);
  lut lut_gate208(0x70, 0898, 0867, 0901, 0866);
  lut lut_gate209(0x8, 0889, 0868, 0867);
  lut lut_gate210(0x8, 0879, 0869, 0868);
  lut lut_gate211(0xc5, 1029, 0878, 0873, 0869);
  lut lut_gate212(0xca, G8, 0871, 0701, 0870);
  lut lut_gate213(0x01, 0804, 0699, 0698, 0871);
  lut lut_gate214(0x6, G8, G9, 0872);
  lut lut_gate215(0x01, 0715, 0874, 0774, 0873);
  lut lut_gate216(0x0, 0707, 0875, 0876, 0874);
  lut lut_gate217(0x8, G29, 0712, 0875);
  lut lut_gate218(0x0, 0877, 0775, G31, 0876);
  lut lut_gate219(0x35, G4, G30, G11, 0877);
  lut lut_gate220(0x01, 0717, 0874, 0774, 0878);
  lut lut_gate221(0xc5, 1032, 0888, 0883, 0879);
  lut lut_gate222(0xb0, G3, 0881, G7, 0880);
  lut lut_gate223(0x1, G8, G9, 0881);
  lut lut_gate224(0xca, G7, 0871, 0701, 0882);
  lut lut_gate225(0x01, 0715, 0884, 0774, 0883);
  lut lut_gate226(0x0, 0707, 0885, 0886, 0884);
  lut lut_gate227(0x8, G28, 0712, 0885);
  lut lut_gate228(0x0, 0887, 0775, G30, 0886);
  lut lut_gate229(0xca, G4, G29, G10, 0887);
  lut lut_gate230(0x01, 0717, 0884, 0774, 0888);
  lut lut_gate231(0x0, 0890, 0897, 1035, 0889);
  lut lut_gate232(0x10, 0893, 0715, 1035, 0890);
  lut lut_gate233(0x8, G9, 0871, 0891);
  lut lut_gate234(0x10, G3, G9, 0746, 0892);
  lut lut_gate235(0x0e, 0774, 0894, 0707, 0893);
  lut lut_gate236(0x0, 0895, 0775, G32, 0894);
  lut lut_gate237(0x70, 0896, 0712, G30, 0895);
  lut lut_gate238(0x35, G4, G31, G12, 0896);
  lut lut_gate239(0x4, 0893, 0717, 0897);
  lut lut_gate240(0x70, 0899, 0868, 0890, 0898);
  lut lut_gate241(0x5c, 0879, 1032, 0900, 0899);
  lut lut_gate242(0x4, 0873, 1029, 0900);
  lut lut_gate243(0x4, 0772, 1016, 0901);
  lut lut_gate244(0x8, 0771, 0867, 0902);
  lut lut_gate245(0x4, 0724, 0902, 0903);
  lut lut_gate246(0x9, 0907, 0905, 0904);
  lut lut_gate247(0x0e, 0906, 0767, 0782, 0905);
  lut lut_gate248(0x4, 0901, 0718, 0906);
  lut lut_gate249(0x78, 0909, G47, 0908, 0907);
  lut lut_gate250(0x01, 0782, 0740, 1045, 0908);
  lut lut_gate251(0xb4, 0889, 0718, 1035, 0909);
  lut lut_gate252(0x69, 0913, 0912, 0911, 0910);
  lut lut_gate253(0x80, G47, 0909, 0908, 0911);
  lut lut_gate254(0xa3, 0909, 0890, 0906, 0912);
  lut lut_gate255(0x4b, 0869, 0914, 1029, 0913);
  lut lut_gate256(0x8, G27, 0691, 0914);
  lut lut_gate257(0x8, 0910, 0916, 0915);
  lut lut_gate258(0x0e, 0690, 0864, 0904, 0916);
  lut lut_gate259(0x80, 0921, 0918, 1063, 0917);
  lut lut_gate260(0x01, 0920, 0919, 0849, 0918);
  lut lut_gate261(0x1, G14, 1066, 0919);
  lut lut_gate262(0x4, G39, 1057, 0920);
  lut lut_gate263(0x10, G4, 0922, 1059, 0921);
  lut lut_gate264(0x0b, 1058, G12, G40, 0922);
  lut lut_gate265(0x0e, 1058, G20, G16, 0923);
  lut lut_gate266(0x0, 0925, 1057, G17, 0924);
  lut lut_gate267(0x4, G18, 1066, 0925);
  lut lut_gate268(0x01, 0929, 0928, 0927, 0926);
  lut lut_gate269(0x4, G22, 1054, 0927);
  lut lut_gate270(0x0b, 1060, G7, G19, 0928);
  lut lut_gate271(0x4, G21, 1065, 0929);
  lut lut_gate272(0xb, 1039, 0930, G3536);
  lut lut_gate273(0x14, 0904, 0864, 0690, 0930);
  lut lut_gate274(0x0e, 1058, G21, G17, 0931);
  lut lut_gate275(0x0, 0933, 1066, G19, 0932);
  lut lut_gate276(0x4, G18, 1057, 0933);
  lut lut_gate277(0x0, 0935, 1065, G22, 0934);
  lut lut_gate278(0x0b, 1060, G8, G20, 0935);
  lut lut_gate279(0x80, 0941, 0939, 0937, 0936);
  lut lut_gate280(0x10, G4, 0938, 0831, 0937);
  lut lut_gate281(0x0, 1058, G41, G13, 0938);
  lut lut_gate282(0x0, 0940, 1057, G40, 0939);
  lut lut_gate283(0x1, G12, 1065, 0940);
  lut lut_gate284(0x0, 0942, 1066, G39, 0941);
  lut lut_gate285(0x07, 1060, G14, G10, 0942);
  lut lut_gate286(0xf4, 1043, 0945, 0943, G3535);
  lut lut_gate287(0x0b, 0803, 0944, 0690, 0943);
  lut lut_gate288(0x1f, 0864, 0910, 0904, 0944);
  lut lut_gate289(0x96, 0949, 0948, 0946, 0945);
  lut lut_gate290(0x8, G47, 0947, 0946);
  lut lut_gate291(0x40, 0908, 0909, 0913, 0947);
  lut lut_gate292(0x5c, 0913, 0912, 0900, 0948);
  lut lut_gate293(0x4b, 0879, 0914, 1032, 0949);
  lut lut_gate294(0x40, 1023, 0951, 0788, 0950);
  lut lut_gate295(0x0e, 0952, 1066, G13, 0951);
  lut lut_gate296(0x1, G14, 1057, 0952);
  lut lut_gate297(0x4, G20, 1065, 0953);
  lut lut_gate298(0x0e, 1058, G19, G15, 0954);
  lut lut_gate299(0x0, 0956, 1057, G16, 0955);
  lut lut_gate300(0x0e, 1060, G22, G18, 0956);
  lut lut_gate301(0x0, 0958, 1066, G17, 0957);
  lut lut_gate302(0x4, G21, 1054, 0958);
  lut lut_gate303(0x4b, 0960, 0959, 0719, G3539);
  lut lut_gate304(0x96, G50, G3535, G3534, 0959);
  lut lut_gate305(0x96, G3529, 0961, G3536, 0960);
  lut lut_gate306(0x69, 0962, G3533, G3531, 0961);
  lut lut_gate307(0x6, G3528, G3532, 0962);
  lut lut_gate308(0x1f, G11, G13, G12, G3520);
  lut lut_gate309(0x70, 0963, 0975, 0976, G3521);
  lut lut_gate310(0x07, 0964, 0691, 0974, 0963);
  lut lut_gate311(0x0e, 0965, G1, G3, 0964);
  lut lut_gate312(0x80, 0972, 0969, 0966, 0965);
  lut lut_gate313(0x0, 0967, G14, G37, 0966);
  lut lut_gate314(0x0, 0968, G11, G34, 0967);
  lut lut_gate315(0x4, G31, G8, 0968);
  lut lut_gate316(0x0, 0970, G12, G35, 0969);
  lut lut_gate317(0x0, 0971, G9, G32, 0970);
  lut lut_gate318(0x4, G33, G10, 0971);
  lut lut_gate319(0x0b, 0973, G36, G13, 0972);
  lut lut_gate320(0x4, G30, G7, 0973);
  lut lut_gate321(0xe0, G34, G35, G36, 0974);
  lut lut_gate322(0x4, 0692, G3, 0975);
  lut lut_gate323(0x1, G7, 0881, 0976);
  lut lut_gate324(0x6, 0979, 0977, G3523);
  lut lut_gate325(0x69, G10, G9, 0978, 0977);
  lut lut_gate326(0x9, G8, G7, 0978);
  lut lut_gate327(0x96, G12, G14, 0980, 0979);
  lut lut_gate328(0x6, G13, G11, 0980);
  lut lut_gate329(0xb, 0866, 0981, G3525);
  lut lut_gate330(0x0, 0902, 0768, 1011, 0981);
  lut lut_gate331(0xef, 0982, G3535, G3534, G3537);
  lut lut_gate332(0x80, 0985, 0984, 0983, 0982);
  lut lut_gate333(0x10, 1039, 0930, G3529, 0983);
  lut lut_gate334(0x1, G3533, G3531, 0984);
  lut lut_gate335(0x1, G3528, G3532, 0985);
  lut lut_gate336(0xbf, G27, G3537, 0986, G3538);
  lut lut_gate337(0x10, G48, G3535, G3534, 0986);
  lut lut_gate338(0x10, 0881, G10, G7, G3519);
  lut lut_gate339(0x9, 0989, 0987, G3522);
  lut lut_gate340(0x96, G30, G31, 0988, 0987);
  lut lut_gate341(0x9, G33, G32, 0988);
  lut lut_gate342(0x69, G34, G36, 0990, 0989);
  lut lut_gate343(0x9, G35, G37, 0990);
  lut lut_gate344(0xf4, 0991, 0767, G1, G3527);
  lut lut_gate345(0x4, 0976, 0690, 0991);
  lut lut_gate346(0xb, 0992, 0998, G3530);
  lut lut_gate347(0x0, 0995, 0993, 0997, 0992);
  lut lut_gate348(0x69, 0948, 0865, 0994, 0993);
  lut lut_gate349(0x60, G47, 0947, 0903, 0994);
  lut lut_gate350(0x10, 0975, G14, 0996, 0995);
  lut lut_gate351(0x6, G13, G12, 0996);
  lut lut_gate352(0xf8, G1, G3, G2, 0997);
  lut lut_gate353(0x01, G1, G2, 0999, 0998);
  lut lut_gate354(0x0b, 1000, G7, G9, 0999);
  lut lut_gate355(0x01, G10, G7, 0872, 1000);
  lut lut_gate356(0x96, 0960, G3535, G3534, G3540);
  lut lut_gate357(0x80, 0694, 0741, 0902, G3524);
  lut lut_gate358(0xac, 0689, G47, 0720, 1001);
  lut lut_gate359(0x9e, 1001, 0693, 0689, 1002);
  lut lut_gate360(0x0, 1002, 1049, 0689, G3528);
  lut lut_gate361(0x2b, 0736, 0732, G24, 1003);
  lut lut_gate362(0xbc, 1003, G24, 0706, 1004);
  lut lut_gate363(0xca, G4, G12, G9, 1005);
  lut lut_gate364(0xca, G3, 0762, 1005, 1006);
  lut lut_gate365(0x0e, 0763, 1006, 0697, 1007);
  lut lut_gate366(0x8, 0700, G11, 1008);
  lut lut_gate367(0x70, 1007, 1008, 0697, 1009);
  lut lut_gate368(0x07, 0769, 0751, 0770, 1010);
  lut lut_gate369(0xca, 0761, 1010, 1009, 1011);
  lut lut_gate370(0xca, G4, G11, G8, 1012);
  lut lut_gate371(0x3a, G3, G1, 1012, 1013);
  lut lut_gate372(0x83, 0697, G3, G10, 1014);
  lut lut_gate373(0xc5, G10, 1014, 0701, 1015);
  lut lut_gate374(0x0, 1015, 1013, 1014, 1016);
  lut lut_gate375(0xb0, 0786, G41, 1057, 1017);
  lut lut_gate376(0xb0, 1048, G19, 1057, 1018);
  lut lut_gate377(0x35, 1017, G13, 1018, 1019);
  lut lut_gate378(0x4b, G3526, 0795, 0769, 1020);
  lut lut_gate379(0x87, 0805, 0799, 1020, 1021);
  lut lut_gate380(0xf4, 0806, 1021, 0790, G3531);
  lut lut_gate381(0xf8, 1060, G12, G8, 1022);
  lut lut_gate382(0x10, 1022, 0834, G4, 1023);
  lut lut_gate383(0x40, 0926, 0924, 0923, 1024);
  lut lut_gate384(0xc5, G4, 0913, 1024, 1025);
  lut lut_gate385(0xbf, 1025, 0689, 0917, 1026);
  lut lut_gate386(0xef, 1026, 0915, 0862, G3534);
  lut lut_gate387(0xc5, G4, G9, G22, 1027);
  lut lut_gate388(0xc5, G3, 0872, 1027, 1028);
  lut lut_gate389(0x0b, 0870, 1028, 0697, 1029);
  lut lut_gate390(0x3a, G4, G8, G21, 1030);
  lut lut_gate391(0xf4, 0880, 1030, G3, 1031);
  lut lut_gate392(0x0b, 0882, 1031, 0697, 1032);
  lut lut_gate393(0xca, G4, G10, G7, 1033);
  lut lut_gate394(0xef, 1033, 0697, G3, 1034);
  lut lut_gate395(0x10, 1034, 0892, 0891, 1035);
  lut lut_gate396(0x40, 0934, 0932, 0931, 1036);
  lut lut_gate397(0x35, G4, 0909, 1036, 1037);
  lut lut_gate398(0xbf, 1037, 0689, 0936, 1038);
  lut lut_gate399(0xb0, 1038, 0803, 0904, 1039);
  lut lut_gate400(0x10, G5, 0954, 0953, 1040);
  lut lut_gate401(0x7f, 0957, 0955, 1040, 1041);
  lut lut_gate402(0x8f, G4, 0949, 1041, 1042);
  lut lut_gate403(0x40, 1042, 0689, 0950, 1043);
  lut lut_gate404(0x18, 0725, 0726, G24, 1044);
  lut lut_gate405(0x40, 1004, 1044, 0718, 1045);
  lut lut_gate406(0xf4, 1060, G9, G21, 1046);
  lut lut_gate407(0x10, 1061, 0785, 0784, 1047);
  lut lut_gate408(0x40, 1047, 1046, G18, 1048);

endmodule
