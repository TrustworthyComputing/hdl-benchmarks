module c1355(G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  lut lut_gate1(0x9, G1, 279, G1324);
  lut lut_gate2(0x1000, 291, 280, 299, 298, 279);
  lut lut_gate3(0x4, 286, 281, 280);
  lut lut_gate4(0x9669, 285, 284, 283, 282, 281);
  lut lut_gate5(0x7887, G25, G29, G37, G41, 282);
  lut lut_gate6(0x9, G21, G17, 283);
  lut lut_gate7(0x9669, G7, G8, G6, G5, 284);
  lut lut_gate8(0x9669, G3, G4, G2, G1, 285);
  lut lut_gate9(0x9669, 290, 289, 288, 287, 286);
  lut lut_gate10(0x7887, G26, G30, G38, G41, 287);
  lut lut_gate11(0x9, G22, G18, 288);
  lut lut_gate12(0x9669, G15, G16, G14, G13, 289);
  lut lut_gate13(0x9669, G11, G12, G10, G9, 290);
  lut lut_gate14(0x1, 295, 292, 291);
  lut lut_gate15(0x9669, 294, 293, 289, 284, 292);
  lut lut_gate16(0x8, G40, G41, 293);
  lut lut_gate17(0x9669, G28, G32, G24, G20, 294);
  lut lut_gate18(0x9669, 297, 296, 290, 285, 295);
  lut lut_gate19(0x7887, G27, G31, G39, G41, 296);
  lut lut_gate20(0x9, G23, G19, 297);
  lut lut_gate21(0x6bbf, 238, 230, 299, 235, 298);
  lut lut_gate22(0x9669, 229, 302, 301, 300, 299);
  lut lut_gate23(0x7887, G9, G13, G33, G41, 300);
  lut lut_gate24(0x9, G1, G5, 301);
  lut lut_gate25(0x9669, G23, G24, G21, G22, 302);
  lut lut_gate26(0x9669, G19, G20, G17, G18, 229);
  lut lut_gate27(0x9669, 234, 233, 232, 231, 230);
  lut lut_gate28(0x7887, G14, G10, G34, G41, 231);
  lut lut_gate29(0x9, G6, G2, 232);
  lut lut_gate30(0x9669, G32, G31, G30, G29, 233);
  lut lut_gate31(0x9669, G28, G27, G26, G25, 234);
  lut lut_gate32(0x9669, 237, 236, 233, 302, 235);
  lut lut_gate33(0x8, G36, G41, 236);
  lut lut_gate34(0x9669, G16, G12, G8, G4, 237);
  lut lut_gate35(0x9669, 240, 239, 234, 229, 238);
  lut lut_gate36(0x7887, G15, G11, G35, G41, 239);
  lut lut_gate37(0x9, G7, G3, 240);
  lut lut_gate38(0x9, G2, 241, G1325);
  lut lut_gate39(0x1000, 291, 280, 230, 298, 241);
  lut lut_gate40(0x9, G3, 242, G1326);
  lut lut_gate41(0x1000, 291, 280, 238, 298, 242);
  lut lut_gate42(0x9, G4, 243, G1327);
  lut lut_gate43(0x4000, 235, 280, 291, 298, 243);
  lut lut_gate44(0x9, G5, 244, G1328);
  lut lut_gate45(0x1000, 280, 245, 299, 298, 244);
  lut lut_gate46(0x8, 295, 292, 245);
  lut lut_gate47(0x9, G6, 246, G1329);
  lut lut_gate48(0x1000, 280, 245, 230, 298, 246);
  lut lut_gate49(0x9, G7, 247, G1330);
  lut lut_gate50(0x1000, 280, 245, 238, 298, 247);
  lut lut_gate51(0x9, G8, 248, G1331);
  lut lut_gate52(0x4000, 235, 245, 280, 298, 248);
  lut lut_gate53(0x9, G9, 249, G1332);
  lut lut_gate54(0x1000, 291, 250, 299, 298, 249);
  lut lut_gate55(0x4, 281, 286, 250);
  lut lut_gate56(0x9, G10, 251, G1333);
  lut lut_gate57(0x1000, 291, 250, 230, 298, 251);
  lut lut_gate58(0x9, G11, 252, G1334);
  lut lut_gate59(0x1000, 291, 250, 238, 298, 252);
  lut lut_gate60(0x9, G12, 253, G1335);
  lut lut_gate61(0x4000, 235, 250, 291, 298, 253);
  lut lut_gate62(0x9, G13, 254, G1336);
  lut lut_gate63(0x1000, 245, 250, 299, 298, 254);
  lut lut_gate64(0x9, G14, 255, G1337);
  lut lut_gate65(0x1000, 245, 250, 230, 298, 255);
  lut lut_gate66(0x9, G15, 256, G1338);
  lut lut_gate67(0x1000, 245, 250, 238, 298, 256);
  lut lut_gate68(0x9, G16, 257, G1339);
  lut lut_gate69(0x4000, 235, 250, 245, 298, 257);
  lut lut_gate70(0x9, G17, 258, G1340);
  lut lut_gate71(0x1000, 260, 259, 281, 261, 258);
  lut lut_gate72(0x4, 230, 299, 259);
  lut lut_gate73(0x1, 238, 235, 260);
  lut lut_gate74(0x6bbf, 295, 286, 281, 292, 261);
  lut lut_gate75(0x9, G18, 262, G1341);
  lut lut_gate76(0x1000, 260, 259, 286, 261, 262);
  lut lut_gate77(0x9, G19, 263, G1342);
  lut lut_gate78(0x1000, 260, 259, 295, 261, 263);
  lut lut_gate79(0x9, G20, 264, G1343);
  lut lut_gate80(0x4000, 292, 259, 260, 261, 264);
  lut lut_gate81(0x9, G21, 265, G1344);
  lut lut_gate82(0x1000, 266, 259, 281, 261, 265);
  lut lut_gate83(0x8, 238, 235, 266);
  lut lut_gate84(0x9, G22, 267, G1345);
  lut lut_gate85(0x1000, 266, 259, 286, 261, 267);
  lut lut_gate86(0x9, G23, 268, G1346);
  lut lut_gate87(0x1000, 266, 259, 295, 261, 268);
  lut lut_gate88(0x9, G24, 269, G1347);
  lut lut_gate89(0x4000, 292, 259, 266, 261, 269);
  lut lut_gate90(0x9, G25, 270, G1348);
  lut lut_gate91(0x1000, 260, 271, 281, 261, 270);
  lut lut_gate92(0x4, 299, 230, 271);
  lut lut_gate93(0x9, G26, 272, G1349);
  lut lut_gate94(0x1000, 260, 271, 286, 261, 272);
  lut lut_gate95(0x9, G27, 273, G1350);
  lut lut_gate96(0x1000, 260, 271, 295, 261, 273);
  lut lut_gate97(0x9, G28, 274, G1351);
  lut lut_gate98(0x4000, 292, 271, 260, 261, 274);
  lut lut_gate99(0x9, G29, 275, G1352);
  lut lut_gate100(0x1000, 266, 271, 281, 261, 275);
  lut lut_gate101(0x9, G30, 276, G1353);
  lut lut_gate102(0x1000, 266, 271, 286, 261, 276);
  lut lut_gate103(0x9, G31, 277, G1354);
  lut lut_gate104(0x1000, 266, 271, 295, 261, 277);
  lut lut_gate105(0x9, G32, 278, G1355);
  lut lut_gate106(0x4000, 292, 271, 266, 261, 278);

endmodule
