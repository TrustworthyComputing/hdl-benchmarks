module c1355(G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  lut lut_gate1(0x4b, G1, 303, 325, G1324);
  lut lut_gate2(0x40, 260, 242, 304, 303);
  lut lut_gate3(0x1, 238, 305, 304);
  lut lut_gate4(0x60, 306, 233, 325, 305);
  lut lut_gate5(0x4, 316, 307, 306);
  lut lut_gate6(0x69, 314, 310, 308, 307);
  lut lut_gate7(0x96, G32, G31, 309, 308);
  lut lut_gate8(0x9, G30, G29, 309);
  lut lut_gate9(0x96, 313, 312, 311, 310);
  lut lut_gate10(0x6, G23, G24, 311);
  lut lut_gate11(0x9, G21, G22, 312);
  lut lut_gate12(0x8, G36, G41, 313);
  lut lut_gate13(0x96, G16, G12, 315, 314);
  lut lut_gate14(0x9, G8, G4, 315);
  lut lut_gate15(0x69, 321, 319, 317, 316);
  lut lut_gate16(0x96, G19, G20, 318, 317);
  lut lut_gate17(0x9, G17, G18, 318);
  lut lut_gate18(0x96, G28, G27, 320, 319);
  lut lut_gate19(0x9, G26, G25, 320);
  lut lut_gate20(0x96, 324, 323, 322, 321);
  lut lut_gate21(0x8, G35, G41, 322);
  lut lut_gate22(0x9, G15, G11, 323);
  lut lut_gate23(0x9, G7, G3, 324);
  lut lut_gate24(0x69, 317, 232, 326, 325);
  lut lut_gate25(0x96, 231, 230, 229, 326);
  lut lut_gate26(0x8, G33, G41, 229);
  lut lut_gate27(0x9, G9, G13, 230);
  lut lut_gate28(0x9, G1, G5, 231);
  lut lut_gate29(0x6, 312, 311, 232);
  lut lut_gate30(0x69, 319, 308, 234, 233);
  lut lut_gate31(0x96, 237, 236, 235, 234);
  lut lut_gate32(0x8, G34, G41, 235);
  lut lut_gate33(0x9, G14, G10, 236);
  lut lut_gate34(0x9, G6, G2, 237);
  lut lut_gate35(0xe0, 241, 239, 240, 238);
  lut lut_gate36(0x8, 316, 307, 239);
  lut lut_gate37(0x1, 316, 307, 240);
  lut lut_gate38(0x8, 233, 325, 241);
  lut lut_gate39(0x4, 252, 243, 242);
  lut lut_gate40(0x9, 247, 244, 243);
  lut lut_gate41(0x69, G21, G17, 245, 244);
  lut lut_gate42(0x78, 246, G37, G41, 245);
  lut lut_gate43(0x9, G25, G29, 246);
  lut lut_gate44(0x96, 251, 250, 248, 247);
  lut lut_gate45(0x96, G3, G4, 249, 248);
  lut lut_gate46(0x9, G2, G1, 249);
  lut lut_gate47(0x6, G7, G8, 250);
  lut lut_gate48(0x9, G6, G5, 251);
  lut lut_gate49(0x69, 258, 256, 253, 252);
  lut lut_gate50(0x69, G22, G18, 254, 253);
  lut lut_gate51(0x78, 255, G38, G41, 254);
  lut lut_gate52(0x9, G26, G30, 255);
  lut lut_gate53(0x96, G15, G16, 257, 256);
  lut lut_gate54(0x9, G14, G13, 257);
  lut lut_gate55(0x96, G11, G12, 259, 258);
  lut lut_gate56(0x9, G10, G9, 259);
  lut lut_gate57(0x1, 266, 261, 260);
  lut lut_gate58(0x69, 264, 262, 256, 261);
  lut lut_gate59(0x96, 263, 251, 250, 262);
  lut lut_gate60(0x8, G40, G41, 263);
  lut lut_gate61(0x96, G28, G32, 265, 264);
  lut lut_gate62(0x9, G24, G20, 265);
  lut lut_gate63(0x69, 267, 258, 248, 266);
  lut lut_gate64(0x96, 270, 269, 268, 267);
  lut lut_gate65(0x8, G39, G41, 268);
  lut lut_gate66(0x9, G27, G31, 269);
  lut lut_gate67(0x9, G23, G19, 270);
  lut lut_gate68(0x4b, G2, 303, 233, G1325);
  lut lut_gate69(0x4b, G3, 303, 316, G1326);
  lut lut_gate70(0x87, G4, 307, 303, G1327);
  lut lut_gate71(0x4b, G5, 271, 325, G1328);
  lut lut_gate72(0x8, 242, 272, 271);
  lut lut_gate73(0xe0, 273, 305, 238, 272);
  lut lut_gate74(0x8, 266, 261, 273);
  lut lut_gate75(0x4b, G6, 271, 233, G1329);
  lut lut_gate76(0x4b, G7, 271, 316, G1330);
  lut lut_gate77(0x9, G8, 274, G1331);
  lut lut_gate78(0x80, 307, 242, 272, 274);
  lut lut_gate79(0x4b, G9, 275, 325, G1332);
  lut lut_gate80(0x40, 260, 276, 304, 275);
  lut lut_gate81(0x4, 243, 252, 276);
  lut lut_gate82(0x4b, G10, 275, 233, G1333);
  lut lut_gate83(0x4b, G11, 275, 316, G1334);
  lut lut_gate84(0x87, G12, 307, 275, G1335);
  lut lut_gate85(0x4b, G13, 277, 325, G1336);
  lut lut_gate86(0x8, 276, 272, 277);
  lut lut_gate87(0x4b, G14, 277, 233, G1337);
  lut lut_gate88(0x4b, G15, 277, 316, G1338);
  lut lut_gate89(0x9, G16, 278, G1339);
  lut lut_gate90(0x80, 307, 276, 272, 278);
  lut lut_gate91(0x9, G17, 279, G1340);
  lut lut_gate92(0x40, 240, 280, 243, 279);
  lut lut_gate93(0xe0, 285, 281, 283, 280);
  lut lut_gate94(0x40, 243, 252, 282, 281);
  lut lut_gate95(0x6, 266, 261, 282);
  lut lut_gate96(0x60, 284, 252, 243, 283);
  lut lut_gate97(0x4, 266, 261, 284);
  lut lut_gate98(0x4, 233, 325, 285);
  lut lut_gate99(0x9, G18, 286, G1341);
  lut lut_gate100(0x40, 240, 280, 252, 286);
  lut lut_gate101(0x9, G19, 287, G1342);
  lut lut_gate102(0x40, 280, 240, 266, 287);
  lut lut_gate103(0x9, G20, 288, G1343);
  lut lut_gate104(0x80, 261, 240, 280, 288);
  lut lut_gate105(0x9, G21, 289, G1344);
  lut lut_gate106(0x40, 239, 280, 243, 289);
  lut lut_gate107(0x9, G22, 290, G1345);
  lut lut_gate108(0x40, 239, 280, 252, 290);
  lut lut_gate109(0x9, G23, 291, G1346);
  lut lut_gate110(0x40, 280, 239, 266, 291);
  lut lut_gate111(0x9, G24, 292, G1347);
  lut lut_gate112(0x80, 261, 239, 280, 292);
  lut lut_gate113(0x9, G25, 293, G1348);
  lut lut_gate114(0x40, 240, 294, 243, 293);
  lut lut_gate115(0xe0, 295, 281, 283, 294);
  lut lut_gate116(0x4, 325, 233, 295);
  lut lut_gate117(0x9, G26, 296, G1349);
  lut lut_gate118(0x40, 240, 294, 252, 296);
  lut lut_gate119(0x9, G27, 297, G1350);
  lut lut_gate120(0x40, 294, 240, 266, 297);
  lut lut_gate121(0x9, G28, 298, G1351);
  lut lut_gate122(0x80, 261, 240, 294, 298);
  lut lut_gate123(0x9, G29, 299, G1352);
  lut lut_gate124(0x40, 239, 294, 243, 299);
  lut lut_gate125(0x9, G30, 300, G1353);
  lut lut_gate126(0x40, 239, 294, 252, 300);
  lut lut_gate127(0x9, G31, 301, G1354);
  lut lut_gate128(0x40, 294, 239, 266, 301);
  lut lut_gate129(0x9, G32, 302, G1355);
  lut lut_gate130(0x80, 261, 239, 294, 302);

endmodule
