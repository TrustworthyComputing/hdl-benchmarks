module euclidean_distance (u_0, v_0, u_1, v_1, u_2, v_2, u_3, v_3, u_4, v_4, u_5, v_5, u_6, v_6, u_7, v_7, u_8, v_8, u_9, v_9, u_10, v_10, u_11, v_11, u_12, v_12, u_13, v_13, u_14, v_14, u_15, v_15, u_16, v_16, u_17, v_17, u_18, v_18, u_19, v_19, u_20, v_20, u_21, v_21, u_22, v_22, u_23, v_23, u_24, v_24, u_25, v_25, u_26, v_26, u_27, v_27, u_28, v_28, u_29, v_29, u_30, v_30, u_31, v_31, dist);

  input [15:0] u_0;
  input [15:0] v_0;
  input [15:0] u_1;
  input [15:0] v_1;
  input [15:0] u_2;
  input [15:0] v_2;
  input [15:0] u_3;
  input [15:0] v_3;
  input [15:0] u_4;
  input [15:0] v_4;
  input [15:0] u_5;
  input [15:0] v_5;
  input [15:0] u_6;
  input [15:0] v_6;
  input [15:0] u_7;
  input [15:0] v_7;
  input [15:0] u_8;
  input [15:0] v_8;
  input [15:0] u_9;
  input [15:0] v_9;
  input [15:0] u_10;
  input [15:0] v_10;
  input [15:0] u_11;
  input [15:0] v_11;
  input [15:0] u_12;
  input [15:0] v_12;
  input [15:0] u_13;
  input [15:0] v_13;
  input [15:0] u_14;
  input [15:0] v_14;
  input [15:0] u_15;
  input [15:0] v_15;
  input [15:0] u_16;
  input [15:0] v_16;
  input [15:0] u_17;
  input [15:0] v_17;
  input [15:0] u_18;
  input [15:0] v_18;
  input [15:0] u_19;
  input [15:0] v_19;
  input [15:0] u_20;
  input [15:0] v_20;
  input [15:0] u_21;
  input [15:0] v_21;
  input [15:0] u_22;
  input [15:0] v_22;
  input [15:0] u_23;
  input [15:0] v_23;
  input [15:0] u_24;
  input [15:0] v_24;
  input [15:0] u_25;
  input [15:0] v_25;
  input [15:0] u_26;
  input [15:0] v_26;
  input [15:0] u_27;
  input [15:0] v_27;
  input [15:0] u_28;
  input [15:0] v_28;
  input [15:0] u_29;
  input [15:0] v_29;
  input [15:0] u_30;
  input [15:0] v_30;
  input [15:0] u_31;
  input [15:0] v_31;

  output [15:0] dist;

  wire [15:0] t_diff_v0;
  wire [15:0] t0_sum_v0;
  wire [15:0] t_diff_v1;
  wire [15:0] t0_sum_v1;
  wire [15:0] t_diff_v2;
  wire [15:0] t0_sum_v2;
  wire [15:0] t_diff_v3;
  wire [15:0] t0_sum_v3;
  wire [15:0] t_diff_v4;
  wire [15:0] t0_sum_v4;
  wire [15:0] t_diff_v5;
  wire [15:0] t0_sum_v5;
  wire [15:0] t_diff_v6;
  wire [15:0] t0_sum_v6;
  wire [15:0] t_diff_v7;
  wire [15:0] t0_sum_v7;
  wire [15:0] t_diff_v8;
  wire [15:0] t0_sum_v8;
  wire [15:0] t_diff_v9;
  wire [15:0] t0_sum_v9;
  wire [15:0] t_diff_v10;
  wire [15:0] t0_sum_v10;
  wire [15:0] t_diff_v11;
  wire [15:0] t0_sum_v11;
  wire [15:0] t_diff_v12;
  wire [15:0] t0_sum_v12;
  wire [15:0] t_diff_v13;
  wire [15:0] t0_sum_v13;
  wire [15:0] t_diff_v14;
  wire [15:0] t0_sum_v14;
  wire [15:0] t_diff_v15;
  wire [15:0] t0_sum_v15;
  wire [15:0] t_diff_v16;
  wire [15:0] t0_sum_v16;
  wire [15:0] t_diff_v17;
  wire [15:0] t0_sum_v17;
  wire [15:0] t_diff_v18;
  wire [15:0] t0_sum_v18;
  wire [15:0] t_diff_v19;
  wire [15:0] t0_sum_v19;
  wire [15:0] t_diff_v20;
  wire [15:0] t0_sum_v20;
  wire [15:0] t_diff_v21;
  wire [15:0] t0_sum_v21;
  wire [15:0] t_diff_v22;
  wire [15:0] t0_sum_v22;
  wire [15:0] t_diff_v23;
  wire [15:0] t0_sum_v23;
  wire [15:0] t_diff_v24;
  wire [15:0] t0_sum_v24;
  wire [15:0] t_diff_v25;
  wire [15:0] t0_sum_v25;
  wire [15:0] t_diff_v26;
  wire [15:0] t0_sum_v26;
  wire [15:0] t_diff_v27;
  wire [15:0] t0_sum_v27;
  wire [15:0] t_diff_v28;
  wire [15:0] t0_sum_v28;
  wire [15:0] t_diff_v29;
  wire [15:0] t0_sum_v29;
  wire [15:0] t_diff_v30;
  wire [15:0] t0_sum_v30;
  wire [15:0] t_diff_v31;
  wire [15:0] t0_sum_v31;
  wire [15:0] t1_sum_v0;
  wire [15:0] t1_sum_v1;
  wire [15:0] t1_sum_v2;
  wire [15:0] t1_sum_v3;
  wire [15:0] t1_sum_v4;
  wire [15:0] t1_sum_v5;
  wire [15:0] t1_sum_v6;
  wire [15:0] t1_sum_v7;
  wire [15:0] t1_sum_v8;
  wire [15:0] t1_sum_v9;
  wire [15:0] t1_sum_v10;
  wire [15:0] t1_sum_v11;
  wire [15:0] t1_sum_v12;
  wire [15:0] t1_sum_v13;
  wire [15:0] t1_sum_v14;
  wire [15:0] t1_sum_v15;
  wire [15:0] t2_sum_v0;
  wire [15:0] t2_sum_v1;
  wire [15:0] t2_sum_v2;
  wire [15:0] t2_sum_v3;
  wire [15:0] t2_sum_v4;
  wire [15:0] t2_sum_v5;
  wire [15:0] t2_sum_v6;
  wire [15:0] t2_sum_v7;
  wire [15:0] t3_sum_v0;
  wire [15:0] t3_sum_v1;
  wire [15:0] t3_sum_v2;
  wire [15:0] t3_sum_v3;
  wire [15:0] t4_sum_v0;
  wire [15:0] t4_sum_v1;
  wire [15:0] t5_sum_v0;
  wire [15:0] t6_sum_v0;

  assign t_diff_v0 = v_0 - u_0;
  assign t0_sum_v0 = t_diff_v0 * t_diff_v0;
  assign t_diff_v1 = v_1 - u_1;
  assign t0_sum_v1 = t_diff_v1 * t_diff_v1;
  assign t_diff_v2 = v_2 - u_2;
  assign t0_sum_v2 = t_diff_v2 * t_diff_v2;
  assign t_diff_v3 = v_3 - u_3;
  assign t0_sum_v3 = t_diff_v3 * t_diff_v3;
  assign t_diff_v4 = v_4 - u_4;
  assign t0_sum_v4 = t_diff_v4 * t_diff_v4;
  assign t_diff_v5 = v_5 - u_5;
  assign t0_sum_v5 = t_diff_v5 * t_diff_v5;
  assign t_diff_v6 = v_6 - u_6;
  assign t0_sum_v6 = t_diff_v6 * t_diff_v6;
  assign t_diff_v7 = v_7 - u_7;
  assign t0_sum_v7 = t_diff_v7 * t_diff_v7;
  assign t_diff_v8 = v_8 - u_8;
  assign t0_sum_v8 = t_diff_v8 * t_diff_v8;
  assign t_diff_v9 = v_9 - u_9;
  assign t0_sum_v9 = t_diff_v9 * t_diff_v9;
  assign t_diff_v10 = v_10 - u_10;
  assign t0_sum_v10 = t_diff_v10 * t_diff_v10;
  assign t_diff_v11 = v_11 - u_11;
  assign t0_sum_v11 = t_diff_v11 * t_diff_v11;
  assign t_diff_v12 = v_12 - u_12;
  assign t0_sum_v12 = t_diff_v12 * t_diff_v12;
  assign t_diff_v13 = v_13 - u_13;
  assign t0_sum_v13 = t_diff_v13 * t_diff_v13;
  assign t_diff_v14 = v_14 - u_14;
  assign t0_sum_v14 = t_diff_v14 * t_diff_v14;
  assign t_diff_v15 = v_15 - u_15;
  assign t0_sum_v15 = t_diff_v15 * t_diff_v15;
  assign t_diff_v16 = v_16 - u_16;
  assign t0_sum_v16 = t_diff_v16 * t_diff_v16;
  assign t_diff_v17 = v_17 - u_17;
  assign t0_sum_v17 = t_diff_v17 * t_diff_v17;
  assign t_diff_v18 = v_18 - u_18;
  assign t0_sum_v18 = t_diff_v18 * t_diff_v18;
  assign t_diff_v19 = v_19 - u_19;
  assign t0_sum_v19 = t_diff_v19 * t_diff_v19;
  assign t_diff_v20 = v_20 - u_20;
  assign t0_sum_v20 = t_diff_v20 * t_diff_v20;
  assign t_diff_v21 = v_21 - u_21;
  assign t0_sum_v21 = t_diff_v21 * t_diff_v21;
  assign t_diff_v22 = v_22 - u_22;
  assign t0_sum_v22 = t_diff_v22 * t_diff_v22;
  assign t_diff_v23 = v_23 - u_23;
  assign t0_sum_v23 = t_diff_v23 * t_diff_v23;
  assign t_diff_v24 = v_24 - u_24;
  assign t0_sum_v24 = t_diff_v24 * t_diff_v24;
  assign t_diff_v25 = v_25 - u_25;
  assign t0_sum_v25 = t_diff_v25 * t_diff_v25;
  assign t_diff_v26 = v_26 - u_26;
  assign t0_sum_v26 = t_diff_v26 * t_diff_v26;
  assign t_diff_v27 = v_27 - u_27;
  assign t0_sum_v27 = t_diff_v27 * t_diff_v27;
  assign t_diff_v28 = v_28 - u_28;
  assign t0_sum_v28 = t_diff_v28 * t_diff_v28;
  assign t_diff_v29 = v_29 - u_29;
  assign t0_sum_v29 = t_diff_v29 * t_diff_v29;
  assign t_diff_v30 = v_30 - u_30;
  assign t0_sum_v30 = t_diff_v30 * t_diff_v30;
  assign t_diff_v31 = v_31 - u_31;
  assign t0_sum_v31 = t_diff_v31 * t_diff_v31;
  assign t1_sum_v0 = t0_sum_v0 + t0_sum_v1;
  assign t1_sum_v1 = t0_sum_v2 + t0_sum_v3;
  assign t1_sum_v2 = t0_sum_v4 + t0_sum_v5;
  assign t1_sum_v3 = t0_sum_v6 + t0_sum_v7;
  assign t1_sum_v4 = t0_sum_v8 + t0_sum_v9;
  assign t1_sum_v5 = t0_sum_v10 + t0_sum_v11;
  assign t1_sum_v6 = t0_sum_v12 + t0_sum_v13;
  assign t1_sum_v7 = t0_sum_v14 + t0_sum_v15;
  assign t1_sum_v8 = t0_sum_v16 + t0_sum_v17;
  assign t1_sum_v9 = t0_sum_v18 + t0_sum_v19;
  assign t1_sum_v10 = t0_sum_v20 + t0_sum_v21;
  assign t1_sum_v11 = t0_sum_v22 + t0_sum_v23;
  assign t1_sum_v12 = t0_sum_v24 + t0_sum_v25;
  assign t1_sum_v13 = t0_sum_v26 + t0_sum_v27;
  assign t1_sum_v14 = t0_sum_v28 + t0_sum_v29;
  assign t1_sum_v15 = t0_sum_v30 + t0_sum_v31;

  assign t2_sum_v0 = t1_sum_v0 + t1_sum_v1;
  assign t2_sum_v1 = t1_sum_v2 + t1_sum_v3;
  assign t2_sum_v2 = t1_sum_v4 + t1_sum_v5;
  assign t2_sum_v3 = t1_sum_v6 + t1_sum_v7;
  assign t2_sum_v4 = t1_sum_v8 + t1_sum_v9;
  assign t2_sum_v5 = t1_sum_v10 + t1_sum_v11;
  assign t2_sum_v6 = t1_sum_v12 + t1_sum_v13;
  assign t2_sum_v7 = t1_sum_v14 + t1_sum_v15;

  assign t3_sum_v0 = t2_sum_v0 + t2_sum_v1;
  assign t3_sum_v1 = t2_sum_v2 + t2_sum_v3;
  assign t3_sum_v2 = t2_sum_v4 + t2_sum_v5;
  assign t3_sum_v3 = t2_sum_v6 + t2_sum_v7;

  assign t4_sum_v0 = t3_sum_v0 + t3_sum_v1;
  assign t4_sum_v1 = t3_sum_v2 + t3_sum_v3;

  assign t5_sum_v0 = t4_sum_v0 + t4_sum_v1;

  assign t6_sum_v0 = t5_sum_v0;

  assign dist = t6_sum_v0;
endmodule
