module multiplier(G11, G12, G14);
  wire _0000_, _0001_, _0002_, _0003_, _0004_, _0005_, _0006_, _0007_, _0008_, _0009_, _0010_, _0011_, _0012_, _0013_, _0014_, _0015_, _0016_, _0017_, _0018_, _0019_, _0020_, _0021_, _0022_, _0023_, _0024_, _0025_, _0026_, _0027_, _0028_, _0029_, _0030_, _0031_, _0032_, _0033_, _0034_, _0035_, _0036_, _0037_, _0038_, _0039_, _0040_, _0041_, _0042_, _0043_, _0044_, _0045_, _0046_, _0047_, _0048_, _0049_, _0050_, _0051_, _0052_, _0053_, _0054_, _0055_, _0056_, _0057_, _0058_, _0059_, _0060_, _0061_, _0062_, _0063_, _0064_, _0065_, _0066_, _0067_, _0068_, _0069_, _0070_, _0071_, _0072_, _0073_, _0074_, _0075_, _0076_, _0077_, _0078_, _0079_, _0080_, _0081_, _0082_, _0083_, _0084_, _0085_, _0086_, _0087_, _0088_, _0089_, _0090_, _0091_, _0092_, _0093_, _0094_, _0095_, _0096_, _0097_, _0098_, _0099_, _0100_, _0101_, _0102_, _0103_, _0104_, _0105_, _0106_, _0107_, _0108_, _0109_, _0110_, _0111_, _0112_, _0113_, _0114_, _0115_, _0116_, _0117_, _0118_, _0119_, _0120_, _0121_, _0122_, _0123_, _0124_, _0125_, _0126_, _0127_, _0128_, _0129_, _0130_, _0131_, _0132_, _0133_, _0134_, _0135_, _0136_, _0137_, _0138_, _0139_, _0140_, _0141_, _0142_, _0143_, _0144_, _0145_, _0146_, _0147_, _0148_, _0149_, _0150_, _0151_, _0152_, _0153_, _0154_, _0155_, _0156_, _0157_, _0158_, _0159_, _0160_, _0161_, _0162_, _0163_, _0164_, _0165_, _0166_, _0167_, _0168_, _0169_, _0170_, _0171_, _0172_, _0173_, _0174_, _0175_, _0176_, _0177_, _0178_, _0179_, _0180_, _0181_, _0182_, _0183_, _0184_, _0185_, _0186_, _0187_, _0188_, _0189_, _0190_, _0191_, _0192_, _0193_, _0194_, _0195_, _0196_, _0197_, _0198_, _0199_, _0200_, _0201_, _0202_, _0203_, _0204_, _0205_, _0206_, _0207_, _0208_, _0209_, _0210_, _0211_, _0212_, _0213_, _0214_, _0215_, _0216_, _0217_, _0218_, _0219_, _0220_, _0221_, _0222_, _0223_, _0224_, _0225_, _0226_, _0227_, _0228_, _0229_, _0230_, _0231_, _0232_, _0233_, _0234_, _0235_, _0236_, _0237_, _0238_, _0239_, _0240_, _0241_, _0242_, _0243_, _0244_, _0245_, _0246_, _0247_, _0248_, _0249_, _0250_, _0251_, _0252_, _0253_, _0254_, _0255_, _0256_, _0257_, _0258_, _0259_, _0260_, _0261_, _0262_, _0263_, _0264_, _0265_, _0266_, _0267_, _0268_, _0269_, _0270_, _0271_, _0272_, _0273_, _0274_, _0275_, _0276_, _0277_, _0278_, _0279_, _0280_, _0281_, _0282_, _0283_, _0284_, _0285_, _0286_, _0287_, _0288_, _0289_, _0290_, _0291_, _0292_, _0293_, _0294_, _0295_, _0296_, _0297_, _0298_, _0299_, _0300_, _0301_, _0302_, _0303_, _0304_, _0305_, _0306_, _0307_, _0308_, _0309_, _0310_, _0311_, _0312_, _0313_, _0314_, _0315_, _0316_, _0317_, _0318_, _0319_, _0320_, _0321_, _0322_, _0323_, _0324_, _0325_, _0326_, _0327_, _0328_, _0329_, _0330_, _0331_, _0332_, _0333_, _0334_, _0335_, _0336_, _0337_, _0338_, _0339_, _0340_, _0341_, _0342_, _0343_, _0344_, _0345_, _0346_, _0347_, _0348_, _0349_, _0350_, _0351_, _0352_, _0353_, _0354_, _0355_, _0356_, _0357_, _0358_, _0359_, _0360_, _0361_, _0362_, _0363_, _0364_, _0365_, _0366_, _0367_, _0368_, _0369_, _0370_, _0371_, _0372_, _0373_, _0374_, _0375_, _0376_, _0377_, _0378_, _0379_, _0380_, _0381_, _0382_, _0383_, _0384_, _0385_, _0386_, _0387_, _0388_, _0389_, _0390_, _0391_, _0392_, _0393_, _0394_, _0395_, _0396_, _0397_, _0398_, _0399_, _0400_, _0401_, _0402_, _0403_, _0404_, _0405_, _0406_, _0407_, _0408_, _0409_, _0410_, _0411_, _0412_, _0413_, _0414_, _0415_, _0416_, _0417_, _0418_, _0419_, _0420_, _0421_, _0422_, _0423_, _0424_, _0425_, _0426_, _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0433_, _0434_, _0435_, _0436_, _0437_, _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_, _0446_, _0447_, _0448_, _0449_, _0450_, _0451_, _0452_, _0453_, _0454_, _0455_, _0456_, _0457_, _0458_, _0459_, _0460_, _0461_, _0462_, _0463_, _0464_, _0465_, _0466_, _0467_, _0468_, _0469_, _0470_, _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_, _0479_, _0480_, _0481_, _0482_, _0483_, _0484_, _0485_, _0486_, _0487_, _0488_, _0489_, _0490_, _0491_, _0492_, _0493_, _0494_, _0495_, _0496_, _0497_, _0498_, _0499_, _0500_, _0501_, _0502_, _0503_, _0504_, _0505_, _0506_, _0507_, _0508_, _0509_, _0510_, _0511_, _0512_, _0513_, _0514_, _0515_, _0516_, _0517_, _0518_, _0519_, _0520_, _0521_, _0522_, _0523_, _0524_, _0525_, _0526_, _0527_, _0528_, _0529_, _0530_, _0531_, _0532_, _0533_, _0534_, _0535_, _0536_, _0537_, _0538_, _0539_, _0540_, _0541_, _0542_, _0543_, _0544_, _0545_, _0546_, _0547_, _0548_, _0549_, _0550_, _0551_, _0552_, _0553_, _0554_, _0555_, _0556_, _0557_, _0558_, _0559_, _0560_, _0561_, _0562_, _0563_, _0564_, _0565_, _0566_, _0567_, _0568_, _0569_, _0570_, _0571_, _0572_, _0573_, _0574_, _0575_, _0576_, _0577_, _0578_, _0579_, _0580_, _0581_, _0582_, _0583_, _0584_, _0585_, _0586_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_, _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0602_, _0603_, _0604_, _0605_, _0606_, _0607_, _0608_, _0609_, _0610_, _0611_, _0612_, _0613_, _0614_, _0615_, _0616_, _0617_, _0618_, _0619_, _0620_, _0621_, _0622_, _0623_, _0624_, _0625_, _0626_, _0627_, _0628_, _0629_, _0630_, _0631_, _0632_, _0633_, _0634_, _0635_, _0636_, _0637_, _0638_, _0639_, _0640_, _0641_, _0642_, _0643_, _0644_, _0645_, _0646_, _0647_, _0648_, _0649_, _0650_, _0651_, _0652_, _0653_, _0654_, _0655_, _0656_, _0657_, _0658_, _0659_, _0660_, _0661_, _0662_, _0663_, _0664_, _0665_, _0666_, _0667_, _0668_, _0669_, _0670_, _0671_, _0672_, _0673_, _0674_, _0675_, _0676_, _0677_, _0678_, _0679_, _0680_, _0681_, _0682_, _0683_, _0684_, _0685_, _0686_, _0687_, _0688_, _0689_, _0690_, _0691_, _0692_, _0693_, _0694_, _0695_, _0696_, _0697_, _0698_, _0699_, _0700_, _0701_, _0702_, _0703_, _0704_, _0705_, _0706_, _0707_, _0708_, _0709_, _0710_, _0711_, _0712_, _0713_, _0714_, _0715_, _0716_, _0717_, _0718_, _0719_, _0720_, _0721_, _0722_, _0723_, _0724_, _0725_, _0726_, _0727_, _0728_, _0729_, _0730_, _0731_, _0732_, _0733_, _0734_, _0735_, _0736_, _0737_, _0738_, _0739_, _0740_, _0741_, _0742_, _0743_, _0744_, _0745_, _0746_, _0747_, _0748_, _0749_, _0750_, _0751_, _0752_, _0753_, _0754_, _0755_, _0756_, _0757_, _0758_, _0759_, _0760_, _0761_, _0762_, _0763_, _0764_, _0765_, _0766_, _0767_, _0768_, _0769_, _0770_, _0771_, _0772_, _0773_, _0774_, _0775_, _0776_, _0777_, _0778_, _0779_, _0780_, _0781_, _0782_, _0783_, _0784_, _0785_, _0786_, _0787_, _0788_, _0789_, _0790_, _0791_, _0792_, _0793_, _0794_, _0795_, _0796_, _0797_, _0798_, _0799_, _0800_, _0801_, _0802_, _0803_, _0804_, _0805_, _0806_, _0807_, _0808_, _0809_, _0810_, _0811_, _0812_, _0813_, _0814_, _0815_, _0816_, _0817_, _0818_, _0819_, _0820_, _0821_, _0822_, _0823_, _0824_, _0825_, _0826_, _0827_, _0828_, _0829_, _0830_, _0831_, _0832_, _0833_, _0834_, _0835_, _0836_, _0837_, _0838_, _0839_, _0840_, _0841_, _0842_, _0843_, _0844_, _0845_, _0846_, _0847_, _0848_, _0849_, _0850_, _0851_, _0852_, _0853_, _0854_, _0855_, _0856_, _0857_, _0858_, _0859_, _0860_, _0861_, _0862_, _0863_, _0864_, _0865_, _0866_, _0867_, _0868_, _0869_, _0870_, _0871_, _0872_, _0873_, _0874_, _0875_, _0876_, _0877_, _0878_, _0879_, _0880_, _0881_, _0882_, _0883_, _0884_, _0885_, _0886_, _0887_, _0888_, _0889_, _0890_, _0891_, _0892_, _0893_, _0894_, _0895_, _0896_, _0897_, _0898_, _0899_, _0900_, _0901_, _0902_, _0903_, _0904_, _0905_, _0906_, _0907_, _0908_, _0909_, _0910_, _0911_, _0912_, _0913_, _0914_, _0915_, _0916_, _0917_, _0918_, _0919_, _0920_, _0921_, _0922_, _0923_, _0924_, _0925_, _0926_, _0927_, _0928_, _0929_, _0930_, _0931_, _0932_, _0933_, _0934_, _0935_, _0936_, _0937_, _0938_, _0939_, _0940_, _0941_, _0942_, _0943_, _0944_, _0945_, _0946_, _0947_, _0948_, _0949_, _0950_, _0951_, _0952_, _0953_, _0954_, _0955_, _0956_, _0957_, _0958_, _0959_, _0960_, _0961_, _0962_, _0963_, _0964_, _0965_, _0966_, _0967_, _0968_, _0969_, _0970_, _0971_, _0972_, _0973_, _0974_, _0975_, _0976_, _0977_, _0978_, _0979_, _0980_, _0981_, _0982_, _0983_, _0984_, _0985_, _0986_, _0987_, _0988_, _0989_, _0990_, _0991_, _0992_, _0993_, _0994_, _0995_, _0996_, _0997_, _0998_, _0999_, _1000_, _1001_, _1002_, _1003_, _1004_, _1005_, _1006_, _1007_, _1008_, _1009_, _1010_, _1011_, _1012_, _1013_, _1014_, _1015_, _1016_, _1017_, _1018_, _1019_, _1020_, _1021_, _1022_, _1023_, _1024_, _1025_, _1026_, _1027_, _1028_, _1029_, _1030_, _1031_, _1032_, _1033_, _1034_, _1035_, _1036_, _1037_, _1038_, _1039_, _1040_, _1041_, _1042_, _1043_, _1044_, _1045_, _1046_, _1047_, _1048_, _1049_, _1050_, _1051_, _1052_, _1053_, _1054_, _1055_, _1056_, _1057_, _1058_, _1059_, _1060_, _1061_, _1062_, _1063_, _1064_, _1065_, _1066_, _1067_, _1068_, _1069_, _1070_, _1071_, _1072_, _1073_, _1074_, _1075_, _1076_, _1077_, _1078_, _1079_, _1080_, _1081_, _1082_, _1083_, _1084_, _1085_, _1086_, _1087_, _1088_, _1089_, _1090_, _1091_, _1092_, _1093_, _1094_, _1095_, _1096_, _1097_, _1098_, _1099_, _1100_, _1101_, _1102_, _1103_, _1104_, _1105_, _1106_, _1107_, _1108_, _1109_, _1110_, _1111_, _1112_, _1113_, _1114_, _1115_, _1116_, _1117_, _1118_, _1119_, _1120_, _1121_, _1122_, _1123_, _1124_, _1125_, _1126_, _1127_, _1128_, _1129_, _1130_, _1131_, _1132_, _1133_, _1134_, _1135_, _1136_, _1137_, _1138_, _1139_, _1140_, _1141_, _1142_, _1143_, _1144_, _1145_, _1146_, _1147_, _1148_, _1149_, _1150_, _1151_, _1152_, _1153_, _1154_, _1155_, _1156_, _1157_, _1158_, _1159_, _1160_, _1161_, _1162_, _1163_, _1164_, _1165_, _1166_, _1167_, _1168_, _1169_, _1170_, _1171_, _1172_, _1173_, _1174_, _1175_, _1176_, _1177_, _1178_, _1179_, _1180_, _1181_, _1182_, _1183_, _1184_, _1185_, _1186_, _1187_, _1188_, _1189_, _1190_, _1191_, _1192_, _1193_, _1194_, _1195_, _1196_, _1197_, _1198_, _1199_, _1200_, _1201_, _1202_, _1203_, _1204_, _1205_, _1206_, _1207_, _1208_, _1209_, _1210_, _1211_, _1212_, _1213_, _1214_, _1215_, _1216_, _1217_, _1218_, _1219_, _1220_, _1221_, _1222_, _1223_, _1224_, _1225_, _1226_, _1227_, _1228_, _1229_, _1230_, _1231_, _1232_, _1233_, _1234_, _1235_, _1236_, _1237_, _1238_, _1239_, _1240_, _1241_, _1242_, _1243_, _1244_, _1245_, _1246_, _1247_, _1248_, _1249_, _1250_, _1251_, _1252_, _1253_, _1254_, _1255_, _1256_, _1257_, _1258_, _1259_, _1260_, _1261_, _1262_, _1263_, _1264_, _1265_, _1266_, _1267_, _1268_, _1269_, _1270_, _1271_, _1272_, _1273_, _1274_, _1275_, _1276_, _1277_, _1278_, _1279_, _1280_, _1281_, _1282_, _1283_, _1284_, _1285_, _1286_, _1287_, _1288_, _1289_, _1290_, _1291_, _1292_, _1293_, _1294_, _1295_, _1296_, _1297_, _1298_, _1299_, _1300_, _1301_, _1302_, _1303_, _1304_, _1305_, _1306_, _1307_, _1308_, _1309_, _1310_, _1311_, _1312_, _1313_, _1314_, _1315_, _1316_, _1317_, _1318_, _1319_, _1320_, _1321_, _1322_, _1323_, _1324_, _1325_, _1326_, _1327_, _1328_, _1329_, _1330_, _1331_, _1332_, _1333_, _1334_, _1335_, _1336_, _1337_;
  input [15:0] G11;
  input [15:0] G12;
  input G11[0], G11[1], G11[2], G11[3], G11[4], G11[5], G11[6], G11[7], G11[8], G11[9], G11[10], G11[11], G11[12], G11[13], G11[14], G11[15], G12[0], G12[1], G12[2], G12[3], G12[4], G12[5], G12[6], G12[7], G12[8], G12[9], G12[10], G12[11], G12[12], G12[13], G12[14], G12[15];
  output G14[0], G14[1], G14[2], G14[3], G14[4], G14[5], G14[6], G14[7], G14[8], G14[9], G14[10], G14[11], G14[12], G14[13], G14[14], G14[15];
  and g_1338_(G12[0], G11[2], _1060_);
  and g_1339_(G12[1], G11[1], _1071_);
  and g_1340_(G12[0], G11[1], _1081_);
  not g_1341_(_1081_, _1092_);
  and g_1342_(G12[1], G11[2], _1103_);
  and g_1343_(_1081_, _1103_, _1114_);
  xor g_1344_(_1060_, _1071_, _1125_);
  and g_1345_(G11[0], G12[1], _1136_);
  and g_1346_(G11[0], G12[0], G14[0]);
  and g_1347_(_1071_, G14[0], _1157_);
  and g_1348_(_1125_, _1157_, _1167_);
  and g_1349_(G11[0], G12[2], _1178_);
  xor g_1350_(_1125_, _1157_, _1189_);
  and g_1351_(_1178_, _1189_, _1200_);
  or g_1352_(_1167_, _1200_, _1211_);
  and g_1353_(G11[1], G12[2], _1222_);
  and g_1354_(G11[3], G12[0], _1233_);
  and g_1355_(G12[3], G11[0], _1244_);
  and g_1356_(G12[3], G11[3], _1254_);
  and g_1357_(G14[0], _1254_, _1265_);
  not g_1358_(_1265_, _1276_);
  or g_1359_(_1233_, _1244_, _1287_);
  not g_1360_(_1287_, _1298_);
  and g_1361_(_1276_, _1287_, _1309_);
  or g_1362_(_1265_, _1298_, _1312_);
  and g_1363_(_1092_, _1103_, _1313_);
  xor g_1364_(_1309_, _1313_, _1314_);
  and g_1365_(_1222_, _1314_, _1315_);
  xor g_1366_(_1222_, _1314_, _1316_);
  and g_1367_(_1211_, _1316_, _1317_);
  xor g_1368_(_1211_, _1316_, G14[3]);
  and g_1369_(_1114_, _1312_, _1318_);
  or g_1370_(_1315_, _1318_, _1319_);
  and g_1371_(G11[0], G12[4], _1320_);
  and g_1372_(G11[2], G12[2], _1321_);
  and g_1373_(G11[2], G12[4], _1322_);
  and g_1374_(_1178_, _1322_, _1323_);
  xor g_1375_(_1320_, _1321_, _1324_);
  and g_1376_(G11[3], G12[1], _1325_);
  and g_1377_(G12[0], G11[4], _1326_);
  and g_1378_(G12[3], G11[1], _1327_);
  and g_1379_(G12[3], G11[4], _1328_);
  and g_1380_(_1081_, _1328_, _1329_);
  xor g_1381_(_1326_, _1327_, _1330_);
  and g_1382_(_1325_, _1330_, _1331_);
  xor g_1383_(_1325_, _1330_, _1332_);
  and g_1384_(_1103_, _1287_, _1333_);
  or g_1385_(_1265_, _1333_, _1334_);
  and g_1386_(_1332_, _1334_, _1335_);
  xor g_1387_(_1332_, _1334_, _1336_);
  and g_1388_(_1324_, _1336_, _1337_);
  xor g_1389_(_1324_, _1336_, _0667_);
  and g_1390_(_1319_, _0667_, _0668_);
  xor g_1391_(_1319_, _0667_, _0669_);
  and g_1392_(_1317_, _0669_, _0670_);
  xor g_1393_(_1317_, _0669_, G14[4]);
  or g_1394_(_1335_, _1337_, _0671_);
  and g_1395_(G11[0], G12[5], _0672_);
  and g_1396_(G11[1], G12[4], _0673_);
  and g_1397_(G11[3], G12[2], _0674_);
  and g_1398_(G11[3], G12[4], _0675_);
  and g_1399_(_1222_, _0675_, _0676_);
  xor g_1400_(_0673_, _0674_, _0677_);
  and g_1401_(_0672_, _0677_, _0678_);
  xor g_1402_(_0672_, _0677_, _0679_);
  or g_1403_(_1329_, _1331_, _0680_);
  and g_1404_(G12[1], G11[4], _0681_);
  and g_1405_(G12[0], G11[5], _0682_);
  and g_1406_(G12[3], G11[2], _0683_);
  and g_1407_(G12[3], G11[5], _0684_);
  and g_1408_(_1060_, _0684_, _0685_);
  xor g_1409_(_0682_, _0683_, _0686_);
  and g_1410_(_0681_, _0686_, _0687_);
  xor g_1411_(_0681_, _0686_, _0688_);
  and g_1412_(_0680_, _0688_, _0689_);
  xor g_1413_(_0680_, _0688_, _0690_);
  and g_1414_(_0679_, _0690_, _0691_);
  xor g_1415_(_0679_, _0690_, _0692_);
  and g_1416_(_0671_, _0692_, _0693_);
  xor g_1417_(_0671_, _0692_, _0694_);
  and g_1418_(_1323_, _0694_, _0695_);
  xor g_1419_(_1323_, _0694_, _0696_);
  and g_1420_(_0668_, _0696_, _0697_);
  xor g_1421_(_0668_, _0696_, _0698_);
  and g_1422_(_0670_, _0698_, _0699_);
  xor g_1423_(_0670_, _0698_, G14[5]);
  or g_1424_(_0693_, _0695_, _0700_);
  and g_1425_(G11[0], G12[6], _0701_);
  or g_1426_(_0676_, _0678_, _0702_);
  and g_1427_(_0701_, _0702_, _0703_);
  xor g_1428_(_0701_, _0702_, _0704_);
  or g_1429_(_0689_, _0691_, _0705_);
  and g_1430_(G11[1], G12[5], _0706_);
  and g_1431_(G12[2], G11[4], _0707_);
  and g_1432_(G11[4], G12[4], _0708_);
  and g_1433_(_1322_, _0707_, _0709_);
  xor g_1434_(_1322_, _0707_, _0710_);
  and g_1435_(_0706_, _0710_, _0711_);
  xor g_1436_(_0706_, _0710_, _0712_);
  or g_1437_(_0685_, _0687_, _0713_);
  and g_1438_(G12[1], G11[5], _0714_);
  and g_1439_(G12[0], G11[6], _0715_);
  and g_1440_(G12[3], G11[6], _0716_);
  and g_1441_(_1254_, _0715_, _0717_);
  xor g_1442_(_1254_, _0715_, _0718_);
  and g_1443_(_0714_, _0718_, _0719_);
  xor g_1444_(_0714_, _0718_, _0720_);
  and g_1445_(_0713_, _0720_, _0721_);
  xor g_1446_(_0713_, _0720_, _0722_);
  and g_1447_(_0712_, _0722_, _0723_);
  xor g_1448_(_0712_, _0722_, _0724_);
  and g_1449_(_0705_, _0724_, _0725_);
  xor g_1450_(_0705_, _0724_, _0726_);
  and g_1451_(_0704_, _0726_, _0727_);
  xor g_1452_(_0704_, _0726_, _0728_);
  and g_1453_(_0700_, _0728_, _0729_);
  xor g_1454_(_0700_, _0728_, _0730_);
  and g_1455_(_0697_, _0730_, _0731_);
  xor g_1456_(_0697_, _0730_, _0732_);
  and g_1457_(_0699_, _0732_, _0733_);
  xor g_1458_(_0699_, _0732_, G14[6]);
  or g_1459_(_0725_, _0727_, _0734_);
  or g_1460_(_0721_, _0723_, _0735_);
  or g_1461_(_0717_, _0719_, _0736_);
  and g_1462_(G12[1], G11[6], _0737_);
  and g_1463_(G12[0], G11[7], _0738_);
  and g_1464_(G12[3], G11[7], _0739_);
  and g_1465_(_1328_, _0738_, _0740_);
  xor g_1466_(_1328_, _0738_, _0741_);
  and g_1467_(_0737_, _0741_, _0742_);
  xor g_1468_(_0737_, _0741_, _0743_);
  and g_1469_(_0736_, _0743_, _0744_);
  xor g_1470_(_0736_, _0743_, _0745_);
  and g_1471_(G11[2], G12[5], _0746_);
  and g_1472_(G12[2], G11[5], _0747_);
  and g_1473_(G12[4], G11[5], _0748_);
  and g_1474_(_0675_, _0747_, _0749_);
  xor g_1475_(_0675_, _0747_, _0750_);
  and g_1476_(_0746_, _0750_, _0751_);
  xor g_1477_(_0746_, _0750_, _0752_);
  and g_1478_(_0745_, _0752_, _0753_);
  xor g_1479_(_0745_, _0752_, _0754_);
  and g_1480_(_0735_, _0754_, _0755_);
  xor g_1481_(_0735_, _0754_, _0756_);
  and g_1482_(G11[0], G12[7], _0757_);
  and g_1483_(G11[1], G12[6], _0758_);
  and g_1484_(G11[1], G12[7], _0759_);
  and g_1485_(_0701_, _0759_, _0760_);
  xor g_1486_(_0757_, _0758_, _0761_);
  or g_1487_(_0709_, _0711_, _0762_);
  and g_1488_(_0761_, _0762_, _0763_);
  xor g_1489_(_0761_, _0762_, _0764_);
  and g_1490_(_0756_, _0764_, _0765_);
  xor g_1491_(_0756_, _0764_, _0766_);
  and g_1492_(_0734_, _0766_, _0767_);
  xor g_1493_(_0734_, _0766_, _0768_);
  and g_1494_(_0703_, _0768_, _0769_);
  xor g_1495_(_0703_, _0768_, _0770_);
  and g_1496_(_0729_, _0770_, _0771_);
  xor g_1497_(_0729_, _0770_, _0772_);
  and g_1498_(_0733_, _0772_, _0773_);
  and g_1499_(_0731_, _0772_, _0774_);
  or g_1500_(_0767_, _0769_, _0775_);
  or g_1501_(_0755_, _0765_, _0776_);
  and g_1502_(G11[0], G12[8], _0777_);
  and g_1503_(G11[2], G12[6], _0778_);
  and g_1504_(G11[2], G12[7], _0779_);
  and g_1505_(_0759_, _0778_, _0780_);
  xor g_1506_(_0759_, _0778_, _0781_);
  and g_1507_(_0777_, _0781_, _0782_);
  xor g_1508_(_0777_, _0781_, _0783_);
  or g_1509_(_0749_, _0751_, _0784_);
  and g_1510_(_0783_, _0784_, _0785_);
  xor g_1511_(_0783_, _0784_, _0786_);
  and g_1512_(_0760_, _0786_, _0787_);
  xor g_1513_(_0760_, _0786_, _0788_);
  or g_1514_(_0744_, _0753_, _0789_);
  and g_1515_(G11[3], G12[5], _0790_);
  and g_1516_(G12[2], G11[6], _0791_);
  and g_1517_(G12[4], G11[6], _0792_);
  and g_1518_(_0708_, _0791_, _0793_);
  xor g_1519_(_0708_, _0791_, _0794_);
  and g_1520_(_0790_, _0794_, _0795_);
  xor g_1521_(_0790_, _0794_, _0796_);
  or g_1522_(_0740_, _0742_, _0797_);
  and g_1523_(G12[1], G11[7], _0798_);
  and g_1524_(G12[0], G11[8], _0799_);
  and g_1525_(G12[3], G11[8], _0800_);
  and g_1526_(_0684_, _0799_, _0801_);
  xor g_1527_(_0684_, _0799_, _0802_);
  and g_1528_(_0798_, _0802_, _0803_);
  xor g_1529_(_0798_, _0802_, _0804_);
  and g_1530_(_0797_, _0804_, _0805_);
  xor g_1531_(_0797_, _0804_, _0806_);
  and g_1532_(_0796_, _0806_, _0807_);
  xor g_1533_(_0796_, _0806_, _0808_);
  and g_1534_(_0789_, _0808_, _0809_);
  xor g_1535_(_0789_, _0808_, _0810_);
  and g_1536_(_0788_, _0810_, _0811_);
  xor g_1537_(_0788_, _0810_, _0812_);
  and g_1538_(_0776_, _0812_, _0813_);
  xor g_1539_(_0776_, _0812_, _0814_);
  and g_1540_(_0763_, _0814_, _0815_);
  xor g_1541_(_0763_, _0814_, _0816_);
  and g_1542_(_0775_, _0816_, _0817_);
  xor g_1543_(_0775_, _0816_, _0818_);
  and g_1544_(_0771_, _0818_, _0819_);
  xor g_1545_(_0771_, _0818_, _0820_);
  and g_1546_(_0774_, _0820_, _0821_);
  xor g_1547_(_0774_, _0820_, _0822_);
  and g_1548_(_0773_, _0822_, _0823_);
  xor g_1549_(_0773_, _0822_, G14[8]);
  or g_1550_(_0821_, _0823_, _0824_);
  or g_1551_(_0813_, _0815_, _0825_);
  and g_1552_(G11[0], G12[9], _0826_);
  or g_1553_(_0785_, _0787_, _0827_);
  and g_1554_(_0826_, _0827_, _0828_);
  xor g_1555_(_0826_, _0827_, _0829_);
  or g_1556_(_0809_, _0811_, _0830_);
  or g_1557_(_0780_, _0782_, _0831_);
  and g_1558_(G11[1], G12[8], _0832_);
  and g_1559_(G11[3], G12[6], _0833_);
  and g_1560_(G11[3], G12[7], _0834_);
  and g_1561_(_0779_, _0833_, _0835_);
  xor g_1562_(_0779_, _0833_, _0836_);
  and g_1563_(_0832_, _0836_, _0837_);
  xor g_1564_(_0832_, _0836_, _0838_);
  or g_1565_(_0793_, _0795_, _0839_);
  and g_1566_(_0838_, _0839_, _0840_);
  xor g_1567_(_0838_, _0839_, _0841_);
  and g_1568_(_0831_, _0841_, _0842_);
  xor g_1569_(_0831_, _0841_, _0843_);
  or g_1570_(_0805_, _0807_, _0844_);
  and g_1571_(G11[4], G12[5], _0845_);
  and g_1572_(G12[2], G11[7], _0846_);
  and g_1573_(G12[4], G11[7], _0847_);
  and g_1574_(_0748_, _0846_, _0848_);
  xor g_1575_(_0748_, _0846_, _0849_);
  and g_1576_(_0845_, _0849_, _0850_);
  xor g_1577_(_0845_, _0849_, _0851_);
  or g_1578_(_0801_, _0803_, _0852_);
  and g_1579_(G12[1], G11[8], _0853_);
  and g_1580_(G12[0], G11[9], _0854_);
  and g_1581_(G12[3], G11[9], _0855_);
  and g_1582_(_0716_, _0854_, _0856_);
  xor g_1583_(_0716_, _0854_, _0857_);
  and g_1584_(_0853_, _0857_, _0858_);
  xor g_1585_(_0853_, _0857_, _0859_);
  and g_1586_(_0852_, _0859_, _0860_);
  xor g_1587_(_0852_, _0859_, _0861_);
  and g_1588_(_0851_, _0861_, _0862_);
  xor g_1589_(_0851_, _0861_, _0863_);
  and g_1590_(_0844_, _0863_, _0864_);
  xor g_1591_(_0844_, _0863_, _0865_);
  and g_1592_(_0843_, _0865_, _0866_);
  xor g_1593_(_0843_, _0865_, _0867_);
  and g_1594_(_0830_, _0867_, _0868_);
  xor g_1595_(_0830_, _0867_, _0869_);
  and g_1596_(_0829_, _0869_, _0870_);
  xor g_1597_(_0829_, _0869_, _0871_);
  and g_1598_(_0825_, _0871_, _0872_);
  xor g_1599_(_0825_, _0871_, _0873_);
  and g_1600_(_0817_, _0873_, _0874_);
  xor g_1601_(_0817_, _0873_, _0875_);
  and g_1602_(_0819_, _0875_, _0876_);
  xor g_1603_(_0819_, _0875_, _0877_);
  and g_1604_(_0824_, _0877_, _0878_);
  xor g_1605_(_0824_, _0877_, G14[9]);
  or g_1606_(_0876_, _0878_, _0879_);
  or g_1607_(_0868_, _0870_, _0880_);
  and g_1608_(G11[0], G12[10], _0881_);
  and g_1609_(G11[1], G12[9], _0882_);
  and g_1610_(G11[1], G12[10], _0883_);
  and g_1611_(_0826_, _0883_, _0884_);
  xor g_1612_(_0881_, _0882_, _0885_);
  or g_1613_(_0840_, _0842_, _0886_);
  and g_1614_(_0885_, _0886_, _0887_);
  xor g_1615_(_0885_, _0886_, _0888_);
  or g_1616_(_0864_, _0866_, _0889_);
  or g_1617_(_0835_, _0837_, _0890_);
  and g_1618_(G11[2], G12[8], _0891_);
  and g_1619_(G11[4], G12[6], _0892_);
  and g_1620_(G11[4], G12[7], _0893_);
  and g_1621_(_0834_, _0892_, _0894_);
  xor g_1622_(_0834_, _0892_, _0895_);
  and g_1623_(_0891_, _0895_, _0896_);
  xor g_1624_(_0891_, _0895_, _0897_);
  or g_1625_(_0848_, _0850_, _0898_);
  and g_1626_(_0897_, _0898_, _0899_);
  xor g_1627_(_0897_, _0898_, _0900_);
  and g_1628_(_0890_, _0900_, _0901_);
  xor g_1629_(_0890_, _0900_, _0902_);
  or g_1630_(_0860_, _0862_, _0903_);
  and g_1631_(G11[5], G12[5], _0904_);
  and g_1632_(G12[2], G11[8], _0905_);
  and g_1633_(G12[4], G11[8], _0906_);
  and g_1634_(_0792_, _0905_, _0907_);
  xor g_1635_(_0792_, _0905_, _0908_);
  and g_1636_(_0904_, _0908_, _0909_);
  xor g_1637_(_0904_, _0908_, _0910_);
  or g_1638_(_0856_, _0858_, _0911_);
  and g_1639_(G12[1], G11[9], _0912_);
  and g_1640_(G12[0], G11[10], _0913_);
  and g_1641_(G12[3], G11[10], _0914_);
  and g_1642_(_0738_, _0914_, _0915_);
  xor g_1643_(_0739_, _0913_, _0916_);
  and g_1644_(_0912_, _0916_, _0917_);
  xor g_1645_(_0912_, _0916_, _0918_);
  and g_1646_(_0911_, _0918_, _0919_);
  xor g_1647_(_0911_, _0918_, _0920_);
  and g_1648_(_0910_, _0920_, _0921_);
  xor g_1649_(_0910_, _0920_, _0922_);
  and g_1650_(_0903_, _0922_, _0923_);
  xor g_1651_(_0903_, _0922_, _0924_);
  and g_1652_(_0902_, _0924_, _0925_);
  xor g_1653_(_0902_, _0924_, _0926_);
  and g_1654_(_0889_, _0926_, _0927_);
  xor g_1655_(_0889_, _0926_, _0928_);
  and g_1656_(_0888_, _0928_, _0929_);
  xor g_1657_(_0888_, _0928_, _0930_);
  and g_1658_(_0880_, _0930_, _0931_);
  xor g_1659_(_0880_, _0930_, _0932_);
  and g_1660_(_0828_, _0932_, _0933_);
  xor g_1661_(_0828_, _0932_, _0934_);
  and g_1662_(_0872_, _0934_, _0935_);
  xor g_1663_(_0872_, _0934_, _0936_);
  and g_1664_(_0874_, _0936_, _0937_);
  xor g_1665_(_0874_, _0936_, _0938_);
  and g_1666_(_0879_, _0938_, _0939_);
  xor g_1667_(_0879_, _0938_, G14[10]);
  or g_1668_(_0937_, _0939_, _0940_);
  or g_1669_(_0931_, _0933_, _0941_);
  or g_1670_(_0927_, _0929_, _0942_);
  and g_1671_(G11[0], G12[11], _0943_);
  and g_1672_(G11[2], G12[9], _0944_);
  and g_1673_(G11[2], G12[10], _0945_);
  and g_1674_(_0883_, _0944_, _0946_);
  xor g_1675_(_0883_, _0944_, _0947_);
  and g_1676_(_0943_, _0947_, _0948_);
  xor g_1677_(_0943_, _0947_, _0949_);
  and g_1678_(_0884_, _0949_, _0950_);
  xor g_1679_(_0884_, _0949_, _0951_);
  or g_1680_(_0899_, _0901_, _0952_);
  and g_1681_(_0951_, _0952_, _0953_);
  xor g_1682_(_0951_, _0952_, _0954_);
  or g_1683_(_0923_, _0925_, _0955_);
  or g_1684_(_0894_, _0896_, _0956_);
  and g_1685_(G11[3], G12[8], _0957_);
  and g_1686_(G11[5], G12[6], _0958_);
  and g_1687_(G11[5], G12[7], _0959_);
  and g_1688_(_0893_, _0958_, _0960_);
  xor g_1689_(_0893_, _0958_, _0961_);
  and g_1690_(_0957_, _0961_, _0962_);
  xor g_1691_(_0957_, _0961_, _0963_);
  or g_1692_(_0907_, _0909_, _0964_);
  and g_1693_(_0963_, _0964_, _0965_);
  xor g_1694_(_0963_, _0964_, _0966_);
  and g_1695_(_0956_, _0966_, _0967_);
  xor g_1696_(_0956_, _0966_, _0968_);
  or g_1697_(_0919_, _0921_, _0969_);
  and g_1698_(G12[5], G11[6], _0970_);
  and g_1699_(G12[2], G11[9], _0971_);
  and g_1700_(G12[4], G11[9], _0972_);
  and g_1701_(_0847_, _0971_, _0973_);
  xor g_1702_(_0847_, _0971_, _0974_);
  and g_1703_(_0970_, _0974_, _0975_);
  xor g_1704_(_0970_, _0974_, _0976_);
  or g_1705_(_0915_, _0917_, _0977_);
  and g_1706_(G12[1], G11[10], _0978_);
  and g_1707_(G12[0], G11[11], _0979_);
  and g_1708_(G12[3], G11[11], _0980_);
  and g_1709_(_0799_, _0980_, _0981_);
  xor g_1710_(_0800_, _0979_, _0982_);
  and g_1711_(_0978_, _0982_, _0983_);
  xor g_1712_(_0978_, _0982_, _0984_);
  and g_1713_(_0977_, _0984_, _0985_);
  xor g_1714_(_0977_, _0984_, _0986_);
  and g_1715_(_0976_, _0986_, _0987_);
  xor g_1716_(_0976_, _0986_, _0988_);
  and g_1717_(_0969_, _0988_, _0989_);
  xor g_1718_(_0969_, _0988_, _0990_);
  and g_1719_(_0968_, _0990_, _0991_);
  xor g_1720_(_0968_, _0990_, _0992_);
  and g_1721_(_0955_, _0992_, _0993_);
  xor g_1722_(_0955_, _0992_, _0994_);
  and g_1723_(_0954_, _0994_, _0995_);
  xor g_1724_(_0954_, _0994_, _0996_);
  and g_1725_(_0942_, _0996_, _0997_);
  xor g_1726_(_0942_, _0996_, _0998_);
  and g_1727_(_0887_, _0998_, _0999_);
  xor g_1728_(_0887_, _0998_, _1000_);
  and g_1729_(_0941_, _1000_, _1001_);
  xor g_1730_(_0941_, _1000_, _1002_);
  and g_1731_(_0935_, _1002_, _1003_);
  xor g_1732_(_0935_, _1002_, _1004_);
  and g_1733_(_0940_, _1004_, _1005_);
  xor g_1734_(_0940_, _1004_, G14[11]);
  or g_1735_(_1003_, _1005_, _1006_);
  or g_1736_(_0997_, _0999_, _1007_);
  or g_1737_(_0993_, _0995_, _1008_);
  and g_1738_(G11[0], G12[12], _1009_);
  or g_1739_(_0946_, _0948_, _1010_);
  and g_1740_(G11[1], G12[11], _1011_);
  and g_1741_(G11[3], G12[9], _1012_);
  and g_1742_(G11[3], G12[10], _1013_);
  and g_1743_(_0945_, _1012_, _1014_);
  xor g_1744_(_0945_, _1012_, _1015_);
  and g_1745_(_1011_, _1015_, _1016_);
  xor g_1746_(_1011_, _1015_, _1017_);
  and g_1747_(_1010_, _1017_, _1018_);
  xor g_1748_(_1010_, _1017_, _1019_);
  and g_1749_(_1009_, _1019_, _1020_);
  xor g_1750_(_1009_, _1019_, _1021_);
  or g_1751_(_0965_, _0967_, _1022_);
  and g_1752_(_1021_, _1022_, _1023_);
  xor g_1753_(_1021_, _1022_, _1024_);
  and g_1754_(_0950_, _1024_, _1025_);
  xor g_1755_(_0950_, _1024_, _1026_);
  or g_1756_(_0989_, _0991_, _1027_);
  or g_1757_(_0960_, _0962_, _1028_);
  and g_1758_(G11[4], G12[8], _1029_);
  and g_1759_(G11[6], G12[6], _1030_);
  and g_1760_(G11[6], G12[7], _1031_);
  and g_1761_(_0959_, _1030_, _1032_);
  xor g_1762_(_0959_, _1030_, _1033_);
  and g_1763_(_1029_, _1033_, _1034_);
  xor g_1764_(_1029_, _1033_, _1035_);
  or g_1765_(_0973_, _0975_, _1036_);
  and g_1766_(_1035_, _1036_, _1037_);
  xor g_1767_(_1035_, _1036_, _1038_);
  and g_1768_(_1028_, _1038_, _1039_);
  xor g_1769_(_1028_, _1038_, _1040_);
  or g_1770_(_0985_, _0987_, _1041_);
  and g_1771_(G12[5], G11[7], _1042_);
  and g_1772_(G12[2], G11[10], _1043_);
  and g_1773_(G12[4], G11[10], _1044_);
  and g_1774_(_0905_, _1044_, _1045_);
  xor g_1775_(_0906_, _1043_, _1046_);
  and g_1776_(_1042_, _1046_, _1047_);
  xor g_1777_(_1042_, _1046_, _1048_);
  or g_1778_(_0981_, _0983_, _1049_);
  and g_1779_(G12[1], G11[11], _1050_);
  and g_1780_(G12[0], G11[12], _1051_);
  and g_1781_(G12[3], G11[12], _1052_);
  and g_1782_(_0854_, _1052_, _1053_);
  xor g_1783_(_0855_, _1051_, _1054_);
  and g_1784_(_1050_, _1054_, _1055_);
  xor g_1785_(_1050_, _1054_, _1056_);
  and g_1786_(_1049_, _1056_, _1057_);
  xor g_1787_(_1049_, _1056_, _1058_);
  and g_1788_(_1048_, _1058_, _1059_);
  xor g_1789_(_1048_, _1058_, _1061_);
  and g_1790_(_1041_, _1061_, _1062_);
  xor g_1791_(_1041_, _1061_, _1063_);
  and g_1792_(_1040_, _1063_, _1064_);
  xor g_1793_(_1040_, _1063_, _1065_);
  and g_1794_(_1027_, _1065_, _1066_);
  xor g_1795_(_1027_, _1065_, _1067_);
  and g_1796_(_1026_, _1067_, _1068_);
  xor g_1797_(_1026_, _1067_, _1069_);
  and g_1798_(_1008_, _1069_, _1070_);
  xor g_1799_(_1008_, _1069_, _1072_);
  and g_1800_(_0953_, _1072_, _1073_);
  xor g_1801_(_0953_, _1072_, _1074_);
  and g_1802_(_1007_, _1074_, _1075_);
  xor g_1803_(_1007_, _1074_, _1076_);
  and g_1804_(_1001_, _1076_, _1077_);
  xor g_1805_(_1001_, _1076_, _1078_);
  and g_1806_(_1006_, _1078_, _1079_);
  xor g_1807_(_1006_, _1078_, G14[12]);
  or g_1808_(_1077_, _1079_, _1080_);
  or g_1809_(_1070_, _1073_, _1082_);
  or g_1810_(_1023_, _1025_, _1083_);
  or g_1811_(_1066_, _1068_, _1084_);
  or g_1812_(_1018_, _1020_, _1085_);
  and g_1813_(G11[0], G12[13], _1086_);
  and g_1814_(G11[1], G12[12], _1087_);
  and g_1815_(G11[1], G12[13], _1088_);
  and g_1816_(_1009_, _1088_, _1089_);
  xor g_1817_(_1086_, _1087_, _1090_);
  or g_1818_(_1014_, _1016_, _1091_);
  and g_1819_(G11[2], G12[11], _1093_);
  and g_1820_(G11[4], G12[9], _1094_);
  and g_1821_(G11[4], G12[10], _1095_);
  and g_1822_(_1013_, _1094_, _1096_);
  xor g_1823_(_1013_, _1094_, _1097_);
  and g_1824_(_1093_, _1097_, _1098_);
  xor g_1825_(_1093_, _1097_, _1099_);
  and g_1826_(_1091_, _1099_, _1100_);
  xor g_1827_(_1091_, _1099_, _1101_);
  and g_1828_(_1090_, _1101_, _1102_);
  xor g_1829_(_1090_, _1101_, _1104_);
  or g_1830_(_1037_, _1039_, _1105_);
  and g_1831_(_1104_, _1105_, _1106_);
  xor g_1832_(_1104_, _1105_, _1107_);
  and g_1833_(_1085_, _1107_, _1108_);
  xor g_1834_(_1085_, _1107_, _1109_);
  or g_1835_(_1062_, _1064_, _1110_);
  or g_1836_(_1032_, _1034_, _1111_);
  and g_1837_(G11[5], G12[8], _1112_);
  and g_1838_(G12[6], G11[7], _1113_);
  and g_1839_(G11[7], G12[7], _1115_);
  and g_1840_(_1031_, _1113_, _1116_);
  xor g_1841_(_1031_, _1113_, _1117_);
  and g_1842_(_1112_, _1117_, _1118_);
  xor g_1843_(_1112_, _1117_, _1119_);
  or g_1844_(_1045_, _1047_, _1120_);
  and g_1845_(_1119_, _1120_, _1121_);
  xor g_1846_(_1119_, _1120_, _1122_);
  and g_1847_(_1111_, _1122_, _1123_);
  xor g_1848_(_1111_, _1122_, _1124_);
  or g_1849_(_1057_, _1059_, _1126_);
  and g_1850_(G12[5], G11[8], _1127_);
  and g_1851_(G12[2], G11[11], _1128_);
  and g_1852_(G12[4], G11[11], _1129_);
  and g_1853_(_0971_, _1129_, _1130_);
  xor g_1854_(_0972_, _1128_, _1131_);
  and g_1855_(_1127_, _1131_, _1132_);
  xor g_1856_(_1127_, _1131_, _1133_);
  or g_1857_(_1053_, _1055_, _1134_);
  and g_1858_(G12[1], G11[12], _1135_);
  and g_1859_(G12[0], G11[13], _1137_);
  and g_1860_(_0914_, _1137_, _1138_);
  xor g_1861_(_0914_, _1137_, _1139_);
  and g_1862_(_1135_, _1139_, _1140_);
  xor g_1863_(_1135_, _1139_, _1141_);
  and g_1864_(_1134_, _1141_, _1142_);
  xor g_1865_(_1134_, _1141_, _1143_);
  and g_1866_(_1133_, _1143_, _1144_);
  xor g_1867_(_1133_, _1143_, _1145_);
  and g_1868_(_1126_, _1145_, _1146_);
  xor g_1869_(_1126_, _1145_, _1147_);
  and g_1870_(_1124_, _1147_, _1148_);
  xor g_1871_(_1124_, _1147_, _1149_);
  and g_1872_(_1110_, _1149_, _1150_);
  xor g_1873_(_1110_, _1149_, _1151_);
  and g_1874_(_1109_, _1151_, _1152_);
  xor g_1875_(_1109_, _1151_, _1153_);
  and g_1876_(_1084_, _1153_, _1154_);
  xor g_1877_(_1084_, _1153_, _1155_);
  and g_1878_(_1083_, _1155_, _1156_);
  xor g_1879_(_1083_, _1155_, _1158_);
  and g_1880_(_1082_, _1158_, _1159_);
  xor g_1881_(_1082_, _1158_, _1160_);
  and g_1882_(_1075_, _1160_, _1161_);
  xor g_1883_(_1075_, _1160_, _1162_);
  and g_1884_(_1080_, _1162_, _1163_);
  xor g_1885_(_1080_, _1162_, G14[13]);
  or g_1886_(_1161_, _1163_, _1164_);
  or g_1887_(_1154_, _1156_, _1165_);
  or g_1888_(_1106_, _1108_, _1166_);
  and g_1889_(_1089_, _1166_, _1168_);
  xor g_1890_(_1089_, _1166_, _1169_);
  or g_1891_(_1150_, _1152_, _1170_);
  or g_1892_(_1100_, _1102_, _1171_);
  and g_1893_(G11[0], G12[14], _1172_);
  and g_1894_(G11[2], G12[12], _1173_);
  and g_1895_(G11[2], G12[13], _1174_);
  and g_1896_(_1087_, _1174_, _1175_);
  xor g_1897_(_1088_, _1173_, _1176_);
  and g_1898_(_1172_, _1176_, _1177_);
  xor g_1899_(_1172_, _1176_, _1179_);
  or g_1900_(_1096_, _1098_, _1180_);
  and g_1901_(G11[3], G12[11], _1181_);
  and g_1902_(G11[5], G12[9], _1182_);
  and g_1903_(G11[5], G12[10], _1183_);
  and g_1904_(_1094_, _1183_, _1184_);
  xor g_1905_(_1095_, _1182_, _1185_);
  and g_1906_(_1181_, _1185_, _1186_);
  xor g_1907_(_1181_, _1185_, _1187_);
  and g_1908_(_1180_, _1187_, _1188_);
  xor g_1909_(_1180_, _1187_, _1190_);
  and g_1910_(_1179_, _1190_, _1191_);
  xor g_1911_(_1179_, _1190_, _1192_);
  or g_1912_(_1121_, _1123_, _1193_);
  and g_1913_(_1192_, _1193_, _1194_);
  xor g_1914_(_1192_, _1193_, _1195_);
  and g_1915_(_1171_, _1195_, _1196_);
  xor g_1916_(_1171_, _1195_, _1197_);
  or g_1917_(_1146_, _1148_, _1198_);
  or g_1918_(_1116_, _1118_, _1199_);
  and g_1919_(G11[6], G12[8], _1201_);
  and g_1920_(G12[6], G11[8], _1202_);
  and g_1921_(G11[8], G12[7], _1203_);
  and g_1922_(_1113_, _1203_, _1204_);
  xor g_1923_(_1115_, _1202_, _1205_);
  and g_1924_(_1201_, _1205_, _1206_);
  xor g_1925_(_1201_, _1205_, _1207_);
  or g_1926_(_1130_, _1132_, _1208_);
  and g_1927_(_1207_, _1208_, _1209_);
  xor g_1928_(_1207_, _1208_, _1210_);
  and g_1929_(_1199_, _1210_, _1212_);
  xor g_1930_(_1199_, _1210_, _1213_);
  or g_1931_(_1142_, _1144_, _1214_);
  and g_1932_(G12[5], G11[9], _1215_);
  and g_1933_(G12[2], G11[12], _1216_);
  and g_1934_(_1044_, _1216_, _1217_);
  xor g_1935_(_1044_, _1216_, _1218_);
  and g_1936_(_1215_, _1218_, _1219_);
  xor g_1937_(_1215_, _1218_, _1220_);
  or g_1938_(_1138_, _1140_, _1221_);
  and g_1939_(G12[1], G11[13], _1223_);
  and g_1940_(G12[0], G11[14], _1224_);
  and g_1941_(_0980_, _1224_, _1225_);
  xor g_1942_(_0980_, _1224_, _1226_);
  and g_1943_(_1223_, _1226_, _1227_);
  xor g_1944_(_1223_, _1226_, _1228_);
  and g_1945_(_1221_, _1228_, _1229_);
  xor g_1946_(_1221_, _1228_, _1230_);
  and g_1947_(_1220_, _1230_, _1231_);
  xor g_1948_(_1220_, _1230_, _1232_);
  and g_1949_(_1214_, _1232_, _1234_);
  xor g_1950_(_1214_, _1232_, _1235_);
  and g_1951_(_1213_, _1235_, _1236_);
  xor g_1952_(_1213_, _1235_, _1237_);
  and g_1953_(_1198_, _1237_, _1238_);
  xor g_1954_(_1198_, _1237_, _1239_);
  and g_1955_(_1197_, _1239_, _1240_);
  xor g_1956_(_1197_, _1239_, _1241_);
  and g_1957_(_1170_, _1241_, _1242_);
  xor g_1958_(_1170_, _1241_, _1243_);
  and g_1959_(_1169_, _1243_, _1245_);
  xor g_1960_(_1169_, _1243_, _1246_);
  and g_1961_(_1165_, _1246_, _1247_);
  xor g_1962_(_1165_, _1246_, _1248_);
  and g_1963_(_1159_, _1248_, _1249_);
  xor g_1964_(_1159_, _1248_, _1250_);
  and g_1965_(_1164_, _1250_, _1251_);
  xor g_1966_(_1164_, _1250_, G14[14]);
  or g_1967_(_1249_, _1251_, _1252_);
  or g_1968_(_1242_, _1245_, _1253_);
  or g_1969_(_1188_, _1191_, _1255_);
  or g_1970_(_1234_, _1236_, _1256_);
  xor g_1971_(_1255_, _1256_, _1257_);
  or g_1972_(_1238_, _1240_, _1258_);
  or g_1973_(_1209_, _1212_, _1259_);
  and g_1974_(G11[1], G12[14], _1260_);
  and g_1975_(G11[6], G12[9], _1261_);
  xor g_1976_(_1183_, _1261_, _1262_);
  and g_1977_(G11[3], G12[12], _1263_);
  xor g_1978_(_1174_, _1263_, _1264_);
  xor g_1979_(_1262_, _1264_, _1266_);
  xor g_1980_(_1260_, _1266_, _1267_);
  or g_1981_(_1184_, _1186_, _1268_);
  and g_1982_(G11[4], G12[11], _1269_);
  xor g_1983_(_1268_, _1269_, _1270_);
  xor g_1984_(_1267_, _1270_, _1271_);
  xor g_1985_(_1259_, _1271_, _1272_);
  and g_1986_(G11[0], G12[15], _1273_);
  or g_1987_(_1175_, _1177_, _1274_);
  xor g_1988_(_1273_, _1274_, _1275_);
  or g_1989_(_1204_, _1206_, _1277_);
  and g_1990_(G12[5], G11[10], _1278_);
  and g_1991_(G12[2], G11[13], _1279_);
  xor g_1992_(_1129_, _1279_, _1280_);
  xor g_1993_(_1278_, _1280_, _1281_);
  or g_1994_(_1217_, _1219_, _1282_);
  and g_1995_(G11[7], G12[8], _1283_);
  and g_1996_(G12[6], G11[9], _1284_);
  xor g_1997_(_1203_, _1284_, _1285_);
  xor g_1998_(_1283_, _1285_, _1286_);
  xor g_1999_(_1282_, _1286_, _1288_);
  or g_2000_(_1225_, _1227_, _1289_);
  and g_2001_(G12[1], G11[14], _1290_);
  and g_2002_(G12[0], G11[15], _1291_);
  xor g_2003_(_1052_, _1291_, _1292_);
  xor g_2004_(_1290_, _1292_, _1293_);
  xor g_2005_(_1289_, _1293_, _1294_);
  xor g_2006_(_1281_, _1294_, _1295_);
  xor g_2007_(_1288_, _1295_, _1296_);
  or g_2008_(_1229_, _1231_, _1297_);
  xor g_2009_(_1272_, _1296_, _1299_);
  xor g_2010_(_1277_, _1297_, _1300_);
  xor g_2011_(_1275_, _1300_, _1301_);
  xor g_2012_(_1299_, _1301_, _1302_);
  or g_2013_(_1194_, _1196_, _1303_);
  xor g_2014_(_1302_, _1303_, _1304_);
  xor g_2015_(_1258_, _1304_, _1305_);
  xor g_2016_(_1257_, _1305_, _1306_);
  xor g_2017_(_1253_, _1306_, _1307_);
  xor g_2018_(_1168_, _1247_, _1308_);
  xor g_2019_(_1307_, _1308_, _1310_);
  xor g_2020_(_1252_, _1310_, G14[15]);
  or g_2021_(_0731_, _0733_, _1311_);
  xor g_2022_(_0772_, _1311_, G14[7]);
  xor g_2023_(_1081_, _1136_, G14[1]);
  xor g_2024_(_1178_, _1189_, G14[2]);

endmodule
