module c499(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491, G492, G493, G494, G495, G496, G497, G498, G499, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491, G492, G493, G494, G495, G496, G497, G498, G499;
  lut lut_gate1(0x6, G1, 350, G468);
  lut lut_gate2(0x4, 351, 353, 350);
  lut lut_gate3(0x8, 281, 352, 351);
  lut lut_gate4(0x4, 254, 345, 352);
  lut lut_gate5(0x9, 359, 354, 353);
  lut lut_gate6(0x6, 358, 355, 354);
  lut lut_gate7(0x6, 357, 356, 355);
  lut lut_gate8(0x8, G33, G41, 356);
  lut lut_gate9(0x9, G9, G13, 357);
  lut lut_gate10(0x9, G1, G5, 358);
  lut lut_gate11(0x6, 363, 360, 359);
  lut lut_gate12(0x6, 362, 361, 360);
  lut lut_gate13(0x6, G23, G24, 361);
  lut lut_gate14(0x9, G21, G22, 362);
  lut lut_gate15(0x6, 365, 364, 363);
  lut lut_gate16(0x6, G19, G20, 364);
  lut lut_gate17(0x9, G17, G18, 365);
  lut lut_gate18(0x9, 232, 367, 366);
  lut lut_gate19(0x6, 231, 368, 367);
  lut lut_gate20(0x6, 370, 369, 368);
  lut lut_gate21(0x8, G34, G41, 369);
  lut lut_gate22(0x9, G14, G10, 370);
  lut lut_gate23(0x9, G6, G2, 231);
  lut lut_gate24(0x6, 236, 233, 232);
  lut lut_gate25(0x6, 235, 234, 233);
  lut lut_gate26(0x6, G32, G31, 234);
  lut lut_gate27(0x9, G30, G29, 235);
  lut lut_gate28(0x6, 238, 237, 236);
  lut lut_gate29(0x6, G28, G27, 237);
  lut lut_gate30(0x9, G26, G25, 238);
  lut lut_gate31(0x6, 242, 240, 239);
  lut lut_gate32(0x6, 241, 360, 240);
  lut lut_gate33(0x8, G36, G41, 241);
  lut lut_gate34(0x9, 243, 233, 242);
  lut lut_gate35(0x6, 245, 244, 243);
  lut lut_gate36(0x6, G16, G12, 244);
  lut lut_gate37(0x9, G8, G4, 245);
  lut lut_gate38(0x9, 252, 247, 246);
  lut lut_gate39(0x6, 251, 248, 247);
  lut lut_gate40(0x6, 250, 249, 248);
  lut lut_gate41(0x8, G35, G41, 249);
  lut lut_gate42(0x9, G15, G11, 250);
  lut lut_gate43(0x9, G7, G3, 251);
  lut lut_gate44(0x6, 236, 363, 252);
  lut lut_gate45(0x8, 366, 353, 253);
  lut lut_gate46(0x1, 268, 255, 254);
  lut lut_gate47(0x6, 261, 256, 255);
  lut lut_gate48(0x6, 260, 257, 256);
  lut lut_gate49(0x6, 259, 258, 257);
  lut lut_gate50(0x6, G7, G8, 258);
  lut lut_gate51(0x9, G6, G5, 259);
  lut lut_gate52(0x8, G40, G41, 260);
  lut lut_gate53(0x9, 265, 262, 261);
  lut lut_gate54(0x6, 264, 263, 262);
  lut lut_gate55(0x6, G15, G16, 263);
  lut lut_gate56(0x9, G14, G13, 264);
  lut lut_gate57(0x6, 267, 266, 265);
  lut lut_gate58(0x6, G28, G32, 266);
  lut lut_gate59(0x9, G24, G20, 267);
  lut lut_gate60(0x9, 274, 269, 268);
  lut lut_gate61(0x6, 273, 270, 269);
  lut lut_gate62(0x6, 272, 271, 270);
  lut lut_gate63(0x8, G39, G41, 271);
  lut lut_gate64(0x9, G27, G31, 272);
  lut lut_gate65(0x9, G23, G19, 273);
  lut lut_gate66(0x6, 278, 275, 274);
  lut lut_gate67(0x6, 277, 276, 275);
  lut lut_gate68(0x6, G3, G4, 276);
  lut lut_gate69(0x9, G2, G1, 277);
  lut lut_gate70(0x6, 280, 279, 278);
  lut lut_gate71(0x6, G11, G12, 279);
  lut lut_gate72(0x9, G10, G9, 280);
  lut lut_gate73(0x4, 289, 282, 281);
  lut lut_gate74(0x9, 288, 283, 282);
  lut lut_gate75(0x6, 287, 284, 283);
  lut lut_gate76(0x6, 286, 285, 284);
  lut lut_gate77(0x8, G37, G41, 285);
  lut lut_gate78(0x9, G25, G29, 286);
  lut lut_gate79(0x9, G21, G17, 287);
  lut lut_gate80(0x6, 275, 257, 288);
  lut lut_gate81(0x9, 295, 290, 289);
  lut lut_gate82(0x6, 294, 291, 290);
  lut lut_gate83(0x6, 293, 292, 291);
  lut lut_gate84(0x8, G38, G41, 292);
  lut lut_gate85(0x9, G26, G30, 293);
  lut lut_gate86(0x9, G22, G18, 294);
  lut lut_gate87(0x6, 278, 262, 295);
  lut lut_gate88(0x6, G2, 296, G469);
  lut lut_gate89(0x4, 351, 366, 296);
  lut lut_gate90(0x6, G3, 297, G470);
  lut lut_gate91(0x4, 351, 246, 297);
  lut lut_gate92(0x6, G4, 298, G471);
  lut lut_gate93(0x8, 239, 351, 298);
  lut lut_gate94(0x6, G5, 299, G472);
  lut lut_gate95(0x4, 300, 353, 299);
  lut lut_gate96(0x8, 281, 301, 300);
  lut lut_gate97(0x4, 302, 345, 301);
  lut lut_gate98(0x8, 268, 255, 302);
  lut lut_gate99(0x6, G6, 303, G473);
  lut lut_gate100(0x4, 300, 366, 303);
  lut lut_gate101(0x6, G7, 304, G474);
  lut lut_gate102(0x4, 300, 246, 304);
  lut lut_gate103(0x6, G8, 305, G475);
  lut lut_gate104(0x8, 239, 300, 305);
  lut lut_gate105(0x6, G9, 306, G476);
  lut lut_gate106(0x4, 307, 353, 306);
  lut lut_gate107(0x8, 308, 352, 307);
  lut lut_gate108(0x4, 282, 289, 308);
  lut lut_gate109(0x6, G10, 309, G477);
  lut lut_gate110(0x4, 307, 366, 309);
  lut lut_gate111(0x6, G11, 310, G478);
  lut lut_gate112(0x4, 307, 246, 310);
  lut lut_gate113(0x6, G12, 311, G479);
  lut lut_gate114(0x8, 239, 307, 311);
  lut lut_gate115(0x6, G13, 312, G480);
  lut lut_gate116(0x4, 313, 353, 312);
  lut lut_gate117(0x8, 308, 301, 313);
  lut lut_gate118(0x6, G14, 314, G481);
  lut lut_gate119(0x4, 313, 366, 314);
  lut lut_gate120(0x6, G15, 315, G482);
  lut lut_gate121(0x4, 313, 246, 315);
  lut lut_gate122(0x6, G16, 316, G483);
  lut lut_gate123(0x8, 239, 313, 316);
  lut lut_gate124(0x6, G17, 317, G484);
  lut lut_gate125(0x4, 318, 282, 317);
  lut lut_gate126(0x8, 322, 319, 318);
  lut lut_gate127(0x4, 321, 347, 319);
  lut lut_gate128(0x8, 289, 282, 320);
  lut lut_gate129(0x4, 366, 353, 321);
  lut lut_gate130(0x1, 246, 239, 322);
  lut lut_gate131(0x6, G18, 323, G485);
  lut lut_gate132(0x4, 318, 289, 323);
  lut lut_gate133(0x6, G19, 324, G486);
  lut lut_gate134(0x4, 318, 268, 324);
  lut lut_gate135(0x6, G20, 325, G487);
  lut lut_gate136(0x8, 255, 318, 325);
  lut lut_gate137(0x6, G21, 326, G488);
  lut lut_gate138(0x4, 327, 282, 326);
  lut lut_gate139(0x8, 328, 319, 327);
  lut lut_gate140(0x8, 246, 239, 328);
  lut lut_gate141(0x6, G22, 329, G489);
  lut lut_gate142(0x4, 327, 289, 329);
  lut lut_gate143(0x6, G23, 330, G490);
  lut lut_gate144(0x4, 327, 268, 330);
  lut lut_gate145(0x6, G24, 331, G491);
  lut lut_gate146(0x8, 255, 327, 331);
  lut lut_gate147(0x6, G25, 332, G492);
  lut lut_gate148(0x4, 333, 282, 332);
  lut lut_gate149(0x8, 322, 334, 333);
  lut lut_gate150(0x4, 335, 347, 334);
  lut lut_gate151(0x4, 353, 366, 335);
  lut lut_gate152(0x6, G26, 336, G493);
  lut lut_gate153(0x4, 333, 289, 336);
  lut lut_gate154(0x6, G27, 337, G494);
  lut lut_gate155(0x4, 333, 268, 337);
  lut lut_gate156(0x6, G28, 338, G495);
  lut lut_gate157(0x8, 255, 333, 338);
  lut lut_gate158(0x6, G29, 339, G496);
  lut lut_gate159(0x4, 340, 282, 339);
  lut lut_gate160(0x8, 328, 334, 340);
  lut lut_gate161(0x6, G30, 341, G497);
  lut lut_gate162(0x4, 340, 289, 341);
  lut lut_gate163(0x6, G31, 342, G498);
  lut lut_gate164(0x4, 340, 268, 342);
  lut lut_gate165(0x6, G32, 343, G499);
  lut lut_gate166(0x8, 255, 340, 343);
  lut lut_gate167(0x8, 253, 246, 344);
  lut lut_gate168(0x5c, 239, 348, 344, 345);
  lut lut_gate169(0x8, 320, 268, 346);
  lut lut_gate170(0x3a, 255, 346, 349, 347);
  lut lut_gate171(0x97, 246, 366, 353, 348);
  lut lut_gate172(0x97, 289, 282, 268, 349);

endmodule
