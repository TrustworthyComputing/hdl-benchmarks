module c17(G1, G16, G17, G2, G3, G4, G5);
  wire 00, 01, 02, 03, 04, 05, 06, 07, 08, 09, 10, 11, 12, 13, 14, 15, 16;
  input G1, G2, G3, G4, G5;
  output G16, G17;
  not g_17_(G3, 11);
  not g_18_(G4, 12);
  or g_19_(11, 12, 07);
  and g_20_(G2, 07, 08);
  or g_21_(G5, G2, 09);
  and g_22_(07, 09, G17);
  and g_23_(G3, G1, 10);
  or g_24_(08, 10, G16);

endmodule
