module c2670(G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, G1014, G1017, G1021, G1026, G1030, G1033, G1036, G1148, G1152, G1159, G1193, G1231, G1237, G1240, G1329, G1336, G1342, G1345, G1348, G1351, G1377, G1478, G1540, G1546, G1563, G1578, G1584, G1650, G1653, G1661, G1663, G1675, G1682, G1683, G1720, G1721, G1722, G1723, G1724, G1725, G1726, G1727, G1734, G1735, G1946, G2418, G2488, G2512, G2515, G2516, G2517, G2520, G2523, G2524, G291, G292, G598, G603, G614, G631, G636, G647, G663, G674, G701, G703, G704, G705, G706, G707, G718, G734, G739, G745, G747, G748, G749, G750, G751, G756, G761, G766, G771, G772, G773, G774, G775, G776, G780, G783, G786, G789, G792, G795, G798, G801, G804, G807, G810, G811, G812, G815, G818, G821, G824, G827;
  input G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594;
  lut lut_gate1(0x00fe, 615, G117, G120, G56, G2570);
  lut lut_gate2(0x3500, G120, G117, G67, G35, 615);
  lut lut_gate3(0x6996, G129, G130, 617, 616, G2583);
  lut lut_gate4(0x6996, G131, G132, G156, G128, 616);
  lut lut_gate5(0x9669, G135, G136, G133, G134, 617);
  lut lut_gate6(0x9, 619, 618, G2582);
  lut lut_gate7(0x9669, G141, G142, G139, G140, 618);
  lut lut_gate8(0x9669, G157, G138, G143, G144, 619);
  lut lut_gate9(0xca, G146, 620, 621, G2557);
  lut lut_gate10(0x35, G145, G109, G79, 620);
  lut lut_gate11(0x35, G145, G99, G89, 621);
  lut lut_gate12(0xca, G146, 622, 623, G2559);
  lut lut_gate13(0x35, G145, G110, G80, 622);
  lut lut_gate14(0x35, G145, G100, G90, 623);
  lut lut_gate15(0xebbe, 628, 625, 624, G29, G2587);
  lut lut_gate16(0x96, 686, G2558, G2557, 624);
  lut lut_gate17(0x53ac, G2559, G146, 627, 626, 625);
  lut lut_gate18(0x35, G145, G114, G84, 626);
  lut lut_gate19(0x35, G145, G104, G94, 627);
  lut lut_gate20(0x9669, 694, 692, 690, 688, 628);
  lut lut_gate21(0xbeeb, 631, 630, 629, G29, G2590);
  lut lut_gate22(0x9, 701, 699, 629);
  lut lut_gate23(0x9669, 703, G2561, G2562, G2566, 630);
  lut lut_gate24(0x6996, G2560, G2572, G2571, G2570, 631);
  lut lut_gate25(0xf, 632, G138, 692, 633, G2591);
  lut lut_gate26(0x001f, 705, 656, 659, 638, 632);
  lut lut_gate27(0x4, 635, 634, 633);
  lut lut_gate28(0x0305, G146, G127, 622, 623, 634);
  lut lut_gate29(0xca00, G30, G146, 620, 621, 635);
  lut lut_gate30(0x4, G136, 694, 636);
  lut lut_gate31(0xbbb0, G135, 688, 694, G136, 637);
  lut lut_gate32(0x00f1, 655, 654, 639, 644, 638);
  lut lut_gate33(0xf800, G8, 640, G2560, 642, 639);
  lut lut_gate34(0x8, G2561, 641, 640);
  lut lut_gate35(0xaccc, 635, 634, G130, G141, 641);
  lut lut_gate36(0xca, 643, G142, G131, 642);
  lut lut_gate37(0x8, 635, 634, 643);
  lut lut_gate38(0x4f00, 652, 650, 648, 645, 644);
  lut lut_gate39(0x0e00, 699, 647, 646, 703, 645);
  lut lut_gate40(0x5333, 635, 634, G126, G138, 646);
  lut lut_gate41(0xaccc, 635, 634, G125, G136, 647);
  lut lut_gate42(0x0777, 703, 646, 649, G2566, 648);
  lut lut_gate43(0x5333, 635, 634, G128, G139, 649);
  lut lut_gate44(0xbbb0, G2566, 649, G2562, 651, 650);
  lut lut_gate45(0x5333, 635, 634, G129, G140, 651);
  lut lut_gate46(0xb0bb, 653, 641, 651, G2562, 652);
  lut lut_gate47(0x4, G8, G2561, 653);
  lut lut_gate48(0x10, G8, G2560, 642, 654);
  lut lut_gate49(0x7000, G8, 643, G2570, G2571, 655);
  lut lut_gate50(0xb, 633, 657, 656);
  lut lut_gate51(0x90, 658, G2572, G134, 657);
  lut lut_gate52(0x07, 636, 688, G135, 658);
  lut lut_gate53(0x0700, G8, 643, G133, G132, 659);
  lut lut_gate54(0x7fff, G141, G142, G139, G140, G2547);
  lut lut_gate55(0x7f, G121, G2, G11, G2548);
  lut lut_gate56(0x7, G7, G121, G2551);
  lut lut_gate57(0xb, G119, G2551, G2552);
  lut lut_gate58(0xb, G147, G2551, G2553);
  lut lut_gate59(0x7, 661, 660, G2554);
  lut lut_gate60(0x8000, G76, G64, G106, G32, 660);
  lut lut_gate61(0x8000, G86, G43, G96, G53, 661);
  lut lut_gate62(0x4f44, G147, 660, G119, 661, G2556);
  lut lut_gate63(0x7, G28, 662, G2564);
  lut lut_gate64(0x10, G116, G121, G2556, 662);
  lut lut_gate65(0x8f, 662, G1, G3, G2565);
  lut lut_gate66(0x3a, G123, G2562, 703, G2573);
  lut lut_gate67(0xac, G123, G2566, G2561, G2575);
  lut lut_gate68(0x44f0, G123, 699, 703, G118, G2578);
  lut lut_gate69(0xbe, G143, 686, G144, G2580);
  lut lut_gate70(0x6f, G10, 665, 663, G2581);
  lut lut_gate71(0x96, G150, G151, 664, 663);
  lut lut_gate72(0x9669, G152, G153, G148, G149, 664);
  lut lut_gate73(0x6996, G154, G155, G125, G126, 665);
  lut lut_gate74(0x5c, G12, G2562, G5, 666);
  lut lut_gate75(0xac, G23, 688, G19, 667);
  lut lut_gate76(0xa3, G23, G2557, G26, 668);
  lut lut_gate77(0x5c, G12, G2561, G15, 669);
  lut lut_gate78(0xc35a, G12, G125, G13, 699, 670);
  lut lut_gate79(0x53, G12, G2572, G18, 671);
  lut lut_gate80(0x3c5a, G12, G132, G17, G2570, 672);
  lut lut_gate81(0xa300, G9, G23, 686, G22, 673);
  lut lut_gate82(0x3ca5, G23, G139, G25, 690, 674);
  lut lut_gate83(0x3ca5, G23, G140, G21, G2559, 675);
  lut lut_gate84(0x3ca5, G23, G136, G24, 694, 676);
  lut lut_gate85(0x3c5a, G12, G133, G6, G2571, 677);
  lut lut_gate86(0xc5, G123, 678, 701, G2588);
  lut lut_gate87(0x96, G2566, 631, 679, 678);
  lut lut_gate88(0x78, 629, G118, 703, 679);
  lut lut_gate89(0x7f, 680, G2590, G2587, G2593);
  lut lut_gate90(0x0100, G2581, G2556, G2582, G2583, 680);
  lut lut_gate91(0x4, G74, G115, G2550);
  lut lut_gate92(0x7, G122, 699, G2563);
  lut lut_gate93(0x4f, 703, G118, G122, G2577);
  lut lut_gate94(0x53, G122, 679, 701, G2586);
  lut lut_gate95(0x1, G2562, G2567);
  lut lut_gate96(0x1, G115, G2531);
  lut lut_gate97(0x1, G124, G2534);
  lut lut_gate98(0x1, G137, G2536);
  lut lut_gate99(0x1, G32, G2539);
  lut lut_gate100(0x1, G106, G2540);
  lut lut_gate101(0x1, G64, G2541);
  lut lut_gate102(0x1, G76, G2542);
  lut lut_gate103(0x1, G53, G2543);
  lut lut_gate104(0x1, G96, G2544);
  lut lut_gate105(0x1, G43, G2545);
  lut lut_gate106(0x1, G86, G2546);
  lut lut_gate107(0x1, G2560, G2569);
  lut lut_gate108(0x1, G2561, G2568);
  lut lut_gate109(0xcfa0, G117, G120, G71, G39, 681);
  lut lut_gate110(0xfc0a, 681, G120, G49, G60, G2566);
  lut lut_gate111(0xcfa0, G117, G120, G66, G34, 682);
  lut lut_gate112(0xfc0a, 682, G120, G45, G55, G2571);
  lut lut_gate113(0xcfa0, G117, G120, G65, G33, 683);
  lut lut_gate114(0xfc0a, 683, G120, G44, G54, G2572);
  lut lut_gate115(0x3f50, G145, G146, G108, G78, 684);
  lut lut_gate116(0xf305, 684, G146, G98, G88, G2558);
  lut lut_gate117(0x3f50, G145, G146, G107, G77, 685);
  lut lut_gate118(0xf305, 685, G146, G97, G87, 686);
  lut lut_gate119(0xcfa0, G145, G146, G105, G75, 687);
  lut lut_gate120(0xfc0a, 687, G146, G95, G85, 688);
  lut lut_gate121(0x3f50, G145, G146, G111, G81, 689);
  lut lut_gate122(0xf305, 689, G146, G101, G91, 690);
  lut lut_gate123(0x3f50, G145, G146, G112, G82, 691);
  lut lut_gate124(0xf305, 691, G146, G102, G92, 692);
  lut lut_gate125(0x3f50, G145, G146, G113, G83, 693);
  lut lut_gate126(0xf305, 693, G146, G103, G93, 694);
  lut lut_gate127(0x3f50, G117, G120, G68, G36, 695);
  lut lut_gate128(0xf305, 695, G120, G46, G57, G2560);
  lut lut_gate129(0x3f50, G117, G120, G70, G38, 696);
  lut lut_gate130(0xf305, 696, G120, G48, G59, G2562);
  lut lut_gate131(0x3f50, G117, G120, G69, G37, 697);
  lut lut_gate132(0xf305, 697, G120, G47, G58, G2561);
  lut lut_gate133(0x3f50, G117, G120, G63, G31, 698);
  lut lut_gate134(0xf305, 698, G120, G42, G52, 699);
  lut lut_gate135(0x3f50, G117, G120, G73, G41, 700);
  lut lut_gate136(0xf305, 700, G120, G51, G62, 701);
  lut lut_gate137(0x3f50, G117, G120, G72, G40, 702);
  lut lut_gate138(0xf305, 702, G120, G50, G61, 703);
  lut lut_gate139(0xf8ff, G2572, G134, G135, 688, 704);
  lut lut_gate140(0x0700, 633, 636, 704, 637, 705);
  lut lut_gate141(0x0990, 666, G129, 667, G135, 706);
  lut lut_gate142(0xa53c, G12, G131, G2560, G16, 707);
  lut lut_gate143(0xa53c, G12, G126, 703, G4, 708);
  lut lut_gate144(0x0100, 673, 675, 674, 672, 709);
  lut lut_gate145(0x1428, 671, 669, G130, G134, 710);
  lut lut_gate146(0x9000, 708, 707, 668, G141, 711);
  lut lut_gate147(0xa5c3, G12, G128, G2566, G14, 712);
  lut lut_gate148(0x8000, 711, 710, 709, 706, 713);
  lut lut_gate149(0xa53c, G23, G138, 692, G20, 714);
  lut lut_gate150(0xa53c, G23, G142, G2558, G27, 715);
  lut lut_gate151(0x1000, 712, 670, 677, 676, 716);
  lut lut_gate152(0x7fff, 713, 716, 715, 714, G2584);

endmodule
