module c1355(G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
  wire 000, 001, 002, 003, 004, 005, 006, 007, 008, 009, 010, 011, 012, 013, 014, 015, 016, 017, 018, 019, 020, 021, 022, 023, 024, 025, 026, 027, 028, 029, 030, 031, 032, 033, 034, 035, 036, 037, 038, 039, 040, 041, 042, 043, 044, 045, 046, 047, 048, 049, 050, 051, 052, 053, 054, 055, 056, 057, 058, 059, 060, 061, 062, 063, 064, 065, 066, 067, 068, 069, 070, 071, 072, 073, 074, 075, 076, 077, 078, 079, 080, 081, 082, 083, 084, 085, 086, 087, 088, 089, 090, 091, 092, 093, 094, 095, 096, 097, 098, 099, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368;
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  lut lut_gate1(0x9, G1, 348, G1324);
  lut lut_gate2(0x4, 349, 351, 348);
  lut lut_gate3(0x8, 279, 350, 349);
  lut lut_gate4(0x4, 252, 343, 350);
  lut lut_gate5(0x9, 357, 352, 351);
  lut lut_gate6(0x6, 356, 353, 352);
  lut lut_gate7(0x6, 355, 354, 353);
  lut lut_gate8(0x8, G33, G41, 354);
  lut lut_gate9(0x9, G9, G13, 355);
  lut lut_gate10(0x9, G1, G5, 356);
  lut lut_gate11(0x6, 361, 358, 357);
  lut lut_gate12(0x6, 360, 359, 358);
  lut lut_gate13(0x6, G23, G24, 359);
  lut lut_gate14(0x9, G21, G22, 360);
  lut lut_gate15(0x6, 363, 362, 361);
  lut lut_gate16(0x6, G19, G20, 362);
  lut lut_gate17(0x9, G17, G18, 363);
  lut lut_gate18(0x9, 230, 365, 364);
  lut lut_gate19(0x6, 229, 366, 365);
  lut lut_gate20(0x6, 368, 367, 366);
  lut lut_gate21(0x8, G34, G41, 367);
  lut lut_gate22(0x9, G14, G10, 368);
  lut lut_gate23(0x9, G6, G2, 229);
  lut lut_gate24(0x6, 234, 231, 230);
  lut lut_gate25(0x6, 233, 232, 231);
  lut lut_gate26(0x6, G32, G31, 232);
  lut lut_gate27(0x9, G30, G29, 233);
  lut lut_gate28(0x6, 236, 235, 234);
  lut lut_gate29(0x6, G28, G27, 235);
  lut lut_gate30(0x9, G26, G25, 236);
  lut lut_gate31(0x6, 240, 238, 237);
  lut lut_gate32(0x6, 239, 358, 238);
  lut lut_gate33(0x8, G36, G41, 239);
  lut lut_gate34(0x9, 241, 231, 240);
  lut lut_gate35(0x6, 243, 242, 241);
  lut lut_gate36(0x6, G16, G12, 242);
  lut lut_gate37(0x9, G8, G4, 243);
  lut lut_gate38(0x9, 250, 245, 244);
  lut lut_gate39(0x6, 249, 246, 245);
  lut lut_gate40(0x6, 248, 247, 246);
  lut lut_gate41(0x8, G35, G41, 247);
  lut lut_gate42(0x9, G15, G11, 248);
  lut lut_gate43(0x9, G7, G3, 249);
  lut lut_gate44(0x6, 234, 361, 250);
  lut lut_gate45(0x8, 364, 351, 251);
  lut lut_gate46(0x1, 266, 253, 252);
  lut lut_gate47(0x6, 259, 254, 253);
  lut lut_gate48(0x6, 258, 255, 254);
  lut lut_gate49(0x6, 257, 256, 255);
  lut lut_gate50(0x6, G7, G8, 256);
  lut lut_gate51(0x9, G6, G5, 257);
  lut lut_gate52(0x8, G40, G41, 258);
  lut lut_gate53(0x9, 263, 260, 259);
  lut lut_gate54(0x6, 262, 261, 260);
  lut lut_gate55(0x6, G15, G16, 261);
  lut lut_gate56(0x9, G14, G13, 262);
  lut lut_gate57(0x6, 265, 264, 263);
  lut lut_gate58(0x6, G28, G32, 264);
  lut lut_gate59(0x9, G24, G20, 265);
  lut lut_gate60(0x9, 272, 267, 266);
  lut lut_gate61(0x6, 271, 268, 267);
  lut lut_gate62(0x6, 270, 269, 268);
  lut lut_gate63(0x8, G39, G41, 269);
  lut lut_gate64(0x9, G27, G31, 270);
  lut lut_gate65(0x9, G23, G19, 271);
  lut lut_gate66(0x6, 276, 273, 272);
  lut lut_gate67(0x6, 275, 274, 273);
  lut lut_gate68(0x6, G3, G4, 274);
  lut lut_gate69(0x9, G2, G1, 275);
  lut lut_gate70(0x6, 278, 277, 276);
  lut lut_gate71(0x6, G11, G12, 277);
  lut lut_gate72(0x9, G10, G9, 278);
  lut lut_gate73(0x4, 287, 280, 279);
  lut lut_gate74(0x9, 286, 281, 280);
  lut lut_gate75(0x6, 285, 282, 281);
  lut lut_gate76(0x6, 284, 283, 282);
  lut lut_gate77(0x8, G37, G41, 283);
  lut lut_gate78(0x9, G25, G29, 284);
  lut lut_gate79(0x9, G21, G17, 285);
  lut lut_gate80(0x6, 273, 255, 286);
  lut lut_gate81(0x9, 293, 288, 287);
  lut lut_gate82(0x6, 292, 289, 288);
  lut lut_gate83(0x6, 291, 290, 289);
  lut lut_gate84(0x8, G38, G41, 290);
  lut lut_gate85(0x9, G26, G30, 291);
  lut lut_gate86(0x9, G22, G18, 292);
  lut lut_gate87(0x6, 276, 260, 293);
  lut lut_gate88(0x9, G2, 294, G1325);
  lut lut_gate89(0x4, 349, 364, 294);
  lut lut_gate90(0x9, G3, 295, G1326);
  lut lut_gate91(0x4, 349, 244, 295);
  lut lut_gate92(0x9, G4, 296, G1327);
  lut lut_gate93(0x8, 237, 349, 296);
  lut lut_gate94(0x9, G5, 297, G1328);
  lut lut_gate95(0x4, 298, 351, 297);
  lut lut_gate96(0x8, 279, 299, 298);
  lut lut_gate97(0x4, 300, 343, 299);
  lut lut_gate98(0x8, 266, 253, 300);
  lut lut_gate99(0x9, G6, 301, G1329);
  lut lut_gate100(0x4, 298, 364, 301);
  lut lut_gate101(0x9, G7, 302, G1330);
  lut lut_gate102(0x4, 298, 244, 302);
  lut lut_gate103(0x9, G8, 303, G1331);
  lut lut_gate104(0x8, 237, 298, 303);
  lut lut_gate105(0x9, G9, 304, G1332);
  lut lut_gate106(0x4, 305, 351, 304);
  lut lut_gate107(0x8, 306, 350, 305);
  lut lut_gate108(0x4, 280, 287, 306);
  lut lut_gate109(0x9, G10, 307, G1333);
  lut lut_gate110(0x4, 305, 364, 307);
  lut lut_gate111(0x9, G11, 308, G1334);
  lut lut_gate112(0x4, 305, 244, 308);
  lut lut_gate113(0x9, G12, 309, G1335);
  lut lut_gate114(0x8, 237, 305, 309);
  lut lut_gate115(0x9, G13, 310, G1336);
  lut lut_gate116(0x4, 311, 351, 310);
  lut lut_gate117(0x8, 306, 299, 311);
  lut lut_gate118(0x9, G14, 312, G1337);
  lut lut_gate119(0x4, 311, 364, 312);
  lut lut_gate120(0x9, G15, 313, G1338);
  lut lut_gate121(0x4, 311, 244, 313);
  lut lut_gate122(0x9, G16, 314, G1339);
  lut lut_gate123(0x8, 237, 311, 314);
  lut lut_gate124(0x9, G17, 315, G1340);
  lut lut_gate125(0x4, 316, 280, 315);
  lut lut_gate126(0x8, 320, 317, 316);
  lut lut_gate127(0x4, 319, 345, 317);
  lut lut_gate128(0x8, 287, 280, 318);
  lut lut_gate129(0x4, 364, 351, 319);
  lut lut_gate130(0x1, 244, 237, 320);
  lut lut_gate131(0x9, G18, 321, G1341);
  lut lut_gate132(0x4, 316, 287, 321);
  lut lut_gate133(0x9, G19, 322, G1342);
  lut lut_gate134(0x4, 316, 266, 322);
  lut lut_gate135(0x9, G20, 323, G1343);
  lut lut_gate136(0x8, 253, 316, 323);
  lut lut_gate137(0x9, G21, 324, G1344);
  lut lut_gate138(0x4, 325, 280, 324);
  lut lut_gate139(0x8, 326, 317, 325);
  lut lut_gate140(0x8, 244, 237, 326);
  lut lut_gate141(0x9, G22, 327, G1345);
  lut lut_gate142(0x4, 325, 287, 327);
  lut lut_gate143(0x9, G23, 328, G1346);
  lut lut_gate144(0x4, 325, 266, 328);
  lut lut_gate145(0x9, G24, 329, G1347);
  lut lut_gate146(0x8, 253, 325, 329);
  lut lut_gate147(0x9, G25, 330, G1348);
  lut lut_gate148(0x4, 331, 280, 330);
  lut lut_gate149(0x8, 320, 332, 331);
  lut lut_gate150(0x4, 333, 345, 332);
  lut lut_gate151(0x4, 351, 364, 333);
  lut lut_gate152(0x9, G26, 334, G1349);
  lut lut_gate153(0x4, 331, 287, 334);
  lut lut_gate154(0x9, G27, 335, G1350);
  lut lut_gate155(0x4, 331, 266, 335);
  lut lut_gate156(0x9, G28, 336, G1351);
  lut lut_gate157(0x8, 253, 331, 336);
  lut lut_gate158(0x9, G29, 337, G1352);
  lut lut_gate159(0x4, 338, 280, 337);
  lut lut_gate160(0x8, 326, 332, 338);
  lut lut_gate161(0x9, G30, 339, G1353);
  lut lut_gate162(0x4, 338, 287, 339);
  lut lut_gate163(0x9, G31, 340, G1354);
  lut lut_gate164(0x4, 338, 266, 340);
  lut lut_gate165(0x9, G32, 341, G1355);
  lut lut_gate166(0x8, 253, 338, 341);
  lut lut_gate167(0x8, 251, 244, 342);
  lut lut_gate168(0x5c, 237, 346, 342, 343);
  lut lut_gate169(0x8, 318, 266, 344);
  lut lut_gate170(0x3a, 253, 344, 347, 345);
  lut lut_gate171(0x97, 244, 364, 351, 346);
  lut lut_gate172(0x97, 287, 280, 266, 347);

endmodule
